magic
tech sky130A
magscale 1 2
timestamp 1657184945
<< obsli1 >>
rect 1104 2159 118864 37553
<< obsm1 >>
rect 658 348 119218 37584
<< metal2 >>
rect 662 0 718 800
rect 2042 0 2098 800
rect 3514 0 3570 800
rect 4894 0 4950 800
rect 6366 0 6422 800
rect 7746 0 7802 800
rect 9218 0 9274 800
rect 10598 0 10654 800
rect 12070 0 12126 800
rect 13450 0 13506 800
rect 14922 0 14978 800
rect 16302 0 16358 800
rect 17774 0 17830 800
rect 19154 0 19210 800
rect 20626 0 20682 800
rect 22006 0 22062 800
rect 23478 0 23534 800
rect 24858 0 24914 800
rect 26330 0 26386 800
rect 27710 0 27766 800
rect 29182 0 29238 800
rect 30654 0 30710 800
rect 32034 0 32090 800
rect 33506 0 33562 800
rect 34886 0 34942 800
rect 36358 0 36414 800
rect 37738 0 37794 800
rect 39210 0 39266 800
rect 40590 0 40646 800
rect 42062 0 42118 800
rect 43442 0 43498 800
rect 44914 0 44970 800
rect 46294 0 46350 800
rect 47766 0 47822 800
rect 49146 0 49202 800
rect 50618 0 50674 800
rect 51998 0 52054 800
rect 53470 0 53526 800
rect 54850 0 54906 800
rect 56322 0 56378 800
rect 57702 0 57758 800
rect 59174 0 59230 800
rect 60646 0 60702 800
rect 62026 0 62082 800
rect 63498 0 63554 800
rect 64878 0 64934 800
rect 66350 0 66406 800
rect 67730 0 67786 800
rect 69202 0 69258 800
rect 70582 0 70638 800
rect 72054 0 72110 800
rect 73434 0 73490 800
rect 74906 0 74962 800
rect 76286 0 76342 800
rect 77758 0 77814 800
rect 79138 0 79194 800
rect 80610 0 80666 800
rect 81990 0 82046 800
rect 83462 0 83518 800
rect 84842 0 84898 800
rect 86314 0 86370 800
rect 87694 0 87750 800
rect 89166 0 89222 800
rect 90638 0 90694 800
rect 92018 0 92074 800
rect 93490 0 93546 800
rect 94870 0 94926 800
rect 96342 0 96398 800
rect 97722 0 97778 800
rect 99194 0 99250 800
rect 100574 0 100630 800
rect 102046 0 102102 800
rect 103426 0 103482 800
rect 104898 0 104954 800
rect 106278 0 106334 800
rect 107750 0 107806 800
rect 109130 0 109186 800
rect 110602 0 110658 800
rect 111982 0 112038 800
rect 113454 0 113510 800
rect 114834 0 114890 800
rect 116306 0 116362 800
rect 117686 0 117742 800
rect 119158 0 119214 800
<< obsm2 >>
rect 664 856 119212 39545
rect 774 342 1986 856
rect 2154 342 3458 856
rect 3626 342 4838 856
rect 5006 342 6310 856
rect 6478 342 7690 856
rect 7858 342 9162 856
rect 9330 342 10542 856
rect 10710 342 12014 856
rect 12182 342 13394 856
rect 13562 342 14866 856
rect 15034 342 16246 856
rect 16414 342 17718 856
rect 17886 342 19098 856
rect 19266 342 20570 856
rect 20738 342 21950 856
rect 22118 342 23422 856
rect 23590 342 24802 856
rect 24970 342 26274 856
rect 26442 342 27654 856
rect 27822 342 29126 856
rect 29294 342 30598 856
rect 30766 342 31978 856
rect 32146 342 33450 856
rect 33618 342 34830 856
rect 34998 342 36302 856
rect 36470 342 37682 856
rect 37850 342 39154 856
rect 39322 342 40534 856
rect 40702 342 42006 856
rect 42174 342 43386 856
rect 43554 342 44858 856
rect 45026 342 46238 856
rect 46406 342 47710 856
rect 47878 342 49090 856
rect 49258 342 50562 856
rect 50730 342 51942 856
rect 52110 342 53414 856
rect 53582 342 54794 856
rect 54962 342 56266 856
rect 56434 342 57646 856
rect 57814 342 59118 856
rect 59286 342 60590 856
rect 60758 342 61970 856
rect 62138 342 63442 856
rect 63610 342 64822 856
rect 64990 342 66294 856
rect 66462 342 67674 856
rect 67842 342 69146 856
rect 69314 342 70526 856
rect 70694 342 71998 856
rect 72166 342 73378 856
rect 73546 342 74850 856
rect 75018 342 76230 856
rect 76398 342 77702 856
rect 77870 342 79082 856
rect 79250 342 80554 856
rect 80722 342 81934 856
rect 82102 342 83406 856
rect 83574 342 84786 856
rect 84954 342 86258 856
rect 86426 342 87638 856
rect 87806 342 89110 856
rect 89278 342 90582 856
rect 90750 342 91962 856
rect 92130 342 93434 856
rect 93602 342 94814 856
rect 94982 342 96286 856
rect 96454 342 97666 856
rect 97834 342 99138 856
rect 99306 342 100518 856
rect 100686 342 101990 856
rect 102158 342 103370 856
rect 103538 342 104842 856
rect 105010 342 106222 856
rect 106390 342 107694 856
rect 107862 342 109074 856
rect 109242 342 110546 856
rect 110714 342 111926 856
rect 112094 342 113398 856
rect 113566 342 114778 856
rect 114946 342 116250 856
rect 116418 342 117630 856
rect 117798 342 119102 856
<< metal3 >>
rect 119200 39448 120000 39568
rect 119200 38496 120000 38616
rect 119200 37544 120000 37664
rect 119200 36592 120000 36712
rect 119200 35640 120000 35760
rect 119200 34688 120000 34808
rect 119200 33872 120000 33992
rect 119200 32920 120000 33040
rect 119200 31968 120000 32088
rect 119200 31016 120000 31136
rect 119200 30064 120000 30184
rect 119200 29112 120000 29232
rect 119200 28296 120000 28416
rect 119200 27344 120000 27464
rect 119200 26392 120000 26512
rect 119200 25440 120000 25560
rect 119200 24488 120000 24608
rect 119200 23536 120000 23656
rect 119200 22720 120000 22840
rect 119200 21768 120000 21888
rect 119200 20816 120000 20936
rect 119200 19864 120000 19984
rect 119200 18912 120000 19032
rect 119200 17960 120000 18080
rect 119200 17144 120000 17264
rect 119200 16192 120000 16312
rect 119200 15240 120000 15360
rect 119200 14288 120000 14408
rect 119200 13336 120000 13456
rect 119200 12384 120000 12504
rect 119200 11568 120000 11688
rect 119200 10616 120000 10736
rect 119200 9664 120000 9784
rect 119200 8712 120000 8832
rect 119200 7760 120000 7880
rect 119200 6808 120000 6928
rect 119200 5992 120000 6112
rect 119200 5040 120000 5160
rect 119200 4088 120000 4208
rect 119200 3136 120000 3256
rect 119200 2184 120000 2304
rect 119200 1232 120000 1352
rect 119200 416 120000 536
<< obsm3 >>
rect 4208 39368 119120 39541
rect 4208 38696 119200 39368
rect 4208 38416 119120 38696
rect 4208 37744 119200 38416
rect 4208 37464 119120 37744
rect 4208 36792 119200 37464
rect 4208 36512 119120 36792
rect 4208 35840 119200 36512
rect 4208 35560 119120 35840
rect 4208 34888 119200 35560
rect 4208 34608 119120 34888
rect 4208 34072 119200 34608
rect 4208 33792 119120 34072
rect 4208 33120 119200 33792
rect 4208 32840 119120 33120
rect 4208 32168 119200 32840
rect 4208 31888 119120 32168
rect 4208 31216 119200 31888
rect 4208 30936 119120 31216
rect 4208 30264 119200 30936
rect 4208 29984 119120 30264
rect 4208 29312 119200 29984
rect 4208 29032 119120 29312
rect 4208 28496 119200 29032
rect 4208 28216 119120 28496
rect 4208 27544 119200 28216
rect 4208 27264 119120 27544
rect 4208 26592 119200 27264
rect 4208 26312 119120 26592
rect 4208 25640 119200 26312
rect 4208 25360 119120 25640
rect 4208 24688 119200 25360
rect 4208 24408 119120 24688
rect 4208 23736 119200 24408
rect 4208 23456 119120 23736
rect 4208 22920 119200 23456
rect 4208 22640 119120 22920
rect 4208 21968 119200 22640
rect 4208 21688 119120 21968
rect 4208 21016 119200 21688
rect 4208 20736 119120 21016
rect 4208 20064 119200 20736
rect 4208 19784 119120 20064
rect 4208 19112 119200 19784
rect 4208 18832 119120 19112
rect 4208 18160 119200 18832
rect 4208 17880 119120 18160
rect 4208 17344 119200 17880
rect 4208 17064 119120 17344
rect 4208 16392 119200 17064
rect 4208 16112 119120 16392
rect 4208 15440 119200 16112
rect 4208 15160 119120 15440
rect 4208 14488 119200 15160
rect 4208 14208 119120 14488
rect 4208 13536 119200 14208
rect 4208 13256 119120 13536
rect 4208 12584 119200 13256
rect 4208 12304 119120 12584
rect 4208 11768 119200 12304
rect 4208 11488 119120 11768
rect 4208 10816 119200 11488
rect 4208 10536 119120 10816
rect 4208 9864 119200 10536
rect 4208 9584 119120 9864
rect 4208 8912 119200 9584
rect 4208 8632 119120 8912
rect 4208 7960 119200 8632
rect 4208 7680 119120 7960
rect 4208 7008 119200 7680
rect 4208 6728 119120 7008
rect 4208 6192 119200 6728
rect 4208 5912 119120 6192
rect 4208 5240 119200 5912
rect 4208 4960 119120 5240
rect 4208 4288 119200 4960
rect 4208 4008 119120 4288
rect 4208 3336 119200 4008
rect 4208 3056 119120 3336
rect 4208 2384 119200 3056
rect 4208 2104 119120 2384
rect 4208 1432 119200 2104
rect 4208 1152 119120 1432
rect 4208 616 119200 1152
rect 4208 443 119120 616
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
rect 65648 2128 65968 37584
rect 81008 2128 81328 37584
rect 96368 2128 96688 37584
rect 111728 2128 112048 37584
<< obsm4 >>
rect 60595 1939 60661 2277
<< labels >>
rlabel metal3 s 119200 1232 120000 1352 6 addr[0]
port 1 nsew signal input
rlabel metal3 s 119200 2184 120000 2304 6 addr[1]
port 2 nsew signal input
rlabel metal3 s 119200 3136 120000 3256 6 addr[2]
port 3 nsew signal input
rlabel metal3 s 119200 4088 120000 4208 6 addr[3]
port 4 nsew signal input
rlabel metal3 s 119200 5040 120000 5160 6 addr[4]
port 5 nsew signal input
rlabel metal3 s 119200 5992 120000 6112 6 addr[5]
port 6 nsew signal input
rlabel metal3 s 119200 6808 120000 6928 6 addr[6]
port 7 nsew signal input
rlabel metal3 s 119200 7760 120000 7880 6 addr[7]
port 8 nsew signal input
rlabel metal3 s 119200 8712 120000 8832 6 addr[8]
port 9 nsew signal input
rlabel metal3 s 119200 9664 120000 9784 6 addr[9]
port 10 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 addr_mem0[0]
port 11 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 addr_mem0[1]
port 12 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 addr_mem0[2]
port 13 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 addr_mem0[3]
port 14 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 addr_mem0[4]
port 15 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 addr_mem0[5]
port 16 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 addr_mem0[6]
port 17 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 addr_mem0[7]
port 18 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 addr_mem0[8]
port 19 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 addr_mem1[0]
port 20 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 addr_mem1[1]
port 21 nsew signal output
rlabel metal2 s 64878 0 64934 800 6 addr_mem1[2]
port 22 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 addr_mem1[3]
port 23 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 addr_mem1[4]
port 24 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 addr_mem1[5]
port 25 nsew signal output
rlabel metal2 s 70582 0 70638 800 6 addr_mem1[6]
port 26 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 addr_mem1[7]
port 27 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 addr_mem1[8]
port 28 nsew signal output
rlabel metal3 s 119200 416 120000 536 6 csb
port 29 nsew signal input
rlabel metal2 s 662 0 718 800 6 csb_mem0
port 30 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 csb_mem1
port 31 nsew signal output
rlabel metal3 s 119200 10616 120000 10736 6 dout[0]
port 32 nsew signal output
rlabel metal3 s 119200 19864 120000 19984 6 dout[10]
port 33 nsew signal output
rlabel metal3 s 119200 20816 120000 20936 6 dout[11]
port 34 nsew signal output
rlabel metal3 s 119200 21768 120000 21888 6 dout[12]
port 35 nsew signal output
rlabel metal3 s 119200 22720 120000 22840 6 dout[13]
port 36 nsew signal output
rlabel metal3 s 119200 23536 120000 23656 6 dout[14]
port 37 nsew signal output
rlabel metal3 s 119200 24488 120000 24608 6 dout[15]
port 38 nsew signal output
rlabel metal3 s 119200 25440 120000 25560 6 dout[16]
port 39 nsew signal output
rlabel metal3 s 119200 26392 120000 26512 6 dout[17]
port 40 nsew signal output
rlabel metal3 s 119200 27344 120000 27464 6 dout[18]
port 41 nsew signal output
rlabel metal3 s 119200 28296 120000 28416 6 dout[19]
port 42 nsew signal output
rlabel metal3 s 119200 11568 120000 11688 6 dout[1]
port 43 nsew signal output
rlabel metal3 s 119200 29112 120000 29232 6 dout[20]
port 44 nsew signal output
rlabel metal3 s 119200 30064 120000 30184 6 dout[21]
port 45 nsew signal output
rlabel metal3 s 119200 31016 120000 31136 6 dout[22]
port 46 nsew signal output
rlabel metal3 s 119200 31968 120000 32088 6 dout[23]
port 47 nsew signal output
rlabel metal3 s 119200 32920 120000 33040 6 dout[24]
port 48 nsew signal output
rlabel metal3 s 119200 33872 120000 33992 6 dout[25]
port 49 nsew signal output
rlabel metal3 s 119200 34688 120000 34808 6 dout[26]
port 50 nsew signal output
rlabel metal3 s 119200 35640 120000 35760 6 dout[27]
port 51 nsew signal output
rlabel metal3 s 119200 36592 120000 36712 6 dout[28]
port 52 nsew signal output
rlabel metal3 s 119200 37544 120000 37664 6 dout[29]
port 53 nsew signal output
rlabel metal3 s 119200 12384 120000 12504 6 dout[2]
port 54 nsew signal output
rlabel metal3 s 119200 38496 120000 38616 6 dout[30]
port 55 nsew signal output
rlabel metal3 s 119200 39448 120000 39568 6 dout[31]
port 56 nsew signal output
rlabel metal3 s 119200 13336 120000 13456 6 dout[3]
port 57 nsew signal output
rlabel metal3 s 119200 14288 120000 14408 6 dout[4]
port 58 nsew signal output
rlabel metal3 s 119200 15240 120000 15360 6 dout[5]
port 59 nsew signal output
rlabel metal3 s 119200 16192 120000 16312 6 dout[6]
port 60 nsew signal output
rlabel metal3 s 119200 17144 120000 17264 6 dout[7]
port 61 nsew signal output
rlabel metal3 s 119200 17960 120000 18080 6 dout[8]
port 62 nsew signal output
rlabel metal3 s 119200 18912 120000 19032 6 dout[9]
port 63 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 dout_mem0[0]
port 64 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 dout_mem0[10]
port 65 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 dout_mem0[11]
port 66 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 dout_mem0[12]
port 67 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 dout_mem0[13]
port 68 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 dout_mem0[14]
port 69 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 dout_mem0[15]
port 70 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 dout_mem0[16]
port 71 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 dout_mem0[17]
port 72 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 dout_mem0[18]
port 73 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 dout_mem0[19]
port 74 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 dout_mem0[1]
port 75 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 dout_mem0[20]
port 76 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 dout_mem0[21]
port 77 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 dout_mem0[22]
port 78 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 dout_mem0[23]
port 79 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 dout_mem0[24]
port 80 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 dout_mem0[25]
port 81 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 dout_mem0[26]
port 82 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 dout_mem0[27]
port 83 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 dout_mem0[28]
port 84 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 dout_mem0[29]
port 85 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 dout_mem0[2]
port 86 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 dout_mem0[30]
port 87 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 dout_mem0[31]
port 88 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 dout_mem0[3]
port 89 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 dout_mem0[4]
port 90 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 dout_mem0[5]
port 91 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 dout_mem0[6]
port 92 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 dout_mem0[7]
port 93 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 dout_mem0[8]
port 94 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 dout_mem0[9]
port 95 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 dout_mem1[0]
port 96 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 dout_mem1[10]
port 97 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 dout_mem1[11]
port 98 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 dout_mem1[12]
port 99 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 dout_mem1[13]
port 100 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 dout_mem1[14]
port 101 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 dout_mem1[15]
port 102 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 dout_mem1[16]
port 103 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 dout_mem1[17]
port 104 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 dout_mem1[18]
port 105 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 dout_mem1[19]
port 106 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 dout_mem1[1]
port 107 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 dout_mem1[20]
port 108 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 dout_mem1[21]
port 109 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 dout_mem1[22]
port 110 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 dout_mem1[23]
port 111 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 dout_mem1[24]
port 112 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 dout_mem1[25]
port 113 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 dout_mem1[26]
port 114 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 dout_mem1[27]
port 115 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 dout_mem1[28]
port 116 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 dout_mem1[29]
port 117 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 dout_mem1[2]
port 118 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 dout_mem1[30]
port 119 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 dout_mem1[31]
port 120 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 dout_mem1[3]
port 121 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 dout_mem1[4]
port 122 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 dout_mem1[5]
port 123 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 dout_mem1[6]
port 124 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 dout_mem1[7]
port 125 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 dout_mem1[8]
port 126 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 dout_mem1[9]
port 127 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 128 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 128 nsew power input
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 128 nsew power input
rlabel metal4 s 96368 2128 96688 37584 6 vccd1
port 128 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 129 nsew ground input
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 129 nsew ground input
rlabel metal4 s 81008 2128 81328 37584 6 vssd1
port 129 nsew ground input
rlabel metal4 s 111728 2128 112048 37584 6 vssd1
port 129 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 120000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1601096
string GDS_FILE /home/leo/Dokumente/caravel_workspace/caravel_wfg/openlane/merge_memory/runs/merge_memory/results/finishing/merge_memory.magic.gds
string GDS_START 62476
<< end >>

