VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wfg_top
  CLASS BLOCK ;
  FOREIGN wfg_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 550.000 ;
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END addr1[8]
  PIN addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END addr1[9]
  PIN csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END csb1
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 4.000 492.280 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END dout1[31]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END dout1[3]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END dout1[4]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END dout1[5]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END dout1[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 546.000 578.590 550.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 546.000 741.430 550.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 546.000 594.690 550.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 546.000 611.250 550.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 546.000 627.350 550.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 546.000 643.450 550.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 546.000 660.010 550.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 546.000 676.110 550.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 546.000 692.670 550.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 546.000 708.770 550.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 546.000 725.330 550.000 ;
    END
  END io_oeb[9]
  PIN io_wbs_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END io_wbs_ack
  PIN io_wbs_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END io_wbs_adr[0]
  PIN io_wbs_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END io_wbs_adr[10]
  PIN io_wbs_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END io_wbs_adr[11]
  PIN io_wbs_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END io_wbs_adr[12]
  PIN io_wbs_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END io_wbs_adr[13]
  PIN io_wbs_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END io_wbs_adr[14]
  PIN io_wbs_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END io_wbs_adr[15]
  PIN io_wbs_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END io_wbs_adr[16]
  PIN io_wbs_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END io_wbs_adr[17]
  PIN io_wbs_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END io_wbs_adr[18]
  PIN io_wbs_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END io_wbs_adr[19]
  PIN io_wbs_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END io_wbs_adr[1]
  PIN io_wbs_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END io_wbs_adr[20]
  PIN io_wbs_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 0.000 510.510 4.000 ;
    END
  END io_wbs_adr[21]
  PIN io_wbs_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END io_wbs_adr[22]
  PIN io_wbs_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END io_wbs_adr[23]
  PIN io_wbs_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END io_wbs_adr[24]
  PIN io_wbs_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 4.000 ;
    END
  END io_wbs_adr[25]
  PIN io_wbs_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END io_wbs_adr[26]
  PIN io_wbs_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END io_wbs_adr[27]
  PIN io_wbs_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 0.000 665.070 4.000 ;
    END
  END io_wbs_adr[28]
  PIN io_wbs_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END io_wbs_adr[29]
  PIN io_wbs_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END io_wbs_adr[2]
  PIN io_wbs_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END io_wbs_adr[30]
  PIN io_wbs_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END io_wbs_adr[31]
  PIN io_wbs_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END io_wbs_adr[3]
  PIN io_wbs_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END io_wbs_adr[4]
  PIN io_wbs_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END io_wbs_adr[5]
  PIN io_wbs_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END io_wbs_adr[6]
  PIN io_wbs_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END io_wbs_adr[7]
  PIN io_wbs_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END io_wbs_adr[8]
  PIN io_wbs_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END io_wbs_adr[9]
  PIN io_wbs_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END io_wbs_clk
  PIN io_wbs_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END io_wbs_cyc
  PIN io_wbs_datrd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END io_wbs_datrd[0]
  PIN io_wbs_datrd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END io_wbs_datrd[10]
  PIN io_wbs_datrd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END io_wbs_datrd[11]
  PIN io_wbs_datrd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END io_wbs_datrd[12]
  PIN io_wbs_datrd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END io_wbs_datrd[13]
  PIN io_wbs_datrd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END io_wbs_datrd[14]
  PIN io_wbs_datrd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END io_wbs_datrd[15]
  PIN io_wbs_datrd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END io_wbs_datrd[16]
  PIN io_wbs_datrd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END io_wbs_datrd[17]
  PIN io_wbs_datrd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END io_wbs_datrd[18]
  PIN io_wbs_datrd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END io_wbs_datrd[19]
  PIN io_wbs_datrd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END io_wbs_datrd[1]
  PIN io_wbs_datrd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END io_wbs_datrd[20]
  PIN io_wbs_datrd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END io_wbs_datrd[21]
  PIN io_wbs_datrd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END io_wbs_datrd[22]
  PIN io_wbs_datrd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END io_wbs_datrd[23]
  PIN io_wbs_datrd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END io_wbs_datrd[24]
  PIN io_wbs_datrd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END io_wbs_datrd[25]
  PIN io_wbs_datrd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END io_wbs_datrd[26]
  PIN io_wbs_datrd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END io_wbs_datrd[27]
  PIN io_wbs_datrd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END io_wbs_datrd[28]
  PIN io_wbs_datrd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END io_wbs_datrd[29]
  PIN io_wbs_datrd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END io_wbs_datrd[2]
  PIN io_wbs_datrd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END io_wbs_datrd[30]
  PIN io_wbs_datrd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END io_wbs_datrd[31]
  PIN io_wbs_datrd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END io_wbs_datrd[3]
  PIN io_wbs_datrd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END io_wbs_datrd[4]
  PIN io_wbs_datrd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END io_wbs_datrd[5]
  PIN io_wbs_datrd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END io_wbs_datrd[6]
  PIN io_wbs_datrd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END io_wbs_datrd[7]
  PIN io_wbs_datrd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END io_wbs_datrd[8]
  PIN io_wbs_datrd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END io_wbs_datrd[9]
  PIN io_wbs_datwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END io_wbs_datwr[0]
  PIN io_wbs_datwr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 0.000 282.810 4.000 ;
    END
  END io_wbs_datwr[10]
  PIN io_wbs_datwr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END io_wbs_datwr[11]
  PIN io_wbs_datwr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END io_wbs_datwr[12]
  PIN io_wbs_datwr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END io_wbs_datwr[13]
  PIN io_wbs_datwr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END io_wbs_datwr[14]
  PIN io_wbs_datwr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END io_wbs_datwr[15]
  PIN io_wbs_datwr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END io_wbs_datwr[16]
  PIN io_wbs_datwr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END io_wbs_datwr[17]
  PIN io_wbs_datwr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END io_wbs_datwr[18]
  PIN io_wbs_datwr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END io_wbs_datwr[19]
  PIN io_wbs_datwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END io_wbs_datwr[1]
  PIN io_wbs_datwr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END io_wbs_datwr[20]
  PIN io_wbs_datwr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END io_wbs_datwr[21]
  PIN io_wbs_datwr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END io_wbs_datwr[22]
  PIN io_wbs_datwr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END io_wbs_datwr[23]
  PIN io_wbs_datwr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END io_wbs_datwr[24]
  PIN io_wbs_datwr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END io_wbs_datwr[25]
  PIN io_wbs_datwr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 4.000 ;
    END
  END io_wbs_datwr[26]
  PIN io_wbs_datwr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END io_wbs_datwr[27]
  PIN io_wbs_datwr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END io_wbs_datwr[28]
  PIN io_wbs_datwr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END io_wbs_datwr[29]
  PIN io_wbs_datwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END io_wbs_datwr[2]
  PIN io_wbs_datwr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END io_wbs_datwr[30]
  PIN io_wbs_datwr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 0.000 746.030 4.000 ;
    END
  END io_wbs_datwr[31]
  PIN io_wbs_datwr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END io_wbs_datwr[3]
  PIN io_wbs_datwr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END io_wbs_datwr[4]
  PIN io_wbs_datwr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END io_wbs_datwr[5]
  PIN io_wbs_datwr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END io_wbs_datwr[6]
  PIN io_wbs_datwr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END io_wbs_datwr[7]
  PIN io_wbs_datwr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END io_wbs_datwr[8]
  PIN io_wbs_datwr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END io_wbs_datwr[9]
  PIN io_wbs_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END io_wbs_rst
  PIN io_wbs_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_wbs_stb
  PIN io_wbs_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END io_wbs_we
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 538.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 538.800 ;
    END
  END vssd1
  PIN wfg_drive_pat_dout_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 546.000 56.950 550.000 ;
    END
  END wfg_drive_pat_dout_o[0]
  PIN wfg_drive_pat_dout_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 546.000 219.790 550.000 ;
    END
  END wfg_drive_pat_dout_o[10]
  PIN wfg_drive_pat_dout_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 546.000 236.350 550.000 ;
    END
  END wfg_drive_pat_dout_o[11]
  PIN wfg_drive_pat_dout_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 546.000 252.450 550.000 ;
    END
  END wfg_drive_pat_dout_o[12]
  PIN wfg_drive_pat_dout_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 546.000 268.550 550.000 ;
    END
  END wfg_drive_pat_dout_o[13]
  PIN wfg_drive_pat_dout_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 546.000 285.110 550.000 ;
    END
  END wfg_drive_pat_dout_o[14]
  PIN wfg_drive_pat_dout_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 546.000 301.210 550.000 ;
    END
  END wfg_drive_pat_dout_o[15]
  PIN wfg_drive_pat_dout_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 546.000 317.770 550.000 ;
    END
  END wfg_drive_pat_dout_o[16]
  PIN wfg_drive_pat_dout_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 546.000 333.870 550.000 ;
    END
  END wfg_drive_pat_dout_o[17]
  PIN wfg_drive_pat_dout_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 546.000 350.430 550.000 ;
    END
  END wfg_drive_pat_dout_o[18]
  PIN wfg_drive_pat_dout_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 546.000 366.530 550.000 ;
    END
  END wfg_drive_pat_dout_o[19]
  PIN wfg_drive_pat_dout_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 546.000 73.050 550.000 ;
    END
  END wfg_drive_pat_dout_o[1]
  PIN wfg_drive_pat_dout_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.810 546.000 383.090 550.000 ;
    END
  END wfg_drive_pat_dout_o[20]
  PIN wfg_drive_pat_dout_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 546.000 399.190 550.000 ;
    END
  END wfg_drive_pat_dout_o[21]
  PIN wfg_drive_pat_dout_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 546.000 415.290 550.000 ;
    END
  END wfg_drive_pat_dout_o[22]
  PIN wfg_drive_pat_dout_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 546.000 431.850 550.000 ;
    END
  END wfg_drive_pat_dout_o[23]
  PIN wfg_drive_pat_dout_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 546.000 447.950 550.000 ;
    END
  END wfg_drive_pat_dout_o[24]
  PIN wfg_drive_pat_dout_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 546.000 464.510 550.000 ;
    END
  END wfg_drive_pat_dout_o[25]
  PIN wfg_drive_pat_dout_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.330 546.000 480.610 550.000 ;
    END
  END wfg_drive_pat_dout_o[26]
  PIN wfg_drive_pat_dout_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 546.000 497.170 550.000 ;
    END
  END wfg_drive_pat_dout_o[27]
  PIN wfg_drive_pat_dout_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 546.000 513.270 550.000 ;
    END
  END wfg_drive_pat_dout_o[28]
  PIN wfg_drive_pat_dout_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 546.000 529.370 550.000 ;
    END
  END wfg_drive_pat_dout_o[29]
  PIN wfg_drive_pat_dout_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 546.000 89.610 550.000 ;
    END
  END wfg_drive_pat_dout_o[2]
  PIN wfg_drive_pat_dout_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 546.000 545.930 550.000 ;
    END
  END wfg_drive_pat_dout_o[30]
  PIN wfg_drive_pat_dout_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 546.000 562.030 550.000 ;
    END
  END wfg_drive_pat_dout_o[31]
  PIN wfg_drive_pat_dout_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 546.000 105.710 550.000 ;
    END
  END wfg_drive_pat_dout_o[3]
  PIN wfg_drive_pat_dout_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 546.000 122.270 550.000 ;
    END
  END wfg_drive_pat_dout_o[4]
  PIN wfg_drive_pat_dout_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 546.000 138.370 550.000 ;
    END
  END wfg_drive_pat_dout_o[5]
  PIN wfg_drive_pat_dout_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 546.000 154.470 550.000 ;
    END
  END wfg_drive_pat_dout_o[6]
  PIN wfg_drive_pat_dout_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 546.000 171.030 550.000 ;
    END
  END wfg_drive_pat_dout_o[7]
  PIN wfg_drive_pat_dout_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 546.000 187.130 550.000 ;
    END
  END wfg_drive_pat_dout_o[8]
  PIN wfg_drive_pat_dout_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 546.000 203.690 550.000 ;
    END
  END wfg_drive_pat_dout_o[9]
  PIN wfg_drive_spi_cs_no
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 546.000 8.190 550.000 ;
    END
  END wfg_drive_spi_cs_no
  PIN wfg_drive_spi_sclk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 546.000 24.290 550.000 ;
    END
  END wfg_drive_spi_sclk_o
  PIN wfg_drive_spi_sdo_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 546.000 40.390 550.000 ;
    END
  END wfg_drive_spi_sdo_o
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 744.280 538.645 ;
      LAYER met1 ;
        RECT 3.290 8.200 746.050 538.800 ;
      LAYER met2 ;
        RECT 3.320 545.720 7.630 546.000 ;
        RECT 8.470 545.720 23.730 546.000 ;
        RECT 24.570 545.720 39.830 546.000 ;
        RECT 40.670 545.720 56.390 546.000 ;
        RECT 57.230 545.720 72.490 546.000 ;
        RECT 73.330 545.720 89.050 546.000 ;
        RECT 89.890 545.720 105.150 546.000 ;
        RECT 105.990 545.720 121.710 546.000 ;
        RECT 122.550 545.720 137.810 546.000 ;
        RECT 138.650 545.720 153.910 546.000 ;
        RECT 154.750 545.720 170.470 546.000 ;
        RECT 171.310 545.720 186.570 546.000 ;
        RECT 187.410 545.720 203.130 546.000 ;
        RECT 203.970 545.720 219.230 546.000 ;
        RECT 220.070 545.720 235.790 546.000 ;
        RECT 236.630 545.720 251.890 546.000 ;
        RECT 252.730 545.720 267.990 546.000 ;
        RECT 268.830 545.720 284.550 546.000 ;
        RECT 285.390 545.720 300.650 546.000 ;
        RECT 301.490 545.720 317.210 546.000 ;
        RECT 318.050 545.720 333.310 546.000 ;
        RECT 334.150 545.720 349.870 546.000 ;
        RECT 350.710 545.720 365.970 546.000 ;
        RECT 366.810 545.720 382.530 546.000 ;
        RECT 383.370 545.720 398.630 546.000 ;
        RECT 399.470 545.720 414.730 546.000 ;
        RECT 415.570 545.720 431.290 546.000 ;
        RECT 432.130 545.720 447.390 546.000 ;
        RECT 448.230 545.720 463.950 546.000 ;
        RECT 464.790 545.720 480.050 546.000 ;
        RECT 480.890 545.720 496.610 546.000 ;
        RECT 497.450 545.720 512.710 546.000 ;
        RECT 513.550 545.720 528.810 546.000 ;
        RECT 529.650 545.720 545.370 546.000 ;
        RECT 546.210 545.720 561.470 546.000 ;
        RECT 562.310 545.720 578.030 546.000 ;
        RECT 578.870 545.720 594.130 546.000 ;
        RECT 594.970 545.720 610.690 546.000 ;
        RECT 611.530 545.720 626.790 546.000 ;
        RECT 627.630 545.720 642.890 546.000 ;
        RECT 643.730 545.720 659.450 546.000 ;
        RECT 660.290 545.720 675.550 546.000 ;
        RECT 676.390 545.720 692.110 546.000 ;
        RECT 692.950 545.720 708.210 546.000 ;
        RECT 709.050 545.720 724.770 546.000 ;
        RECT 725.610 545.720 740.870 546.000 ;
        RECT 741.710 545.720 746.020 546.000 ;
        RECT 3.320 4.280 746.020 545.720 ;
        RECT 3.870 3.670 9.930 4.280 ;
        RECT 10.770 3.670 17.290 4.280 ;
        RECT 18.130 3.670 24.650 4.280 ;
        RECT 25.490 3.670 32.010 4.280 ;
        RECT 32.850 3.670 39.370 4.280 ;
        RECT 40.210 3.670 46.730 4.280 ;
        RECT 47.570 3.670 54.090 4.280 ;
        RECT 54.930 3.670 61.450 4.280 ;
        RECT 62.290 3.670 68.810 4.280 ;
        RECT 69.650 3.670 76.170 4.280 ;
        RECT 77.010 3.670 83.530 4.280 ;
        RECT 84.370 3.670 90.890 4.280 ;
        RECT 91.730 3.670 98.250 4.280 ;
        RECT 99.090 3.670 105.610 4.280 ;
        RECT 106.450 3.670 112.970 4.280 ;
        RECT 113.810 3.670 120.330 4.280 ;
        RECT 121.170 3.670 127.690 4.280 ;
        RECT 128.530 3.670 135.050 4.280 ;
        RECT 135.890 3.670 142.410 4.280 ;
        RECT 143.250 3.670 149.770 4.280 ;
        RECT 150.610 3.670 157.130 4.280 ;
        RECT 157.970 3.670 164.490 4.280 ;
        RECT 165.330 3.670 171.850 4.280 ;
        RECT 172.690 3.670 179.210 4.280 ;
        RECT 180.050 3.670 186.570 4.280 ;
        RECT 187.410 3.670 193.930 4.280 ;
        RECT 194.770 3.670 201.290 4.280 ;
        RECT 202.130 3.670 208.650 4.280 ;
        RECT 209.490 3.670 216.010 4.280 ;
        RECT 216.850 3.670 223.370 4.280 ;
        RECT 224.210 3.670 230.730 4.280 ;
        RECT 231.570 3.670 238.090 4.280 ;
        RECT 238.930 3.670 245.450 4.280 ;
        RECT 246.290 3.670 252.810 4.280 ;
        RECT 253.650 3.670 260.170 4.280 ;
        RECT 261.010 3.670 267.530 4.280 ;
        RECT 268.370 3.670 274.890 4.280 ;
        RECT 275.730 3.670 282.250 4.280 ;
        RECT 283.090 3.670 289.610 4.280 ;
        RECT 290.450 3.670 296.970 4.280 ;
        RECT 297.810 3.670 304.330 4.280 ;
        RECT 305.170 3.670 311.690 4.280 ;
        RECT 312.530 3.670 319.050 4.280 ;
        RECT 319.890 3.670 326.410 4.280 ;
        RECT 327.250 3.670 333.770 4.280 ;
        RECT 334.610 3.670 341.130 4.280 ;
        RECT 341.970 3.670 348.490 4.280 ;
        RECT 349.330 3.670 355.850 4.280 ;
        RECT 356.690 3.670 363.210 4.280 ;
        RECT 364.050 3.670 370.570 4.280 ;
        RECT 371.410 3.670 377.930 4.280 ;
        RECT 378.770 3.670 384.830 4.280 ;
        RECT 385.670 3.670 392.190 4.280 ;
        RECT 393.030 3.670 399.550 4.280 ;
        RECT 400.390 3.670 406.910 4.280 ;
        RECT 407.750 3.670 414.270 4.280 ;
        RECT 415.110 3.670 421.630 4.280 ;
        RECT 422.470 3.670 428.990 4.280 ;
        RECT 429.830 3.670 436.350 4.280 ;
        RECT 437.190 3.670 443.710 4.280 ;
        RECT 444.550 3.670 451.070 4.280 ;
        RECT 451.910 3.670 458.430 4.280 ;
        RECT 459.270 3.670 465.790 4.280 ;
        RECT 466.630 3.670 473.150 4.280 ;
        RECT 473.990 3.670 480.510 4.280 ;
        RECT 481.350 3.670 487.870 4.280 ;
        RECT 488.710 3.670 495.230 4.280 ;
        RECT 496.070 3.670 502.590 4.280 ;
        RECT 503.430 3.670 509.950 4.280 ;
        RECT 510.790 3.670 517.310 4.280 ;
        RECT 518.150 3.670 524.670 4.280 ;
        RECT 525.510 3.670 532.030 4.280 ;
        RECT 532.870 3.670 539.390 4.280 ;
        RECT 540.230 3.670 546.750 4.280 ;
        RECT 547.590 3.670 554.110 4.280 ;
        RECT 554.950 3.670 561.470 4.280 ;
        RECT 562.310 3.670 568.830 4.280 ;
        RECT 569.670 3.670 576.190 4.280 ;
        RECT 577.030 3.670 583.550 4.280 ;
        RECT 584.390 3.670 590.910 4.280 ;
        RECT 591.750 3.670 598.270 4.280 ;
        RECT 599.110 3.670 605.630 4.280 ;
        RECT 606.470 3.670 612.990 4.280 ;
        RECT 613.830 3.670 620.350 4.280 ;
        RECT 621.190 3.670 627.710 4.280 ;
        RECT 628.550 3.670 635.070 4.280 ;
        RECT 635.910 3.670 642.430 4.280 ;
        RECT 643.270 3.670 649.790 4.280 ;
        RECT 650.630 3.670 657.150 4.280 ;
        RECT 657.990 3.670 664.510 4.280 ;
        RECT 665.350 3.670 671.870 4.280 ;
        RECT 672.710 3.670 679.230 4.280 ;
        RECT 680.070 3.670 686.590 4.280 ;
        RECT 687.430 3.670 693.950 4.280 ;
        RECT 694.790 3.670 701.310 4.280 ;
        RECT 702.150 3.670 708.670 4.280 ;
        RECT 709.510 3.670 716.030 4.280 ;
        RECT 716.870 3.670 723.390 4.280 ;
        RECT 724.230 3.670 730.750 4.280 ;
        RECT 731.590 3.670 738.110 4.280 ;
        RECT 738.950 3.670 745.470 4.280 ;
      LAYER met3 ;
        RECT 4.400 542.960 732.715 543.825 ;
        RECT 4.000 531.440 732.715 542.960 ;
        RECT 4.400 530.040 732.715 531.440 ;
        RECT 4.000 518.520 732.715 530.040 ;
        RECT 4.400 517.120 732.715 518.520 ;
        RECT 4.000 505.600 732.715 517.120 ;
        RECT 4.400 504.200 732.715 505.600 ;
        RECT 4.000 492.680 732.715 504.200 ;
        RECT 4.400 491.280 732.715 492.680 ;
        RECT 4.000 480.440 732.715 491.280 ;
        RECT 4.400 479.040 732.715 480.440 ;
        RECT 4.000 467.520 732.715 479.040 ;
        RECT 4.400 466.120 732.715 467.520 ;
        RECT 4.000 454.600 732.715 466.120 ;
        RECT 4.400 453.200 732.715 454.600 ;
        RECT 4.000 441.680 732.715 453.200 ;
        RECT 4.400 440.280 732.715 441.680 ;
        RECT 4.000 428.760 732.715 440.280 ;
        RECT 4.400 427.360 732.715 428.760 ;
        RECT 4.000 416.520 732.715 427.360 ;
        RECT 4.400 415.120 732.715 416.520 ;
        RECT 4.000 403.600 732.715 415.120 ;
        RECT 4.400 402.200 732.715 403.600 ;
        RECT 4.000 390.680 732.715 402.200 ;
        RECT 4.400 389.280 732.715 390.680 ;
        RECT 4.000 377.760 732.715 389.280 ;
        RECT 4.400 376.360 732.715 377.760 ;
        RECT 4.000 364.840 732.715 376.360 ;
        RECT 4.400 363.440 732.715 364.840 ;
        RECT 4.000 351.920 732.715 363.440 ;
        RECT 4.400 350.520 732.715 351.920 ;
        RECT 4.000 339.680 732.715 350.520 ;
        RECT 4.400 338.280 732.715 339.680 ;
        RECT 4.000 326.760 732.715 338.280 ;
        RECT 4.400 325.360 732.715 326.760 ;
        RECT 4.000 313.840 732.715 325.360 ;
        RECT 4.400 312.440 732.715 313.840 ;
        RECT 4.000 300.920 732.715 312.440 ;
        RECT 4.400 299.520 732.715 300.920 ;
        RECT 4.000 288.000 732.715 299.520 ;
        RECT 4.400 286.600 732.715 288.000 ;
        RECT 4.000 275.760 732.715 286.600 ;
        RECT 4.400 274.360 732.715 275.760 ;
        RECT 4.000 262.840 732.715 274.360 ;
        RECT 4.400 261.440 732.715 262.840 ;
        RECT 4.000 249.920 732.715 261.440 ;
        RECT 4.400 248.520 732.715 249.920 ;
        RECT 4.000 237.000 732.715 248.520 ;
        RECT 4.400 235.600 732.715 237.000 ;
        RECT 4.000 224.080 732.715 235.600 ;
        RECT 4.400 222.680 732.715 224.080 ;
        RECT 4.000 211.840 732.715 222.680 ;
        RECT 4.400 210.440 732.715 211.840 ;
        RECT 4.000 198.920 732.715 210.440 ;
        RECT 4.400 197.520 732.715 198.920 ;
        RECT 4.000 186.000 732.715 197.520 ;
        RECT 4.400 184.600 732.715 186.000 ;
        RECT 4.000 173.080 732.715 184.600 ;
        RECT 4.400 171.680 732.715 173.080 ;
        RECT 4.000 160.160 732.715 171.680 ;
        RECT 4.400 158.760 732.715 160.160 ;
        RECT 4.000 147.240 732.715 158.760 ;
        RECT 4.400 145.840 732.715 147.240 ;
        RECT 4.000 135.000 732.715 145.840 ;
        RECT 4.400 133.600 732.715 135.000 ;
        RECT 4.000 122.080 732.715 133.600 ;
        RECT 4.400 120.680 732.715 122.080 ;
        RECT 4.000 109.160 732.715 120.680 ;
        RECT 4.400 107.760 732.715 109.160 ;
        RECT 4.000 96.240 732.715 107.760 ;
        RECT 4.400 94.840 732.715 96.240 ;
        RECT 4.000 83.320 732.715 94.840 ;
        RECT 4.400 81.920 732.715 83.320 ;
        RECT 4.000 71.080 732.715 81.920 ;
        RECT 4.400 69.680 732.715 71.080 ;
        RECT 4.000 58.160 732.715 69.680 ;
        RECT 4.400 56.760 732.715 58.160 ;
        RECT 4.000 45.240 732.715 56.760 ;
        RECT 4.400 43.840 732.715 45.240 ;
        RECT 4.000 32.320 732.715 43.840 ;
        RECT 4.400 30.920 732.715 32.320 ;
        RECT 4.000 19.400 732.715 30.920 ;
        RECT 4.400 18.000 732.715 19.400 ;
        RECT 4.000 7.160 732.715 18.000 ;
        RECT 4.400 6.295 732.715 7.160 ;
      LAYER met4 ;
        RECT 28.815 14.455 97.440 537.025 ;
        RECT 99.840 14.455 174.240 537.025 ;
        RECT 176.640 14.455 251.040 537.025 ;
        RECT 253.440 14.455 327.840 537.025 ;
        RECT 330.240 14.455 404.640 537.025 ;
        RECT 407.040 14.455 481.440 537.025 ;
        RECT 483.840 14.455 558.240 537.025 ;
        RECT 560.640 14.455 635.040 537.025 ;
        RECT 637.440 14.455 647.385 537.025 ;
  END
END wfg_top
END LIBRARY

