magic
tech sky130B
magscale 1 2
timestamp 1657870539
<< nwell >>
rect 1066 37253 148894 37574
rect 1066 36165 148894 36731
rect 1066 35077 148894 35643
rect 1066 33989 148894 34555
rect 1066 32901 148894 33467
rect 1066 31813 148894 32379
rect 1066 30725 148894 31291
rect 1066 29637 148894 30203
rect 1066 28549 148894 29115
rect 1066 27461 148894 28027
rect 1066 26373 148894 26939
rect 1066 25285 148894 25851
rect 1066 24197 148894 24763
rect 1066 23109 148894 23675
rect 1066 22021 148894 22587
rect 1066 20933 148894 21499
rect 1066 19845 148894 20411
rect 1066 18757 148894 19323
rect 1066 17669 148894 18235
rect 1066 16581 148894 17147
rect 1066 15493 148894 16059
rect 1066 14405 148894 14971
rect 1066 13317 148894 13883
rect 1066 12229 148894 12795
rect 1066 11141 148894 11707
rect 1066 10053 148894 10619
rect 1066 8965 148894 9531
rect 1066 7877 148894 8443
rect 1066 6789 148894 7355
rect 1066 5701 148894 6267
rect 1066 4613 148894 5179
rect 1066 3525 148894 4091
rect 1066 2437 148894 3003
<< obsli1 >>
rect 1104 2159 148856 37553
<< obsm1 >>
rect 1104 484 148856 37584
<< metal2 >>
rect 2410 0 2466 800
rect 4158 0 4214 800
rect 5906 0 5962 800
rect 7654 0 7710 800
rect 9402 0 9458 800
rect 11150 0 11206 800
rect 12898 0 12954 800
rect 14646 0 14702 800
rect 16394 0 16450 800
rect 18142 0 18198 800
rect 19890 0 19946 800
rect 21638 0 21694 800
rect 23386 0 23442 800
rect 25134 0 25190 800
rect 26882 0 26938 800
rect 28630 0 28686 800
rect 30378 0 30434 800
rect 32126 0 32182 800
rect 33874 0 33930 800
rect 35622 0 35678 800
rect 37370 0 37426 800
rect 39118 0 39174 800
rect 40866 0 40922 800
rect 42614 0 42670 800
rect 44362 0 44418 800
rect 46110 0 46166 800
rect 47858 0 47914 800
rect 49606 0 49662 800
rect 51354 0 51410 800
rect 53102 0 53158 800
rect 54850 0 54906 800
rect 56598 0 56654 800
rect 58346 0 58402 800
rect 60094 0 60150 800
rect 61842 0 61898 800
rect 63590 0 63646 800
rect 65338 0 65394 800
rect 67086 0 67142 800
rect 68834 0 68890 800
rect 70582 0 70638 800
rect 72330 0 72386 800
rect 74078 0 74134 800
rect 75826 0 75882 800
rect 77574 0 77630 800
rect 79322 0 79378 800
rect 81070 0 81126 800
rect 82818 0 82874 800
rect 84566 0 84622 800
rect 86314 0 86370 800
rect 88062 0 88118 800
rect 89810 0 89866 800
rect 91558 0 91614 800
rect 93306 0 93362 800
rect 95054 0 95110 800
rect 96802 0 96858 800
rect 98550 0 98606 800
rect 100298 0 100354 800
rect 102046 0 102102 800
rect 103794 0 103850 800
rect 105542 0 105598 800
rect 107290 0 107346 800
rect 109038 0 109094 800
rect 110786 0 110842 800
rect 112534 0 112590 800
rect 114282 0 114338 800
rect 116030 0 116086 800
rect 117778 0 117834 800
rect 119526 0 119582 800
rect 121274 0 121330 800
rect 123022 0 123078 800
rect 124770 0 124826 800
rect 126518 0 126574 800
rect 128266 0 128322 800
rect 130014 0 130070 800
rect 131762 0 131818 800
rect 133510 0 133566 800
rect 135258 0 135314 800
rect 137006 0 137062 800
rect 138754 0 138810 800
rect 140502 0 140558 800
rect 142250 0 142306 800
rect 143998 0 144054 800
rect 145746 0 145802 800
rect 147494 0 147550 800
<< obsm2 >>
rect 2412 856 148194 37573
rect 2522 478 4102 856
rect 4270 478 5850 856
rect 6018 478 7598 856
rect 7766 478 9346 856
rect 9514 478 11094 856
rect 11262 478 12842 856
rect 13010 478 14590 856
rect 14758 478 16338 856
rect 16506 478 18086 856
rect 18254 478 19834 856
rect 20002 478 21582 856
rect 21750 478 23330 856
rect 23498 478 25078 856
rect 25246 478 26826 856
rect 26994 478 28574 856
rect 28742 478 30322 856
rect 30490 478 32070 856
rect 32238 478 33818 856
rect 33986 478 35566 856
rect 35734 478 37314 856
rect 37482 478 39062 856
rect 39230 478 40810 856
rect 40978 478 42558 856
rect 42726 478 44306 856
rect 44474 478 46054 856
rect 46222 478 47802 856
rect 47970 478 49550 856
rect 49718 478 51298 856
rect 51466 478 53046 856
rect 53214 478 54794 856
rect 54962 478 56542 856
rect 56710 478 58290 856
rect 58458 478 60038 856
rect 60206 478 61786 856
rect 61954 478 63534 856
rect 63702 478 65282 856
rect 65450 478 67030 856
rect 67198 478 68778 856
rect 68946 478 70526 856
rect 70694 478 72274 856
rect 72442 478 74022 856
rect 74190 478 75770 856
rect 75938 478 77518 856
rect 77686 478 79266 856
rect 79434 478 81014 856
rect 81182 478 82762 856
rect 82930 478 84510 856
rect 84678 478 86258 856
rect 86426 478 88006 856
rect 88174 478 89754 856
rect 89922 478 91502 856
rect 91670 478 93250 856
rect 93418 478 94998 856
rect 95166 478 96746 856
rect 96914 478 98494 856
rect 98662 478 100242 856
rect 100410 478 101990 856
rect 102158 478 103738 856
rect 103906 478 105486 856
rect 105654 478 107234 856
rect 107402 478 108982 856
rect 109150 478 110730 856
rect 110898 478 112478 856
rect 112646 478 114226 856
rect 114394 478 115974 856
rect 116142 478 117722 856
rect 117890 478 119470 856
rect 119638 478 121218 856
rect 121386 478 122966 856
rect 123134 478 124714 856
rect 124882 478 126462 856
rect 126630 478 128210 856
rect 128378 478 129958 856
rect 130126 478 131706 856
rect 131874 478 133454 856
rect 133622 478 135202 856
rect 135370 478 136950 856
rect 137118 478 138698 856
rect 138866 478 140446 856
rect 140614 478 142194 856
rect 142362 478 143942 856
rect 144110 478 145690 856
rect 145858 478 147438 856
rect 147606 478 148194 856
<< metal3 >>
rect 149200 37000 150000 37120
rect 149200 36184 150000 36304
rect 149200 35368 150000 35488
rect 149200 34552 150000 34672
rect 149200 33736 150000 33856
rect 149200 32920 150000 33040
rect 149200 32104 150000 32224
rect 149200 31288 150000 31408
rect 149200 30472 150000 30592
rect 149200 29656 150000 29776
rect 149200 28840 150000 28960
rect 149200 28024 150000 28144
rect 149200 27208 150000 27328
rect 149200 26392 150000 26512
rect 149200 25576 150000 25696
rect 149200 24760 150000 24880
rect 149200 23944 150000 24064
rect 149200 23128 150000 23248
rect 149200 22312 150000 22432
rect 149200 21496 150000 21616
rect 149200 20680 150000 20800
rect 149200 19864 150000 19984
rect 149200 19048 150000 19168
rect 149200 18232 150000 18352
rect 149200 17416 150000 17536
rect 149200 16600 150000 16720
rect 149200 15784 150000 15904
rect 149200 14968 150000 15088
rect 149200 14152 150000 14272
rect 149200 13336 150000 13456
rect 149200 12520 150000 12640
rect 149200 11704 150000 11824
rect 149200 10888 150000 11008
rect 149200 10072 150000 10192
rect 149200 9256 150000 9376
rect 149200 8440 150000 8560
rect 149200 7624 150000 7744
rect 149200 6808 150000 6928
rect 149200 5992 150000 6112
rect 149200 5176 150000 5296
rect 149200 4360 150000 4480
rect 149200 3544 150000 3664
rect 149200 2728 150000 2848
<< obsm3 >>
rect 4210 37200 149200 37569
rect 4210 36920 149120 37200
rect 4210 36384 149200 36920
rect 4210 36104 149120 36384
rect 4210 35568 149200 36104
rect 4210 35288 149120 35568
rect 4210 34752 149200 35288
rect 4210 34472 149120 34752
rect 4210 33936 149200 34472
rect 4210 33656 149120 33936
rect 4210 33120 149200 33656
rect 4210 32840 149120 33120
rect 4210 32304 149200 32840
rect 4210 32024 149120 32304
rect 4210 31488 149200 32024
rect 4210 31208 149120 31488
rect 4210 30672 149200 31208
rect 4210 30392 149120 30672
rect 4210 29856 149200 30392
rect 4210 29576 149120 29856
rect 4210 29040 149200 29576
rect 4210 28760 149120 29040
rect 4210 28224 149200 28760
rect 4210 27944 149120 28224
rect 4210 27408 149200 27944
rect 4210 27128 149120 27408
rect 4210 26592 149200 27128
rect 4210 26312 149120 26592
rect 4210 25776 149200 26312
rect 4210 25496 149120 25776
rect 4210 24960 149200 25496
rect 4210 24680 149120 24960
rect 4210 24144 149200 24680
rect 4210 23864 149120 24144
rect 4210 23328 149200 23864
rect 4210 23048 149120 23328
rect 4210 22512 149200 23048
rect 4210 22232 149120 22512
rect 4210 21696 149200 22232
rect 4210 21416 149120 21696
rect 4210 20880 149200 21416
rect 4210 20600 149120 20880
rect 4210 20064 149200 20600
rect 4210 19784 149120 20064
rect 4210 19248 149200 19784
rect 4210 18968 149120 19248
rect 4210 18432 149200 18968
rect 4210 18152 149120 18432
rect 4210 17616 149200 18152
rect 4210 17336 149120 17616
rect 4210 16800 149200 17336
rect 4210 16520 149120 16800
rect 4210 15984 149200 16520
rect 4210 15704 149120 15984
rect 4210 15168 149200 15704
rect 4210 14888 149120 15168
rect 4210 14352 149200 14888
rect 4210 14072 149120 14352
rect 4210 13536 149200 14072
rect 4210 13256 149120 13536
rect 4210 12720 149200 13256
rect 4210 12440 149120 12720
rect 4210 11904 149200 12440
rect 4210 11624 149120 11904
rect 4210 11088 149200 11624
rect 4210 10808 149120 11088
rect 4210 10272 149200 10808
rect 4210 9992 149120 10272
rect 4210 9456 149200 9992
rect 4210 9176 149120 9456
rect 4210 8640 149200 9176
rect 4210 8360 149120 8640
rect 4210 7824 149200 8360
rect 4210 7544 149120 7824
rect 4210 7008 149200 7544
rect 4210 6728 149120 7008
rect 4210 6192 149200 6728
rect 4210 5912 149120 6192
rect 4210 5376 149200 5912
rect 4210 5096 149120 5376
rect 4210 4560 149200 5096
rect 4210 4280 149120 4560
rect 4210 3744 149200 4280
rect 4210 3464 149120 3744
rect 4210 2928 149200 3464
rect 4210 2648 149120 2928
rect 4210 851 149200 2648
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
rect 65648 2128 65968 37584
rect 81008 2128 81328 37584
rect 96368 2128 96688 37584
rect 111728 2128 112048 37584
rect 127088 2128 127408 37584
rect 142448 2128 142768 37584
<< labels >>
rlabel metal3 s 149200 3544 150000 3664 6 addr[0]
port 1 nsew signal input
rlabel metal3 s 149200 4360 150000 4480 6 addr[1]
port 2 nsew signal input
rlabel metal3 s 149200 5176 150000 5296 6 addr[2]
port 3 nsew signal input
rlabel metal3 s 149200 5992 150000 6112 6 addr[3]
port 4 nsew signal input
rlabel metal3 s 149200 6808 150000 6928 6 addr[4]
port 5 nsew signal input
rlabel metal3 s 149200 7624 150000 7744 6 addr[5]
port 6 nsew signal input
rlabel metal3 s 149200 8440 150000 8560 6 addr[6]
port 7 nsew signal input
rlabel metal3 s 149200 9256 150000 9376 6 addr[7]
port 8 nsew signal input
rlabel metal3 s 149200 10072 150000 10192 6 addr[8]
port 9 nsew signal input
rlabel metal3 s 149200 10888 150000 11008 6 addr[9]
port 10 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 addr_mem0[0]
port 11 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 addr_mem0[1]
port 12 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 addr_mem0[2]
port 13 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 addr_mem0[3]
port 14 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 addr_mem0[4]
port 15 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 addr_mem0[5]
port 16 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 addr_mem0[6]
port 17 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 addr_mem0[7]
port 18 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 addr_mem0[8]
port 19 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 addr_mem1[0]
port 20 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 addr_mem1[1]
port 21 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 addr_mem1[2]
port 22 nsew signal output
rlabel metal2 s 82818 0 82874 800 6 addr_mem1[3]
port 23 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 addr_mem1[4]
port 24 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 addr_mem1[5]
port 25 nsew signal output
rlabel metal2 s 88062 0 88118 800 6 addr_mem1[6]
port 26 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 addr_mem1[7]
port 27 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 addr_mem1[8]
port 28 nsew signal output
rlabel metal3 s 149200 2728 150000 2848 6 csb
port 29 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 csb_mem0
port 30 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 csb_mem1
port 31 nsew signal output
rlabel metal3 s 149200 11704 150000 11824 6 dout[0]
port 32 nsew signal output
rlabel metal3 s 149200 19864 150000 19984 6 dout[10]
port 33 nsew signal output
rlabel metal3 s 149200 20680 150000 20800 6 dout[11]
port 34 nsew signal output
rlabel metal3 s 149200 21496 150000 21616 6 dout[12]
port 35 nsew signal output
rlabel metal3 s 149200 22312 150000 22432 6 dout[13]
port 36 nsew signal output
rlabel metal3 s 149200 23128 150000 23248 6 dout[14]
port 37 nsew signal output
rlabel metal3 s 149200 23944 150000 24064 6 dout[15]
port 38 nsew signal output
rlabel metal3 s 149200 24760 150000 24880 6 dout[16]
port 39 nsew signal output
rlabel metal3 s 149200 25576 150000 25696 6 dout[17]
port 40 nsew signal output
rlabel metal3 s 149200 26392 150000 26512 6 dout[18]
port 41 nsew signal output
rlabel metal3 s 149200 27208 150000 27328 6 dout[19]
port 42 nsew signal output
rlabel metal3 s 149200 12520 150000 12640 6 dout[1]
port 43 nsew signal output
rlabel metal3 s 149200 28024 150000 28144 6 dout[20]
port 44 nsew signal output
rlabel metal3 s 149200 28840 150000 28960 6 dout[21]
port 45 nsew signal output
rlabel metal3 s 149200 29656 150000 29776 6 dout[22]
port 46 nsew signal output
rlabel metal3 s 149200 30472 150000 30592 6 dout[23]
port 47 nsew signal output
rlabel metal3 s 149200 31288 150000 31408 6 dout[24]
port 48 nsew signal output
rlabel metal3 s 149200 32104 150000 32224 6 dout[25]
port 49 nsew signal output
rlabel metal3 s 149200 32920 150000 33040 6 dout[26]
port 50 nsew signal output
rlabel metal3 s 149200 33736 150000 33856 6 dout[27]
port 51 nsew signal output
rlabel metal3 s 149200 34552 150000 34672 6 dout[28]
port 52 nsew signal output
rlabel metal3 s 149200 35368 150000 35488 6 dout[29]
port 53 nsew signal output
rlabel metal3 s 149200 13336 150000 13456 6 dout[2]
port 54 nsew signal output
rlabel metal3 s 149200 36184 150000 36304 6 dout[30]
port 55 nsew signal output
rlabel metal3 s 149200 37000 150000 37120 6 dout[31]
port 56 nsew signal output
rlabel metal3 s 149200 14152 150000 14272 6 dout[3]
port 57 nsew signal output
rlabel metal3 s 149200 14968 150000 15088 6 dout[4]
port 58 nsew signal output
rlabel metal3 s 149200 15784 150000 15904 6 dout[5]
port 59 nsew signal output
rlabel metal3 s 149200 16600 150000 16720 6 dout[6]
port 60 nsew signal output
rlabel metal3 s 149200 17416 150000 17536 6 dout[7]
port 61 nsew signal output
rlabel metal3 s 149200 18232 150000 18352 6 dout[8]
port 62 nsew signal output
rlabel metal3 s 149200 19048 150000 19168 6 dout[9]
port 63 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 dout_mem0[0]
port 64 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 dout_mem0[10]
port 65 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 dout_mem0[11]
port 66 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 dout_mem0[12]
port 67 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 dout_mem0[13]
port 68 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 dout_mem0[14]
port 69 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 dout_mem0[15]
port 70 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 dout_mem0[16]
port 71 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 dout_mem0[17]
port 72 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 dout_mem0[18]
port 73 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 dout_mem0[19]
port 74 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 dout_mem0[1]
port 75 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 dout_mem0[20]
port 76 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 dout_mem0[21]
port 77 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 dout_mem0[22]
port 78 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 dout_mem0[23]
port 79 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 dout_mem0[24]
port 80 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 dout_mem0[25]
port 81 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 dout_mem0[26]
port 82 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 dout_mem0[27]
port 83 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 dout_mem0[28]
port 84 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 dout_mem0[29]
port 85 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 dout_mem0[2]
port 86 nsew signal input
rlabel metal2 s 72330 0 72386 800 6 dout_mem0[30]
port 87 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 dout_mem0[31]
port 88 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 dout_mem0[3]
port 89 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 dout_mem0[4]
port 90 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 dout_mem0[5]
port 91 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 dout_mem0[6]
port 92 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 dout_mem0[7]
port 93 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 dout_mem0[8]
port 94 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 dout_mem0[9]
port 95 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 dout_mem1[0]
port 96 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 dout_mem1[10]
port 97 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 dout_mem1[11]
port 98 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 dout_mem1[12]
port 99 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 dout_mem1[13]
port 100 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 dout_mem1[14]
port 101 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 dout_mem1[15]
port 102 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 dout_mem1[16]
port 103 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 dout_mem1[17]
port 104 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 dout_mem1[18]
port 105 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 dout_mem1[19]
port 106 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 dout_mem1[1]
port 107 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 dout_mem1[20]
port 108 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 dout_mem1[21]
port 109 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 dout_mem1[22]
port 110 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 dout_mem1[23]
port 111 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 dout_mem1[24]
port 112 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 dout_mem1[25]
port 113 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 dout_mem1[26]
port 114 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 dout_mem1[27]
port 115 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 dout_mem1[28]
port 116 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 dout_mem1[29]
port 117 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 dout_mem1[2]
port 118 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 dout_mem1[30]
port 119 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 dout_mem1[31]
port 120 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 dout_mem1[3]
port 121 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 dout_mem1[4]
port 122 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 dout_mem1[5]
port 123 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 dout_mem1[6]
port 124 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 dout_mem1[7]
port 125 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 dout_mem1[8]
port 126 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 dout_mem1[9]
port 127 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 128 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 128 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 128 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 37584 6 vccd1
port 128 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 37584 6 vccd1
port 128 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 129 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 129 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 37584 6 vssd1
port 129 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 37584 6 vssd1
port 129 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 37584 6 vssd1
port 129 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 150000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1911542
string GDS_FILE /home/leo/Dokumente/caravel_workspace_mpw7/caravel_wfg/openlane/merge_memory/runs/22_07_15_09_34/results/signoff/merge_memory.magic.gds
string GDS_START 56722
<< end >>

