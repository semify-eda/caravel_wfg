magic
tech sky130A
magscale 1 2
timestamp 1657004106
<< viali >>
rect 1593 19465 1627 19499
rect 2329 19465 2363 19499
rect 3985 19465 4019 19499
rect 5181 19465 5215 19499
rect 6653 19465 6687 19499
rect 8033 19465 8067 19499
rect 9505 19465 9539 19499
rect 10885 19465 10919 19499
rect 12357 19465 12391 19499
rect 14289 19465 14323 19499
rect 16681 19465 16715 19499
rect 20729 19465 20763 19499
rect 22109 19465 22143 19499
rect 26985 19465 27019 19499
rect 29561 19465 29595 19499
rect 30757 19465 30791 19499
rect 32137 19465 32171 19499
rect 33609 19465 33643 19499
rect 34989 19465 35023 19499
rect 39865 19465 39899 19499
rect 40693 19465 40727 19499
rect 42441 19465 42475 19499
rect 43545 19465 43579 19499
rect 45017 19465 45051 19499
rect 49249 19465 49283 19499
rect 50721 19465 50755 19499
rect 53205 19465 53239 19499
rect 53849 19465 53883 19499
rect 54677 19465 54711 19499
rect 56517 19465 56551 19499
rect 58081 19465 58115 19499
rect 1409 19329 1443 19363
rect 2145 19329 2179 19363
rect 3801 19329 3835 19363
rect 4997 19329 5031 19363
rect 6469 19329 6503 19363
rect 7849 19329 7883 19363
rect 9321 19329 9355 19363
rect 10701 19329 10735 19363
rect 12173 19329 12207 19363
rect 14105 19329 14139 19363
rect 15209 19329 15243 19363
rect 16865 19329 16899 19363
rect 18061 19329 18095 19363
rect 19441 19329 19475 19363
rect 20913 19329 20947 19363
rect 22293 19329 22327 19363
rect 23765 19329 23799 19363
rect 25145 19329 25179 19363
rect 27169 19329 27203 19363
rect 27997 19329 28031 19363
rect 29745 19329 29779 19363
rect 30941 19329 30975 19363
rect 32321 19329 32355 19363
rect 33793 19329 33827 19363
rect 35173 19329 35207 19363
rect 36645 19329 36679 19363
rect 38025 19329 38059 19363
rect 40049 19329 40083 19363
rect 40877 19329 40911 19363
rect 42625 19329 42659 19363
rect 43729 19329 43763 19363
rect 45201 19329 45235 19363
rect 46581 19329 46615 19363
rect 48053 19329 48087 19363
rect 49433 19329 49467 19363
rect 50905 19329 50939 19363
rect 52193 19329 52227 19363
rect 53389 19329 53423 19363
rect 54033 19329 54067 19363
rect 54493 19329 54527 19363
rect 55597 19329 55631 19363
rect 56333 19329 56367 19363
rect 57069 19329 57103 19363
rect 57897 19329 57931 19363
rect 55781 19193 55815 19227
rect 15025 19125 15059 19159
rect 17877 19125 17911 19159
rect 19257 19125 19291 19159
rect 23581 19125 23615 19159
rect 24961 19125 24995 19159
rect 27813 19125 27847 19159
rect 36461 19125 36495 19159
rect 37841 19125 37875 19159
rect 46397 19125 46431 19159
rect 47869 19125 47903 19159
rect 52009 19125 52043 19159
rect 57253 19125 57287 19159
rect 53205 18921 53239 18955
rect 54585 18921 54619 18955
rect 51457 18785 51491 18819
rect 52653 18785 52687 18819
rect 53757 18785 53791 18819
rect 55965 18785 55999 18819
rect 57069 18785 57103 18819
rect 51181 18717 51215 18751
rect 52469 18717 52503 18751
rect 54769 18717 54803 18751
rect 57897 18717 57931 18751
rect 55781 18649 55815 18683
rect 56977 18649 57011 18683
rect 50813 18581 50847 18615
rect 51273 18581 51307 18615
rect 52009 18581 52043 18615
rect 52377 18581 52411 18615
rect 53573 18581 53607 18615
rect 53665 18581 53699 18615
rect 55321 18581 55355 18615
rect 55689 18581 55723 18615
rect 56517 18581 56551 18615
rect 56885 18581 56919 18615
rect 58081 18581 58115 18615
rect 51549 18377 51583 18411
rect 53573 18377 53607 18411
rect 54585 18377 54619 18411
rect 56057 18377 56091 18411
rect 57069 18309 57103 18343
rect 51733 18241 51767 18275
rect 52929 18241 52963 18275
rect 53757 18241 53791 18275
rect 54769 18241 54803 18275
rect 55413 18241 55447 18275
rect 55873 18241 55907 18275
rect 56977 18241 57011 18275
rect 57897 18241 57931 18275
rect 57161 18173 57195 18207
rect 52745 18105 52779 18139
rect 55229 18105 55263 18139
rect 56609 18037 56643 18071
rect 58081 18037 58115 18071
rect 47961 17833 47995 17867
rect 55873 17833 55907 17867
rect 56609 17833 56643 17867
rect 57161 17833 57195 17867
rect 48605 17765 48639 17799
rect 49157 17697 49191 17731
rect 57713 17697 57747 17731
rect 46949 17629 46983 17663
rect 48145 17629 48179 17663
rect 48973 17629 49007 17663
rect 50353 17629 50387 17663
rect 56425 17629 56459 17663
rect 55781 17561 55815 17595
rect 57621 17561 57655 17595
rect 46765 17493 46799 17527
rect 49065 17493 49099 17527
rect 50169 17493 50203 17527
rect 57529 17493 57563 17527
rect 46029 17289 46063 17323
rect 46397 17289 46431 17323
rect 47593 17289 47627 17323
rect 47961 17289 47995 17323
rect 44925 17153 44959 17187
rect 56609 17153 56643 17187
rect 57069 17153 57103 17187
rect 57897 17153 57931 17187
rect 46489 17085 46523 17119
rect 46581 17085 46615 17119
rect 48053 17085 48087 17119
rect 48237 17085 48271 17119
rect 56425 17017 56459 17051
rect 57253 17017 57287 17051
rect 45017 16949 45051 16983
rect 58081 16949 58115 16983
rect 57253 16745 57287 16779
rect 44097 16609 44131 16643
rect 44281 16609 44315 16643
rect 45477 16609 45511 16643
rect 45569 16609 45603 16643
rect 44005 16541 44039 16575
rect 45385 16541 45419 16575
rect 46397 16541 46431 16575
rect 56793 16541 56827 16575
rect 57437 16541 57471 16575
rect 57897 16541 57931 16575
rect 43637 16405 43671 16439
rect 45017 16405 45051 16439
rect 46213 16405 46247 16439
rect 56609 16405 56643 16439
rect 58081 16405 58115 16439
rect 57161 16201 57195 16235
rect 44557 16065 44591 16099
rect 57345 16065 57379 16099
rect 57897 16065 57931 16099
rect 44373 15861 44407 15895
rect 58081 15861 58115 15895
rect 42073 15521 42107 15555
rect 41889 15453 41923 15487
rect 57897 15453 57931 15487
rect 41521 15317 41555 15351
rect 41981 15317 42015 15351
rect 58081 15317 58115 15351
rect 39313 15113 39347 15147
rect 39405 14977 39439 15011
rect 41337 14977 41371 15011
rect 42717 14977 42751 15011
rect 57897 14977 57931 15011
rect 39589 14909 39623 14943
rect 41061 14909 41095 14943
rect 42441 14909 42475 14943
rect 38945 14773 38979 14807
rect 58081 14773 58115 14807
rect 41153 14569 41187 14603
rect 38117 14433 38151 14467
rect 39865 14433 39899 14467
rect 41797 14433 41831 14467
rect 37841 14365 37875 14399
rect 40141 14365 40175 14399
rect 57897 14365 57931 14399
rect 41521 14297 41555 14331
rect 37473 14229 37507 14263
rect 37933 14229 37967 14263
rect 41613 14229 41647 14263
rect 58081 14229 58115 14263
rect 58081 14025 58115 14059
rect 38209 13889 38243 13923
rect 57897 13889 57931 13923
rect 38485 13821 38519 13855
rect 36093 13413 36127 13447
rect 36737 13345 36771 13379
rect 37289 13345 37323 13379
rect 36461 13277 36495 13311
rect 37565 13277 37599 13311
rect 57897 13277 57931 13311
rect 36553 13141 36587 13175
rect 58081 13141 58115 13175
rect 38301 12937 38335 12971
rect 35173 12801 35207 12835
rect 38209 12801 38243 12835
rect 57437 12801 57471 12835
rect 57897 12801 57931 12835
rect 35357 12665 35391 12699
rect 58081 12597 58115 12631
rect 34713 12393 34747 12427
rect 31401 12325 31435 12359
rect 33977 12257 34011 12291
rect 35265 12257 35299 12291
rect 33701 12189 33735 12223
rect 35081 12189 35115 12223
rect 38669 12189 38703 12223
rect 57897 12189 57931 12223
rect 31217 12121 31251 12155
rect 32597 12121 32631 12155
rect 32781 12121 32815 12155
rect 33333 12053 33367 12087
rect 33793 12053 33827 12087
rect 35173 12053 35207 12087
rect 38853 12053 38887 12087
rect 58081 12053 58115 12087
rect 29837 11849 29871 11883
rect 30665 11849 30699 11883
rect 31033 11849 31067 11883
rect 32137 11849 32171 11883
rect 32505 11849 32539 11883
rect 34069 11781 34103 11815
rect 34253 11781 34287 11815
rect 57897 11713 57931 11747
rect 29929 11645 29963 11679
rect 30113 11645 30147 11679
rect 31125 11645 31159 11679
rect 31217 11645 31251 11679
rect 32597 11645 32631 11679
rect 32781 11645 32815 11679
rect 29469 11509 29503 11543
rect 58081 11509 58115 11543
rect 31033 11305 31067 11339
rect 58081 11237 58115 11271
rect 30205 11101 30239 11135
rect 30389 11101 30423 11135
rect 39865 11101 39899 11135
rect 57897 11101 57931 11135
rect 30941 11033 30975 11067
rect 40141 11033 40175 11067
rect 57069 10625 57103 10659
rect 57897 10625 57931 10659
rect 57253 10421 57287 10455
rect 58081 10421 58115 10455
rect 28089 10217 28123 10251
rect 27077 10013 27111 10047
rect 57897 10013 57931 10047
rect 26893 9945 26927 9979
rect 27997 9945 28031 9979
rect 57529 9877 57563 9911
rect 58081 9877 58115 9911
rect 26985 9673 27019 9707
rect 24961 9605 24995 9639
rect 26065 9605 26099 9639
rect 27353 9605 27387 9639
rect 25881 9537 25915 9571
rect 57897 9537 57931 9571
rect 25053 9469 25087 9503
rect 25145 9469 25179 9503
rect 27445 9469 27479 9503
rect 27537 9469 27571 9503
rect 24593 9401 24627 9435
rect 58081 9333 58115 9367
rect 10609 9129 10643 9163
rect 12081 9129 12115 9163
rect 14105 9129 14139 9163
rect 27169 9129 27203 9163
rect 24593 9061 24627 9095
rect 9413 8993 9447 9027
rect 22845 8993 22879 9027
rect 26709 8993 26743 9027
rect 27721 8993 27755 9027
rect 9137 8925 9171 8959
rect 10793 8925 10827 8959
rect 12265 8925 12299 8959
rect 14289 8925 14323 8959
rect 22569 8925 22603 8959
rect 24409 8925 24443 8959
rect 27537 8925 27571 8959
rect 57897 8925 57931 8959
rect 26525 8857 26559 8891
rect 22201 8789 22235 8823
rect 22661 8789 22695 8823
rect 27629 8789 27663 8823
rect 58081 8789 58115 8823
rect 9505 8585 9539 8619
rect 23213 8585 23247 8619
rect 23581 8585 23615 8619
rect 57437 8585 57471 8619
rect 9689 8449 9723 8483
rect 13645 8449 13679 8483
rect 22477 8449 22511 8483
rect 57897 8449 57931 8483
rect 23673 8381 23707 8415
rect 23765 8381 23799 8415
rect 22661 8313 22695 8347
rect 58081 8313 58115 8347
rect 13461 8245 13495 8279
rect 9873 8041 9907 8075
rect 10977 8041 11011 8075
rect 12541 8041 12575 8075
rect 13461 8041 13495 8075
rect 21005 8041 21039 8075
rect 9781 7973 9815 8007
rect 10241 7973 10275 8007
rect 10885 7973 10919 8007
rect 12357 7973 12391 8007
rect 13369 7973 13403 8007
rect 10517 7905 10551 7939
rect 12081 7905 12115 7939
rect 13001 7905 13035 7939
rect 9413 7837 9447 7871
rect 20821 7837 20855 7871
rect 57897 7837 57931 7871
rect 19901 7769 19935 7803
rect 19993 7701 20027 7735
rect 57529 7701 57563 7735
rect 58081 7701 58115 7735
rect 9873 7497 9907 7531
rect 9413 7429 9447 7463
rect 19349 7429 19383 7463
rect 20545 7429 20579 7463
rect 20637 7429 20671 7463
rect 57897 7361 57931 7395
rect 19441 7293 19475 7327
rect 19533 7293 19567 7327
rect 20729 7293 20763 7327
rect 9781 7225 9815 7259
rect 20177 7225 20211 7259
rect 18981 7157 19015 7191
rect 57437 7157 57471 7191
rect 58081 7157 58115 7191
rect 16681 6817 16715 6851
rect 18061 6817 18095 6851
rect 16405 6749 16439 6783
rect 17877 6749 17911 6783
rect 19625 6749 19659 6783
rect 57897 6749 57931 6783
rect 16037 6613 16071 6647
rect 16497 6613 16531 6647
rect 17509 6613 17543 6647
rect 17969 6613 18003 6647
rect 19809 6613 19843 6647
rect 58081 6613 58115 6647
rect 15577 6409 15611 6443
rect 18429 6409 18463 6443
rect 16681 6273 16715 6307
rect 17417 6273 17451 6307
rect 18245 6273 18279 6307
rect 57897 6273 57931 6307
rect 15669 6205 15703 6239
rect 15853 6205 15887 6239
rect 15209 6137 15243 6171
rect 16865 6137 16899 6171
rect 17601 6137 17635 6171
rect 58081 6069 58115 6103
rect 56977 5865 57011 5899
rect 57989 5797 58023 5831
rect 56885 5593 56919 5627
rect 57805 5593 57839 5627
rect 56977 5185 57011 5219
rect 57069 4981 57103 5015
rect 57621 4641 57655 4675
rect 57345 4573 57379 4607
rect 56517 4505 56551 4539
rect 56609 4437 56643 4471
rect 56057 4165 56091 4199
rect 56977 4165 57011 4199
rect 3249 4097 3283 4131
rect 4537 4097 4571 4131
rect 6653 4097 6687 4131
rect 7941 4097 7975 4131
rect 2973 4029 3007 4063
rect 4261 4029 4295 4063
rect 6377 4029 6411 4063
rect 7665 4029 7699 4063
rect 56241 3961 56275 3995
rect 57069 3893 57103 3927
rect 4261 3689 4295 3723
rect 56609 3689 56643 3723
rect 4077 3621 4111 3655
rect 7205 3621 7239 3655
rect 55781 3621 55815 3655
rect 5089 3553 5123 3587
rect 57345 3553 57379 3587
rect 3249 3485 3283 3519
rect 4813 3485 4847 3519
rect 6377 3485 6411 3519
rect 7941 3485 7975 3519
rect 9321 3485 9355 3519
rect 10885 3485 10919 3519
rect 11529 3485 11563 3519
rect 57621 3485 57655 3519
rect 3801 3417 3835 3451
rect 6837 3417 6871 3451
rect 55597 3417 55631 3451
rect 56517 3417 56551 3451
rect 3065 3349 3099 3383
rect 6193 3349 6227 3383
rect 7297 3349 7331 3383
rect 7757 3349 7791 3383
rect 9137 3349 9171 3383
rect 10701 3349 10735 3383
rect 11345 3349 11379 3383
rect 3985 3145 4019 3179
rect 4997 3145 5031 3179
rect 6837 3145 6871 3179
rect 7665 3145 7699 3179
rect 10885 3145 10919 3179
rect 13553 3145 13587 3179
rect 55689 3145 55723 3179
rect 3525 3077 3559 3111
rect 4537 3077 4571 3111
rect 6377 3077 6411 3111
rect 10057 3077 10091 3111
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 5641 3009 5675 3043
rect 7481 3009 7515 3043
rect 8309 3009 8343 3043
rect 9229 3009 9263 3043
rect 9873 3009 9907 3043
rect 10701 3009 10735 3043
rect 11805 3009 11839 3043
rect 12265 3009 12299 3043
rect 13093 3009 13127 3043
rect 13277 3009 13311 3043
rect 13921 3009 13955 3043
rect 49525 3009 49559 3043
rect 53849 3009 53883 3043
rect 55597 3009 55631 3043
rect 56701 3009 56735 3043
rect 7297 2941 7331 2975
rect 9689 2941 9723 2975
rect 10517 2941 10551 2975
rect 12081 2941 12115 2975
rect 12909 2941 12943 2975
rect 49249 2941 49283 2975
rect 53573 2941 53607 2975
rect 56425 2941 56459 2975
rect 2145 2873 2179 2907
rect 3893 2873 3927 2907
rect 4905 2873 4939 2907
rect 6745 2873 6779 2907
rect 8125 2873 8159 2907
rect 2973 2805 3007 2839
rect 5457 2805 5491 2839
rect 9045 2805 9079 2839
rect 12449 2805 12483 2839
rect 13737 2805 13771 2839
rect 3249 2601 3283 2635
rect 4169 2601 4203 2635
rect 5089 2601 5123 2635
rect 16681 2601 16715 2635
rect 17877 2601 17911 2635
rect 19257 2601 19291 2635
rect 20729 2601 20763 2635
rect 22109 2601 22143 2635
rect 23581 2601 23615 2635
rect 24961 2601 24995 2635
rect 26985 2601 27019 2635
rect 27813 2601 27847 2635
rect 29561 2601 29595 2635
rect 30757 2601 30791 2635
rect 32137 2601 32171 2635
rect 33609 2601 33643 2635
rect 34989 2601 35023 2635
rect 36461 2601 36495 2635
rect 37841 2601 37875 2635
rect 39865 2601 39899 2635
rect 40693 2601 40727 2635
rect 42441 2601 42475 2635
rect 43545 2601 43579 2635
rect 45017 2601 45051 2635
rect 46397 2601 46431 2635
rect 57069 2601 57103 2635
rect 7389 2533 7423 2567
rect 10609 2533 10643 2567
rect 13001 2533 13035 2567
rect 15025 2533 15059 2567
rect 6745 2465 6779 2499
rect 9597 2465 9631 2499
rect 9965 2465 9999 2499
rect 48145 2465 48179 2499
rect 50997 2465 51031 2499
rect 53021 2465 53055 2499
rect 55597 2465 55631 2499
rect 1409 2397 1443 2431
rect 2145 2397 2179 2431
rect 2973 2397 3007 2431
rect 3065 2397 3099 2431
rect 3893 2397 3927 2431
rect 3985 2397 4019 2431
rect 4813 2397 4847 2431
rect 4905 2397 4939 2431
rect 5549 2397 5583 2431
rect 6469 2397 6503 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 7941 2397 7975 2431
rect 9137 2397 9171 2431
rect 9781 2397 9815 2431
rect 10425 2397 10459 2431
rect 11529 2397 11563 2431
rect 12265 2397 12299 2431
rect 13185 2397 13219 2431
rect 14105 2397 14139 2431
rect 15209 2397 15243 2431
rect 16865 2397 16899 2431
rect 18061 2397 18095 2431
rect 19441 2397 19475 2431
rect 20913 2397 20947 2431
rect 22293 2397 22327 2431
rect 23765 2397 23799 2431
rect 25145 2397 25179 2431
rect 27169 2397 27203 2431
rect 27997 2397 28031 2431
rect 29745 2397 29779 2431
rect 30941 2397 30975 2431
rect 32321 2397 32355 2431
rect 33793 2397 33827 2431
rect 35173 2397 35207 2431
rect 36645 2397 36679 2431
rect 38025 2397 38059 2431
rect 40049 2397 40083 2431
rect 40877 2397 40911 2431
rect 42625 2397 42659 2431
rect 43729 2397 43763 2431
rect 45201 2397 45235 2431
rect 46581 2397 46615 2431
rect 47869 2397 47903 2431
rect 50721 2397 50755 2431
rect 52745 2397 52779 2431
rect 55321 2397 55355 2431
rect 54401 2329 54435 2363
rect 56977 2329 57011 2363
rect 1593 2261 1627 2295
rect 2329 2261 2363 2295
rect 5733 2261 5767 2295
rect 8125 2261 8159 2295
rect 8953 2261 8987 2295
rect 11713 2261 11747 2295
rect 12449 2261 12483 2295
rect 14289 2261 14323 2295
rect 54493 2261 54527 2295
<< metal1 >>
rect 53006 19796 53012 19848
rect 53064 19836 53070 19848
rect 57146 19836 57152 19848
rect 53064 19808 57152 19836
rect 53064 19796 53070 19808
rect 57146 19796 57152 19808
rect 57204 19796 57210 19848
rect 53374 19728 53380 19780
rect 53432 19768 53438 19780
rect 56962 19768 56968 19780
rect 53432 19740 56968 19768
rect 53432 19728 53438 19740
rect 56962 19728 56968 19740
rect 57020 19728 57026 19780
rect 53926 19660 53932 19712
rect 53984 19700 53990 19712
rect 57054 19700 57060 19712
rect 53984 19672 57060 19700
rect 53984 19660 53990 19672
rect 57054 19660 57060 19672
rect 57112 19660 57118 19712
rect 1104 19610 58880 19632
rect 1104 19558 20214 19610
rect 20266 19558 20278 19610
rect 20330 19558 20342 19610
rect 20394 19558 20406 19610
rect 20458 19558 20470 19610
rect 20522 19558 39478 19610
rect 39530 19558 39542 19610
rect 39594 19558 39606 19610
rect 39658 19558 39670 19610
rect 39722 19558 39734 19610
rect 39786 19558 58880 19610
rect 1104 19536 58880 19558
rect 1026 19456 1032 19508
rect 1084 19496 1090 19508
rect 1581 19499 1639 19505
rect 1581 19496 1593 19499
rect 1084 19468 1593 19496
rect 1084 19456 1090 19468
rect 1581 19465 1593 19468
rect 1627 19465 1639 19499
rect 2314 19496 2320 19508
rect 2275 19468 2320 19496
rect 1581 19459 1639 19465
rect 2314 19456 2320 19468
rect 2372 19456 2378 19508
rect 3510 19456 3516 19508
rect 3568 19496 3574 19508
rect 3973 19499 4031 19505
rect 3973 19496 3985 19499
rect 3568 19468 3985 19496
rect 3568 19456 3574 19468
rect 3973 19465 3985 19468
rect 4019 19465 4031 19499
rect 5166 19496 5172 19508
rect 5127 19468 5172 19496
rect 3973 19459 4031 19465
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 6638 19496 6644 19508
rect 6599 19468 6644 19496
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 8018 19496 8024 19508
rect 7979 19468 8024 19496
rect 8018 19456 8024 19468
rect 8076 19456 8082 19508
rect 9490 19496 9496 19508
rect 9451 19468 9496 19496
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 10870 19496 10876 19508
rect 10831 19468 10876 19496
rect 10870 19456 10876 19468
rect 10928 19456 10934 19508
rect 12342 19496 12348 19508
rect 12303 19468 12348 19496
rect 12342 19456 12348 19468
rect 12400 19456 12406 19508
rect 13446 19456 13452 19508
rect 13504 19496 13510 19508
rect 14277 19499 14335 19505
rect 14277 19496 14289 19499
rect 13504 19468 14289 19496
rect 13504 19456 13510 19468
rect 14277 19465 14289 19468
rect 14323 19465 14335 19499
rect 14277 19459 14335 19465
rect 16390 19456 16396 19508
rect 16448 19496 16454 19508
rect 16669 19499 16727 19505
rect 16669 19496 16681 19499
rect 16448 19468 16681 19496
rect 16448 19456 16454 19468
rect 16669 19465 16681 19468
rect 16715 19465 16727 19499
rect 16669 19459 16727 19465
rect 20070 19456 20076 19508
rect 20128 19496 20134 19508
rect 20717 19499 20775 19505
rect 20717 19496 20729 19499
rect 20128 19468 20729 19496
rect 20128 19456 20134 19468
rect 20717 19465 20729 19468
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 22097 19499 22155 19505
rect 22097 19465 22109 19499
rect 22143 19496 22155 19499
rect 22554 19496 22560 19508
rect 22143 19468 22560 19496
rect 22143 19465 22155 19468
rect 22097 19459 22155 19465
rect 22554 19456 22560 19468
rect 22612 19456 22618 19508
rect 26973 19499 27031 19505
rect 26973 19465 26985 19499
rect 27019 19496 27031 19499
rect 27338 19496 27344 19508
rect 27019 19468 27344 19496
rect 27019 19465 27031 19468
rect 26973 19459 27031 19465
rect 27338 19456 27344 19468
rect 27396 19456 27402 19508
rect 29549 19499 29607 19505
rect 29549 19465 29561 19499
rect 29595 19496 29607 19499
rect 29638 19496 29644 19508
rect 29595 19468 29644 19496
rect 29595 19465 29607 19468
rect 29549 19459 29607 19465
rect 29638 19456 29644 19468
rect 29696 19456 29702 19508
rect 30745 19499 30803 19505
rect 30745 19465 30757 19499
rect 30791 19496 30803 19499
rect 31018 19496 31024 19508
rect 30791 19468 31024 19496
rect 30791 19465 30803 19468
rect 30745 19459 30803 19465
rect 31018 19456 31024 19468
rect 31076 19456 31082 19508
rect 32125 19499 32183 19505
rect 32125 19465 32137 19499
rect 32171 19496 32183 19499
rect 32490 19496 32496 19508
rect 32171 19468 32496 19496
rect 32171 19465 32183 19468
rect 32125 19459 32183 19465
rect 32490 19456 32496 19468
rect 32548 19456 32554 19508
rect 33597 19499 33655 19505
rect 33597 19465 33609 19499
rect 33643 19496 33655 19499
rect 33686 19496 33692 19508
rect 33643 19468 33692 19496
rect 33643 19465 33655 19468
rect 33597 19459 33655 19465
rect 33686 19456 33692 19468
rect 33744 19456 33750 19508
rect 34977 19499 35035 19505
rect 34977 19465 34989 19499
rect 35023 19496 35035 19499
rect 35066 19496 35072 19508
rect 35023 19468 35072 19496
rect 35023 19465 35035 19468
rect 34977 19459 35035 19465
rect 35066 19456 35072 19468
rect 35124 19456 35130 19508
rect 39298 19456 39304 19508
rect 39356 19496 39362 19508
rect 39853 19499 39911 19505
rect 39853 19496 39865 19499
rect 39356 19468 39865 19496
rect 39356 19456 39362 19468
rect 39853 19465 39865 19468
rect 39899 19465 39911 19499
rect 39853 19459 39911 19465
rect 40681 19499 40739 19505
rect 40681 19465 40693 19499
rect 40727 19496 40739 19499
rect 41506 19496 41512 19508
rect 40727 19468 41512 19496
rect 40727 19465 40739 19468
rect 40681 19459 40739 19465
rect 41506 19456 41512 19468
rect 41564 19456 41570 19508
rect 41874 19456 41880 19508
rect 41932 19496 41938 19508
rect 42429 19499 42487 19505
rect 42429 19496 42441 19499
rect 41932 19468 42441 19496
rect 41932 19456 41938 19468
rect 42429 19465 42441 19468
rect 42475 19465 42487 19499
rect 42429 19459 42487 19465
rect 43533 19499 43591 19505
rect 43533 19465 43545 19499
rect 43579 19496 43591 19499
rect 43990 19496 43996 19508
rect 43579 19468 43996 19496
rect 43579 19465 43591 19468
rect 43533 19459 43591 19465
rect 43990 19456 43996 19468
rect 44048 19456 44054 19508
rect 45005 19499 45063 19505
rect 45005 19465 45017 19499
rect 45051 19496 45063 19499
rect 45370 19496 45376 19508
rect 45051 19468 45376 19496
rect 45051 19465 45063 19468
rect 45005 19459 45063 19465
rect 45370 19456 45376 19468
rect 45428 19456 45434 19508
rect 48958 19456 48964 19508
rect 49016 19496 49022 19508
rect 49237 19499 49295 19505
rect 49237 19496 49249 19499
rect 49016 19468 49249 19496
rect 49016 19456 49022 19468
rect 49237 19465 49249 19468
rect 49283 19465 49295 19499
rect 49237 19459 49295 19465
rect 50709 19499 50767 19505
rect 50709 19465 50721 19499
rect 50755 19496 50767 19499
rect 51166 19496 51172 19508
rect 50755 19468 51172 19496
rect 50755 19465 50767 19468
rect 50709 19459 50767 19465
rect 51166 19456 51172 19468
rect 51224 19456 51230 19508
rect 53193 19499 53251 19505
rect 53193 19465 53205 19499
rect 53239 19465 53251 19499
rect 53193 19459 53251 19465
rect 53837 19499 53895 19505
rect 53837 19465 53849 19499
rect 53883 19496 53895 19499
rect 54665 19499 54723 19505
rect 53883 19468 54616 19496
rect 53883 19465 53895 19468
rect 53837 19459 53895 19465
rect 53208 19428 53236 19459
rect 54588 19428 54616 19468
rect 54665 19465 54677 19499
rect 54711 19496 54723 19499
rect 56226 19496 56232 19508
rect 54711 19468 56232 19496
rect 54711 19465 54723 19468
rect 54665 19459 54723 19465
rect 56226 19456 56232 19468
rect 56284 19456 56290 19508
rect 56502 19496 56508 19508
rect 56463 19468 56508 19496
rect 56502 19456 56508 19468
rect 56560 19456 56566 19508
rect 57882 19456 57888 19508
rect 57940 19496 57946 19508
rect 58069 19499 58127 19505
rect 58069 19496 58081 19499
rect 57940 19468 58081 19496
rect 57940 19456 57946 19468
rect 58069 19465 58081 19468
rect 58115 19465 58127 19499
rect 58069 19459 58127 19465
rect 53208 19400 54524 19428
rect 54588 19400 56364 19428
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19320 1458 19372
rect 2130 19360 2136 19372
rect 2091 19332 2136 19360
rect 2130 19320 2136 19332
rect 2188 19320 2194 19372
rect 3786 19360 3792 19372
rect 3747 19332 3792 19360
rect 3786 19320 3792 19332
rect 3844 19320 3850 19372
rect 4985 19363 5043 19369
rect 4985 19329 4997 19363
rect 5031 19360 5043 19363
rect 5074 19360 5080 19372
rect 5031 19332 5080 19360
rect 5031 19329 5043 19332
rect 4985 19323 5043 19329
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 6457 19363 6515 19369
rect 6457 19329 6469 19363
rect 6503 19360 6515 19363
rect 6546 19360 6552 19372
rect 6503 19332 6552 19360
rect 6503 19329 6515 19332
rect 6457 19323 6515 19329
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19360 7895 19363
rect 7926 19360 7932 19372
rect 7883 19332 7932 19360
rect 7883 19329 7895 19332
rect 7837 19323 7895 19329
rect 7926 19320 7932 19332
rect 7984 19320 7990 19372
rect 9309 19363 9367 19369
rect 9309 19329 9321 19363
rect 9355 19360 9367 19363
rect 9398 19360 9404 19372
rect 9355 19332 9404 19360
rect 9355 19329 9367 19332
rect 9309 19323 9367 19329
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 10502 19320 10508 19372
rect 10560 19360 10566 19372
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 10560 19332 10701 19360
rect 10560 19320 10566 19332
rect 10689 19329 10701 19332
rect 10735 19329 10747 19363
rect 10689 19323 10747 19329
rect 12066 19320 12072 19372
rect 12124 19360 12130 19372
rect 12161 19363 12219 19369
rect 12161 19360 12173 19363
rect 12124 19332 12173 19360
rect 12124 19320 12130 19332
rect 12161 19329 12173 19332
rect 12207 19329 12219 19363
rect 14090 19360 14096 19372
rect 14051 19332 14096 19360
rect 12161 19323 12219 19329
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 14918 19320 14924 19372
rect 14976 19360 14982 19372
rect 15197 19363 15255 19369
rect 15197 19360 15209 19363
rect 14976 19332 15209 19360
rect 14976 19320 14982 19332
rect 15197 19329 15209 19332
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 16298 19320 16304 19372
rect 16356 19360 16362 19372
rect 16853 19363 16911 19369
rect 16853 19360 16865 19363
rect 16356 19332 16865 19360
rect 16356 19320 16362 19332
rect 16853 19329 16865 19332
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 18049 19363 18107 19369
rect 18049 19360 18061 19363
rect 17828 19332 18061 19360
rect 17828 19320 17834 19332
rect 18049 19329 18061 19332
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 19150 19320 19156 19372
rect 19208 19360 19214 19372
rect 19429 19363 19487 19369
rect 19429 19360 19441 19363
rect 19208 19332 19441 19360
rect 19208 19320 19214 19332
rect 19429 19329 19441 19332
rect 19475 19329 19487 19363
rect 19429 19323 19487 19329
rect 20622 19320 20628 19372
rect 20680 19360 20686 19372
rect 20901 19363 20959 19369
rect 20901 19360 20913 19363
rect 20680 19332 20913 19360
rect 20680 19320 20686 19332
rect 20901 19329 20913 19332
rect 20947 19329 20959 19363
rect 20901 19323 20959 19329
rect 22002 19320 22008 19372
rect 22060 19360 22066 19372
rect 22281 19363 22339 19369
rect 22281 19360 22293 19363
rect 22060 19332 22293 19360
rect 22060 19320 22066 19332
rect 22281 19329 22293 19332
rect 22327 19329 22339 19363
rect 23750 19360 23756 19372
rect 23711 19332 23756 19360
rect 22281 19323 22339 19329
rect 23750 19320 23756 19332
rect 23808 19320 23814 19372
rect 25130 19360 25136 19372
rect 25091 19332 25136 19360
rect 25130 19320 25136 19332
rect 25188 19320 25194 19372
rect 26326 19320 26332 19372
rect 26384 19360 26390 19372
rect 27157 19363 27215 19369
rect 27157 19360 27169 19363
rect 26384 19332 27169 19360
rect 26384 19320 26390 19332
rect 27157 19329 27169 19332
rect 27203 19329 27215 19363
rect 27982 19360 27988 19372
rect 27943 19332 27988 19360
rect 27157 19323 27215 19329
rect 27982 19320 27988 19332
rect 28040 19320 28046 19372
rect 29178 19320 29184 19372
rect 29236 19360 29242 19372
rect 29733 19363 29791 19369
rect 29733 19360 29745 19363
rect 29236 19332 29745 19360
rect 29236 19320 29242 19332
rect 29733 19329 29745 19332
rect 29779 19329 29791 19363
rect 30926 19360 30932 19372
rect 30887 19332 30932 19360
rect 29733 19323 29791 19329
rect 30926 19320 30932 19332
rect 30984 19320 30990 19372
rect 32306 19360 32312 19372
rect 32267 19332 32312 19360
rect 32306 19320 32312 19332
rect 32364 19320 32370 19372
rect 33778 19360 33784 19372
rect 33739 19332 33784 19360
rect 33778 19320 33784 19332
rect 33836 19320 33842 19372
rect 35158 19360 35164 19372
rect 35119 19332 35164 19360
rect 35158 19320 35164 19332
rect 35216 19320 35222 19372
rect 36630 19360 36636 19372
rect 36591 19332 36636 19360
rect 36630 19320 36636 19332
rect 36688 19320 36694 19372
rect 38010 19360 38016 19372
rect 37971 19332 38016 19360
rect 38010 19320 38016 19332
rect 38068 19320 38074 19372
rect 39206 19320 39212 19372
rect 39264 19360 39270 19372
rect 40037 19363 40095 19369
rect 40037 19360 40049 19363
rect 39264 19332 40049 19360
rect 39264 19320 39270 19332
rect 40037 19329 40049 19332
rect 40083 19329 40095 19363
rect 40862 19360 40868 19372
rect 40823 19332 40868 19360
rect 40037 19323 40095 19329
rect 40862 19320 40868 19332
rect 40920 19320 40926 19372
rect 42058 19320 42064 19372
rect 42116 19360 42122 19372
rect 42613 19363 42671 19369
rect 42613 19360 42625 19363
rect 42116 19332 42625 19360
rect 42116 19320 42122 19332
rect 42613 19329 42625 19332
rect 42659 19329 42671 19363
rect 43714 19360 43720 19372
rect 43675 19332 43720 19360
rect 42613 19323 42671 19329
rect 43714 19320 43720 19332
rect 43772 19320 43778 19372
rect 44910 19320 44916 19372
rect 44968 19360 44974 19372
rect 45189 19363 45247 19369
rect 45189 19360 45201 19363
rect 44968 19332 45201 19360
rect 44968 19320 44974 19332
rect 45189 19329 45201 19332
rect 45235 19329 45247 19363
rect 46566 19360 46572 19372
rect 46527 19332 46572 19360
rect 45189 19323 45247 19329
rect 46566 19320 46572 19332
rect 46624 19320 46630 19372
rect 48038 19360 48044 19372
rect 47999 19332 48044 19360
rect 48038 19320 48044 19332
rect 48096 19320 48102 19372
rect 49418 19360 49424 19372
rect 49379 19332 49424 19360
rect 49418 19320 49424 19332
rect 49476 19320 49482 19372
rect 50890 19360 50896 19372
rect 50851 19332 50896 19360
rect 50890 19320 50896 19332
rect 50948 19320 50954 19372
rect 52178 19360 52184 19372
rect 52139 19332 52184 19360
rect 52178 19320 52184 19332
rect 52236 19320 52242 19372
rect 53374 19360 53380 19372
rect 53335 19332 53380 19360
rect 53374 19320 53380 19332
rect 53432 19320 53438 19372
rect 54018 19360 54024 19372
rect 53979 19332 54024 19360
rect 54018 19320 54024 19332
rect 54076 19320 54082 19372
rect 54496 19369 54524 19400
rect 54481 19363 54539 19369
rect 54481 19329 54493 19363
rect 54527 19329 54539 19363
rect 55582 19360 55588 19372
rect 55543 19332 55588 19360
rect 54481 19323 54539 19329
rect 55582 19320 55588 19332
rect 55640 19320 55646 19372
rect 55766 19320 55772 19372
rect 55824 19320 55830 19372
rect 56336 19369 56364 19400
rect 56321 19363 56379 19369
rect 56321 19329 56333 19363
rect 56367 19329 56379 19363
rect 57054 19360 57060 19372
rect 57015 19332 57060 19360
rect 56321 19323 56379 19329
rect 57054 19320 57060 19332
rect 57112 19320 57118 19372
rect 57146 19320 57152 19372
rect 57204 19360 57210 19372
rect 57885 19363 57943 19369
rect 57885 19360 57897 19363
rect 57204 19332 57897 19360
rect 57204 19320 57210 19332
rect 57885 19329 57897 19332
rect 57931 19329 57943 19363
rect 57885 19323 57943 19329
rect 55784 19233 55812 19320
rect 55769 19227 55827 19233
rect 55769 19193 55781 19227
rect 55815 19193 55827 19227
rect 55769 19187 55827 19193
rect 15010 19156 15016 19168
rect 14971 19128 15016 19156
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 17862 19156 17868 19168
rect 17823 19128 17868 19156
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 19242 19156 19248 19168
rect 19203 19128 19248 19156
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 23566 19156 23572 19168
rect 23527 19128 23572 19156
rect 23566 19116 23572 19128
rect 23624 19116 23630 19168
rect 24946 19156 24952 19168
rect 24907 19128 24952 19156
rect 24946 19116 24952 19128
rect 25004 19116 25010 19168
rect 27798 19156 27804 19168
rect 27759 19128 27804 19156
rect 27798 19116 27804 19128
rect 27856 19116 27862 19168
rect 36446 19156 36452 19168
rect 36407 19128 36452 19156
rect 36446 19116 36452 19128
rect 36504 19116 36510 19168
rect 37826 19156 37832 19168
rect 37787 19128 37832 19156
rect 37826 19116 37832 19128
rect 37884 19116 37890 19168
rect 46382 19156 46388 19168
rect 46343 19128 46388 19156
rect 46382 19116 46388 19128
rect 46440 19116 46446 19168
rect 47854 19156 47860 19168
rect 47815 19128 47860 19156
rect 47854 19116 47860 19128
rect 47912 19116 47918 19168
rect 51997 19159 52055 19165
rect 51997 19125 52009 19159
rect 52043 19156 52055 19159
rect 52270 19156 52276 19168
rect 52043 19128 52276 19156
rect 52043 19125 52055 19128
rect 51997 19119 52055 19125
rect 52270 19116 52276 19128
rect 52328 19116 52334 19168
rect 57238 19156 57244 19168
rect 57199 19128 57244 19156
rect 57238 19116 57244 19128
rect 57296 19116 57302 19168
rect 1104 19066 58880 19088
rect 1104 19014 10582 19066
rect 10634 19014 10646 19066
rect 10698 19014 10710 19066
rect 10762 19014 10774 19066
rect 10826 19014 10838 19066
rect 10890 19014 29846 19066
rect 29898 19014 29910 19066
rect 29962 19014 29974 19066
rect 30026 19014 30038 19066
rect 30090 19014 30102 19066
rect 30154 19014 49110 19066
rect 49162 19014 49174 19066
rect 49226 19014 49238 19066
rect 49290 19014 49302 19066
rect 49354 19014 49366 19066
rect 49418 19014 58880 19066
rect 1104 18992 58880 19014
rect 53193 18955 53251 18961
rect 53193 18921 53205 18955
rect 53239 18952 53251 18955
rect 54018 18952 54024 18964
rect 53239 18924 54024 18952
rect 53239 18921 53251 18924
rect 53193 18915 53251 18921
rect 54018 18912 54024 18924
rect 54076 18912 54082 18964
rect 54573 18955 54631 18961
rect 54573 18921 54585 18955
rect 54619 18952 54631 18955
rect 55582 18952 55588 18964
rect 54619 18924 55588 18952
rect 54619 18921 54631 18924
rect 54573 18915 54631 18921
rect 55582 18912 55588 18924
rect 55640 18912 55646 18964
rect 51074 18844 51080 18896
rect 51132 18884 51138 18896
rect 51132 18856 57928 18884
rect 51132 18844 51138 18856
rect 51445 18819 51503 18825
rect 51445 18785 51457 18819
rect 51491 18816 51503 18819
rect 52641 18819 52699 18825
rect 52641 18816 52653 18819
rect 51491 18788 52653 18816
rect 51491 18785 51503 18788
rect 51445 18779 51503 18785
rect 52641 18785 52653 18788
rect 52687 18816 52699 18819
rect 53745 18819 53803 18825
rect 53745 18816 53757 18819
rect 52687 18788 53757 18816
rect 52687 18785 52699 18788
rect 52641 18779 52699 18785
rect 53745 18785 53757 18788
rect 53791 18816 53803 18819
rect 55858 18816 55864 18828
rect 53791 18788 55864 18816
rect 53791 18785 53803 18788
rect 53745 18779 53803 18785
rect 55858 18776 55864 18788
rect 55916 18816 55922 18828
rect 55953 18819 56011 18825
rect 55953 18816 55965 18819
rect 55916 18788 55965 18816
rect 55916 18776 55922 18788
rect 55953 18785 55965 18788
rect 55999 18816 56011 18819
rect 57057 18819 57115 18825
rect 57057 18816 57069 18819
rect 55999 18788 57069 18816
rect 55999 18785 56011 18788
rect 55953 18779 56011 18785
rect 57057 18785 57069 18788
rect 57103 18785 57115 18819
rect 57057 18779 57115 18785
rect 51166 18748 51172 18760
rect 51127 18720 51172 18748
rect 51166 18708 51172 18720
rect 51224 18708 51230 18760
rect 52362 18708 52368 18760
rect 52420 18748 52426 18760
rect 57900 18757 57928 18856
rect 52457 18751 52515 18757
rect 52457 18748 52469 18751
rect 52420 18720 52469 18748
rect 52420 18708 52426 18720
rect 52457 18717 52469 18720
rect 52503 18717 52515 18751
rect 52457 18711 52515 18717
rect 54757 18751 54815 18757
rect 54757 18717 54769 18751
rect 54803 18748 54815 18751
rect 57885 18751 57943 18757
rect 54803 18720 55214 18748
rect 54803 18717 54815 18720
rect 54757 18711 54815 18717
rect 50798 18612 50804 18624
rect 50759 18584 50804 18612
rect 50798 18572 50804 18584
rect 50856 18572 50862 18624
rect 50982 18572 50988 18624
rect 51040 18612 51046 18624
rect 51261 18615 51319 18621
rect 51261 18612 51273 18615
rect 51040 18584 51273 18612
rect 51040 18572 51046 18584
rect 51261 18581 51273 18584
rect 51307 18581 51319 18615
rect 51994 18612 52000 18624
rect 51955 18584 52000 18612
rect 51261 18575 51319 18581
rect 51994 18572 52000 18584
rect 52052 18572 52058 18624
rect 52270 18572 52276 18624
rect 52328 18612 52334 18624
rect 52365 18615 52423 18621
rect 52365 18612 52377 18615
rect 52328 18584 52377 18612
rect 52328 18572 52334 18584
rect 52365 18581 52377 18584
rect 52411 18581 52423 18615
rect 53558 18612 53564 18624
rect 53519 18584 53564 18612
rect 52365 18575 52423 18581
rect 53558 18572 53564 18584
rect 53616 18572 53622 18624
rect 53653 18615 53711 18621
rect 53653 18581 53665 18615
rect 53699 18612 53711 18615
rect 53834 18612 53840 18624
rect 53699 18584 53840 18612
rect 53699 18581 53711 18584
rect 53653 18575 53711 18581
rect 53834 18572 53840 18584
rect 53892 18572 53898 18624
rect 55186 18612 55214 18720
rect 57885 18717 57897 18751
rect 57931 18717 57943 18751
rect 57885 18711 57943 18717
rect 55490 18640 55496 18692
rect 55548 18680 55554 18692
rect 55769 18683 55827 18689
rect 55769 18680 55781 18683
rect 55548 18652 55781 18680
rect 55548 18640 55554 18652
rect 55769 18649 55781 18652
rect 55815 18649 55827 18683
rect 55769 18643 55827 18649
rect 56686 18640 56692 18692
rect 56744 18680 56750 18692
rect 56965 18683 57023 18689
rect 56965 18680 56977 18683
rect 56744 18652 56977 18680
rect 56744 18640 56750 18652
rect 56965 18649 56977 18652
rect 57011 18649 57023 18683
rect 56965 18643 57023 18649
rect 55309 18615 55367 18621
rect 55309 18612 55321 18615
rect 55186 18584 55321 18612
rect 55309 18581 55321 18584
rect 55355 18581 55367 18615
rect 55674 18612 55680 18624
rect 55635 18584 55680 18612
rect 55309 18575 55367 18581
rect 55674 18572 55680 18584
rect 55732 18572 55738 18624
rect 56502 18612 56508 18624
rect 56463 18584 56508 18612
rect 56502 18572 56508 18584
rect 56560 18572 56566 18624
rect 56870 18612 56876 18624
rect 56831 18584 56876 18612
rect 56870 18572 56876 18584
rect 56928 18572 56934 18624
rect 58066 18612 58072 18624
rect 58027 18584 58072 18612
rect 58066 18572 58072 18584
rect 58124 18572 58130 18624
rect 1104 18522 58880 18544
rect 1104 18470 20214 18522
rect 20266 18470 20278 18522
rect 20330 18470 20342 18522
rect 20394 18470 20406 18522
rect 20458 18470 20470 18522
rect 20522 18470 39478 18522
rect 39530 18470 39542 18522
rect 39594 18470 39606 18522
rect 39658 18470 39670 18522
rect 39722 18470 39734 18522
rect 39786 18470 58880 18522
rect 1104 18448 58880 18470
rect 51537 18411 51595 18417
rect 51537 18377 51549 18411
rect 51583 18408 51595 18411
rect 53006 18408 53012 18420
rect 51583 18380 53012 18408
rect 51583 18377 51595 18380
rect 51537 18371 51595 18377
rect 53006 18368 53012 18380
rect 53064 18368 53070 18420
rect 53558 18408 53564 18420
rect 53519 18380 53564 18408
rect 53558 18368 53564 18380
rect 53616 18368 53622 18420
rect 54573 18411 54631 18417
rect 54573 18377 54585 18411
rect 54619 18408 54631 18411
rect 55674 18408 55680 18420
rect 54619 18380 55680 18408
rect 54619 18377 54631 18380
rect 54573 18371 54631 18377
rect 55674 18368 55680 18380
rect 55732 18368 55738 18420
rect 56042 18408 56048 18420
rect 56003 18380 56048 18408
rect 56042 18368 56048 18380
rect 56100 18368 56106 18420
rect 56502 18340 56508 18352
rect 55416 18312 56508 18340
rect 50798 18232 50804 18284
rect 50856 18272 50862 18284
rect 51721 18275 51779 18281
rect 51721 18272 51733 18275
rect 50856 18244 51733 18272
rect 50856 18232 50862 18244
rect 51721 18241 51733 18244
rect 51767 18241 51779 18275
rect 51721 18235 51779 18241
rect 51994 18232 52000 18284
rect 52052 18272 52058 18284
rect 52917 18275 52975 18281
rect 52917 18272 52929 18275
rect 52052 18244 52929 18272
rect 52052 18232 52058 18244
rect 52917 18241 52929 18244
rect 52963 18241 52975 18275
rect 53742 18272 53748 18284
rect 53703 18244 53748 18272
rect 52917 18235 52975 18241
rect 53742 18232 53748 18244
rect 53800 18232 53806 18284
rect 54754 18272 54760 18284
rect 54715 18244 54760 18272
rect 54754 18232 54760 18244
rect 54812 18232 54818 18284
rect 55416 18281 55444 18312
rect 56502 18300 56508 18312
rect 56560 18300 56566 18352
rect 57057 18343 57115 18349
rect 57057 18309 57069 18343
rect 57103 18340 57115 18343
rect 57698 18340 57704 18352
rect 57103 18312 57704 18340
rect 57103 18309 57115 18312
rect 57057 18303 57115 18309
rect 57698 18300 57704 18312
rect 57756 18300 57762 18352
rect 55401 18275 55459 18281
rect 55401 18241 55413 18275
rect 55447 18241 55459 18275
rect 55401 18235 55459 18241
rect 55861 18275 55919 18281
rect 55861 18241 55873 18275
rect 55907 18241 55919 18275
rect 55861 18235 55919 18241
rect 55876 18204 55904 18235
rect 56594 18232 56600 18284
rect 56652 18272 56658 18284
rect 56965 18275 57023 18281
rect 56965 18272 56977 18275
rect 56652 18244 56977 18272
rect 56652 18232 56658 18244
rect 56965 18241 56977 18244
rect 57011 18241 57023 18275
rect 56965 18235 57023 18241
rect 57238 18232 57244 18284
rect 57296 18272 57302 18284
rect 57885 18275 57943 18281
rect 57885 18272 57897 18275
rect 57296 18244 57897 18272
rect 57296 18232 57302 18244
rect 57885 18241 57897 18244
rect 57931 18241 57943 18275
rect 57885 18235 57943 18241
rect 55232 18176 55904 18204
rect 52733 18139 52791 18145
rect 52733 18105 52745 18139
rect 52779 18136 52791 18139
rect 53926 18136 53932 18148
rect 52779 18108 53932 18136
rect 52779 18105 52791 18108
rect 52733 18099 52791 18105
rect 53926 18096 53932 18108
rect 53984 18096 53990 18148
rect 55232 18145 55260 18176
rect 56778 18164 56784 18216
rect 56836 18204 56842 18216
rect 57149 18207 57207 18213
rect 57149 18204 57161 18207
rect 56836 18176 57161 18204
rect 56836 18164 56842 18176
rect 57149 18173 57161 18176
rect 57195 18173 57207 18207
rect 57149 18167 57207 18173
rect 55217 18139 55275 18145
rect 55217 18105 55229 18139
rect 55263 18105 55275 18139
rect 55217 18099 55275 18105
rect 56597 18071 56655 18077
rect 56597 18037 56609 18071
rect 56643 18068 56655 18071
rect 57422 18068 57428 18080
rect 56643 18040 57428 18068
rect 56643 18037 56655 18040
rect 56597 18031 56655 18037
rect 57422 18028 57428 18040
rect 57480 18028 57486 18080
rect 57882 18028 57888 18080
rect 57940 18068 57946 18080
rect 58069 18071 58127 18077
rect 58069 18068 58081 18071
rect 57940 18040 58081 18068
rect 57940 18028 57946 18040
rect 58069 18037 58081 18040
rect 58115 18037 58127 18071
rect 58069 18031 58127 18037
rect 1104 17978 58880 18000
rect 1104 17926 10582 17978
rect 10634 17926 10646 17978
rect 10698 17926 10710 17978
rect 10762 17926 10774 17978
rect 10826 17926 10838 17978
rect 10890 17926 29846 17978
rect 29898 17926 29910 17978
rect 29962 17926 29974 17978
rect 30026 17926 30038 17978
rect 30090 17926 30102 17978
rect 30154 17926 49110 17978
rect 49162 17926 49174 17978
rect 49226 17926 49238 17978
rect 49290 17926 49302 17978
rect 49354 17926 49366 17978
rect 49418 17926 58880 17978
rect 1104 17904 58880 17926
rect 47949 17867 48007 17873
rect 47949 17833 47961 17867
rect 47995 17864 48007 17867
rect 55858 17864 55864 17876
rect 47995 17836 55214 17864
rect 55819 17836 55864 17864
rect 47995 17833 48007 17836
rect 47949 17827 48007 17833
rect 48593 17799 48651 17805
rect 48593 17765 48605 17799
rect 48639 17796 48651 17799
rect 48639 17768 50384 17796
rect 48639 17765 48651 17768
rect 48593 17759 48651 17765
rect 48222 17688 48228 17740
rect 48280 17728 48286 17740
rect 49145 17731 49203 17737
rect 49145 17728 49157 17731
rect 48280 17700 49157 17728
rect 48280 17688 48286 17700
rect 49145 17697 49157 17700
rect 49191 17697 49203 17731
rect 49145 17691 49203 17697
rect 46014 17620 46020 17672
rect 46072 17660 46078 17672
rect 46937 17663 46995 17669
rect 46937 17660 46949 17663
rect 46072 17632 46949 17660
rect 46072 17620 46078 17632
rect 46937 17629 46949 17632
rect 46983 17629 46995 17663
rect 46937 17623 46995 17629
rect 47578 17620 47584 17672
rect 47636 17660 47642 17672
rect 48133 17663 48191 17669
rect 48133 17660 48145 17663
rect 47636 17632 48145 17660
rect 47636 17620 47642 17632
rect 48133 17629 48145 17632
rect 48179 17629 48191 17663
rect 48958 17660 48964 17672
rect 48919 17632 48964 17660
rect 48133 17623 48191 17629
rect 48958 17620 48964 17632
rect 49016 17620 49022 17672
rect 50356 17669 50384 17768
rect 55186 17728 55214 17836
rect 55858 17824 55864 17836
rect 55916 17824 55922 17876
rect 55950 17824 55956 17876
rect 56008 17864 56014 17876
rect 56597 17867 56655 17873
rect 56597 17864 56609 17867
rect 56008 17836 56609 17864
rect 56008 17824 56014 17836
rect 56597 17833 56609 17836
rect 56643 17833 56655 17867
rect 56597 17827 56655 17833
rect 56962 17824 56968 17876
rect 57020 17864 57026 17876
rect 57149 17867 57207 17873
rect 57149 17864 57161 17867
rect 57020 17836 57161 17864
rect 57020 17824 57026 17836
rect 57149 17833 57161 17836
rect 57195 17833 57207 17867
rect 57149 17827 57207 17833
rect 56778 17756 56784 17808
rect 56836 17796 56842 17808
rect 56836 17768 57744 17796
rect 56836 17756 56842 17768
rect 57238 17728 57244 17740
rect 55186 17700 57244 17728
rect 57238 17688 57244 17700
rect 57296 17688 57302 17740
rect 57716 17737 57744 17768
rect 57701 17731 57759 17737
rect 57701 17697 57713 17731
rect 57747 17697 57759 17731
rect 57701 17691 57759 17697
rect 50341 17663 50399 17669
rect 50341 17629 50353 17663
rect 50387 17629 50399 17663
rect 50341 17623 50399 17629
rect 56413 17663 56471 17669
rect 56413 17629 56425 17663
rect 56459 17660 56471 17663
rect 57146 17660 57152 17672
rect 56459 17632 57152 17660
rect 56459 17629 56471 17632
rect 56413 17623 56471 17629
rect 57146 17620 57152 17632
rect 57204 17620 57210 17672
rect 55766 17592 55772 17604
rect 55727 17564 55772 17592
rect 55766 17552 55772 17564
rect 55824 17552 55830 17604
rect 56962 17552 56968 17604
rect 57020 17592 57026 17604
rect 57609 17595 57667 17601
rect 57609 17592 57621 17595
rect 57020 17564 57621 17592
rect 57020 17552 57026 17564
rect 57609 17561 57621 17564
rect 57655 17561 57667 17595
rect 57609 17555 57667 17561
rect 46750 17524 46756 17536
rect 46711 17496 46756 17524
rect 46750 17484 46756 17496
rect 46808 17484 46814 17536
rect 49053 17527 49111 17533
rect 49053 17493 49065 17527
rect 49099 17524 49111 17527
rect 49510 17524 49516 17536
rect 49099 17496 49516 17524
rect 49099 17493 49111 17496
rect 49053 17487 49111 17493
rect 49510 17484 49516 17496
rect 49568 17484 49574 17536
rect 50157 17527 50215 17533
rect 50157 17493 50169 17527
rect 50203 17524 50215 17527
rect 51074 17524 51080 17536
rect 50203 17496 51080 17524
rect 50203 17493 50215 17496
rect 50157 17487 50215 17493
rect 51074 17484 51080 17496
rect 51132 17484 51138 17536
rect 57514 17524 57520 17536
rect 57475 17496 57520 17524
rect 57514 17484 57520 17496
rect 57572 17484 57578 17536
rect 1104 17434 58880 17456
rect 1104 17382 20214 17434
rect 20266 17382 20278 17434
rect 20330 17382 20342 17434
rect 20394 17382 20406 17434
rect 20458 17382 20470 17434
rect 20522 17382 39478 17434
rect 39530 17382 39542 17434
rect 39594 17382 39606 17434
rect 39658 17382 39670 17434
rect 39722 17382 39734 17434
rect 39786 17382 58880 17434
rect 1104 17360 58880 17382
rect 46014 17320 46020 17332
rect 45975 17292 46020 17320
rect 46014 17280 46020 17292
rect 46072 17280 46078 17332
rect 46382 17320 46388 17332
rect 46343 17292 46388 17320
rect 46382 17280 46388 17292
rect 46440 17280 46446 17332
rect 47578 17320 47584 17332
rect 47539 17292 47584 17320
rect 47578 17280 47584 17292
rect 47636 17280 47642 17332
rect 47854 17280 47860 17332
rect 47912 17320 47918 17332
rect 47949 17323 48007 17329
rect 47949 17320 47961 17323
rect 47912 17292 47961 17320
rect 47912 17280 47918 17292
rect 47949 17289 47961 17292
rect 47995 17289 48007 17323
rect 47949 17283 48007 17289
rect 55186 17292 57100 17320
rect 46750 17212 46756 17264
rect 46808 17252 46814 17264
rect 55186 17252 55214 17292
rect 46808 17224 55214 17252
rect 46808 17212 46814 17224
rect 42978 17144 42984 17196
rect 43036 17184 43042 17196
rect 44913 17187 44971 17193
rect 44913 17184 44925 17187
rect 43036 17156 44925 17184
rect 43036 17144 43042 17156
rect 44913 17153 44925 17156
rect 44959 17184 44971 17187
rect 44959 17156 46796 17184
rect 44959 17153 44971 17156
rect 44913 17147 44971 17153
rect 46290 17076 46296 17128
rect 46348 17116 46354 17128
rect 46477 17119 46535 17125
rect 46477 17116 46489 17119
rect 46348 17088 46489 17116
rect 46348 17076 46354 17088
rect 46477 17085 46489 17088
rect 46523 17085 46535 17119
rect 46477 17079 46535 17085
rect 46569 17119 46627 17125
rect 46569 17085 46581 17119
rect 46615 17085 46627 17119
rect 46569 17079 46627 17085
rect 45002 16980 45008 16992
rect 44963 16952 45008 16980
rect 45002 16940 45008 16952
rect 45060 16980 45066 16992
rect 46584 16980 46612 17079
rect 46768 17048 46796 17156
rect 56318 17144 56324 17196
rect 56376 17184 56382 17196
rect 57072 17193 57100 17292
rect 56597 17187 56655 17193
rect 56597 17184 56609 17187
rect 56376 17156 56609 17184
rect 56376 17144 56382 17156
rect 56597 17153 56609 17156
rect 56643 17153 56655 17187
rect 56597 17147 56655 17153
rect 57057 17187 57115 17193
rect 57057 17153 57069 17187
rect 57103 17153 57115 17187
rect 57057 17147 57115 17153
rect 57606 17144 57612 17196
rect 57664 17184 57670 17196
rect 57885 17187 57943 17193
rect 57885 17184 57897 17187
rect 57664 17156 57897 17184
rect 57664 17144 57670 17156
rect 57885 17153 57897 17156
rect 57931 17153 57943 17187
rect 57885 17147 57943 17153
rect 48038 17116 48044 17128
rect 47999 17088 48044 17116
rect 48038 17076 48044 17088
rect 48096 17076 48102 17128
rect 48222 17116 48228 17128
rect 48183 17088 48228 17116
rect 48222 17076 48228 17088
rect 48280 17076 48286 17128
rect 55766 17048 55772 17060
rect 46768 17020 55772 17048
rect 55766 17008 55772 17020
rect 55824 17008 55830 17060
rect 56413 17051 56471 17057
rect 56413 17017 56425 17051
rect 56459 17048 56471 17051
rect 56870 17048 56876 17060
rect 56459 17020 56876 17048
rect 56459 17017 56471 17020
rect 56413 17011 56471 17017
rect 56870 17008 56876 17020
rect 56928 17008 56934 17060
rect 57238 17048 57244 17060
rect 57199 17020 57244 17048
rect 57238 17008 57244 17020
rect 57296 17008 57302 17060
rect 48222 16980 48228 16992
rect 45060 16952 48228 16980
rect 45060 16940 45066 16952
rect 48222 16940 48228 16952
rect 48280 16940 48286 16992
rect 58066 16980 58072 16992
rect 58027 16952 58072 16980
rect 58066 16940 58072 16952
rect 58124 16940 58130 16992
rect 1104 16890 58880 16912
rect 1104 16838 10582 16890
rect 10634 16838 10646 16890
rect 10698 16838 10710 16890
rect 10762 16838 10774 16890
rect 10826 16838 10838 16890
rect 10890 16838 29846 16890
rect 29898 16838 29910 16890
rect 29962 16838 29974 16890
rect 30026 16838 30038 16890
rect 30090 16838 30102 16890
rect 30154 16838 49110 16890
rect 49162 16838 49174 16890
rect 49226 16838 49238 16890
rect 49290 16838 49302 16890
rect 49354 16838 49366 16890
rect 49418 16838 58880 16890
rect 1104 16816 58880 16838
rect 45002 16736 45008 16788
rect 45060 16736 45066 16788
rect 57146 16736 57152 16788
rect 57204 16776 57210 16788
rect 57241 16779 57299 16785
rect 57241 16776 57253 16779
rect 57204 16748 57253 16776
rect 57204 16736 57210 16748
rect 57241 16745 57253 16748
rect 57287 16745 57299 16779
rect 57241 16739 57299 16745
rect 45020 16708 45048 16736
rect 44284 16680 45600 16708
rect 43530 16600 43536 16652
rect 43588 16640 43594 16652
rect 44284 16649 44312 16680
rect 44085 16643 44143 16649
rect 44085 16640 44097 16643
rect 43588 16612 44097 16640
rect 43588 16600 43594 16612
rect 44085 16609 44097 16612
rect 44131 16609 44143 16643
rect 44085 16603 44143 16609
rect 44269 16643 44327 16649
rect 44269 16609 44281 16643
rect 44315 16609 44327 16643
rect 44269 16603 44327 16609
rect 45002 16600 45008 16652
rect 45060 16640 45066 16652
rect 45572 16649 45600 16680
rect 57054 16668 57060 16720
rect 57112 16708 57118 16720
rect 59170 16708 59176 16720
rect 57112 16680 59176 16708
rect 57112 16668 57118 16680
rect 59170 16668 59176 16680
rect 59228 16668 59234 16720
rect 45465 16643 45523 16649
rect 45465 16640 45477 16643
rect 45060 16612 45477 16640
rect 45060 16600 45066 16612
rect 45465 16609 45477 16612
rect 45511 16609 45523 16643
rect 45465 16603 45523 16609
rect 45557 16643 45615 16649
rect 45557 16609 45569 16643
rect 45603 16609 45615 16643
rect 45557 16603 45615 16609
rect 43990 16572 43996 16584
rect 43951 16544 43996 16572
rect 43990 16532 43996 16544
rect 44048 16532 44054 16584
rect 45370 16572 45376 16584
rect 45331 16544 45376 16572
rect 45370 16532 45376 16544
rect 45428 16532 45434 16584
rect 46385 16575 46443 16581
rect 46385 16572 46397 16575
rect 45526 16544 46397 16572
rect 45526 16504 45554 16544
rect 46385 16541 46397 16544
rect 46431 16541 46443 16575
rect 46385 16535 46443 16541
rect 56781 16575 56839 16581
rect 56781 16541 56793 16575
rect 56827 16572 56839 16575
rect 57054 16572 57060 16584
rect 56827 16544 57060 16572
rect 56827 16541 56839 16544
rect 56781 16535 56839 16541
rect 57054 16532 57060 16544
rect 57112 16532 57118 16584
rect 57422 16572 57428 16584
rect 57383 16544 57428 16572
rect 57422 16532 57428 16544
rect 57480 16532 57486 16584
rect 57882 16572 57888 16584
rect 57843 16544 57888 16572
rect 57882 16532 57888 16544
rect 57940 16532 57946 16584
rect 57606 16504 57612 16516
rect 45020 16476 45554 16504
rect 46216 16476 57612 16504
rect 43622 16436 43628 16448
rect 43583 16408 43628 16436
rect 43622 16396 43628 16408
rect 43680 16396 43686 16448
rect 45020 16445 45048 16476
rect 46216 16445 46244 16476
rect 57606 16464 57612 16476
rect 57664 16464 57670 16516
rect 45005 16439 45063 16445
rect 45005 16405 45017 16439
rect 45051 16405 45063 16439
rect 45005 16399 45063 16405
rect 46201 16439 46259 16445
rect 46201 16405 46213 16439
rect 46247 16405 46259 16439
rect 56594 16436 56600 16448
rect 56555 16408 56600 16436
rect 46201 16399 46259 16405
rect 56594 16396 56600 16408
rect 56652 16396 56658 16448
rect 58066 16436 58072 16448
rect 58027 16408 58072 16436
rect 58066 16396 58072 16408
rect 58124 16396 58130 16448
rect 1104 16346 58880 16368
rect 1104 16294 20214 16346
rect 20266 16294 20278 16346
rect 20330 16294 20342 16346
rect 20394 16294 20406 16346
rect 20458 16294 20470 16346
rect 20522 16294 39478 16346
rect 39530 16294 39542 16346
rect 39594 16294 39606 16346
rect 39658 16294 39670 16346
rect 39722 16294 39734 16346
rect 39786 16294 58880 16346
rect 1104 16272 58880 16294
rect 57149 16235 57207 16241
rect 57149 16201 57161 16235
rect 57195 16232 57207 16235
rect 57514 16232 57520 16244
rect 57195 16204 57520 16232
rect 57195 16201 57207 16204
rect 57149 16195 57207 16201
rect 57514 16192 57520 16204
rect 57572 16192 57578 16244
rect 43622 16056 43628 16108
rect 43680 16096 43686 16108
rect 44545 16099 44603 16105
rect 44545 16096 44557 16099
rect 43680 16068 44557 16096
rect 43680 16056 43686 16068
rect 44545 16065 44557 16068
rect 44591 16065 44603 16099
rect 57330 16096 57336 16108
rect 57291 16068 57336 16096
rect 44545 16059 44603 16065
rect 57330 16056 57336 16068
rect 57388 16056 57394 16108
rect 57422 16056 57428 16108
rect 57480 16096 57486 16108
rect 57885 16099 57943 16105
rect 57885 16096 57897 16099
rect 57480 16068 57897 16096
rect 57480 16056 57486 16068
rect 57885 16065 57897 16068
rect 57931 16065 57943 16099
rect 57885 16059 57943 16065
rect 44361 15895 44419 15901
rect 44361 15861 44373 15895
rect 44407 15892 44419 15895
rect 57882 15892 57888 15904
rect 44407 15864 57888 15892
rect 44407 15861 44419 15864
rect 44361 15855 44419 15861
rect 57882 15852 57888 15864
rect 57940 15852 57946 15904
rect 58066 15892 58072 15904
rect 58027 15864 58072 15892
rect 58066 15852 58072 15864
rect 58124 15852 58130 15904
rect 1104 15802 58880 15824
rect 1104 15750 10582 15802
rect 10634 15750 10646 15802
rect 10698 15750 10710 15802
rect 10762 15750 10774 15802
rect 10826 15750 10838 15802
rect 10890 15750 29846 15802
rect 29898 15750 29910 15802
rect 29962 15750 29974 15802
rect 30026 15750 30038 15802
rect 30090 15750 30102 15802
rect 30154 15750 49110 15802
rect 49162 15750 49174 15802
rect 49226 15750 49238 15802
rect 49290 15750 49302 15802
rect 49354 15750 49366 15802
rect 49418 15750 58880 15802
rect 1104 15728 58880 15750
rect 42058 15552 42064 15564
rect 42019 15524 42064 15552
rect 42058 15512 42064 15524
rect 42116 15512 42122 15564
rect 41874 15484 41880 15496
rect 41835 15456 41880 15484
rect 41874 15444 41880 15456
rect 41932 15444 41938 15496
rect 56594 15444 56600 15496
rect 56652 15484 56658 15496
rect 57885 15487 57943 15493
rect 57885 15484 57897 15487
rect 56652 15456 57897 15484
rect 56652 15444 56658 15456
rect 57885 15453 57897 15456
rect 57931 15453 57943 15487
rect 57885 15447 57943 15453
rect 41509 15351 41567 15357
rect 41509 15317 41521 15351
rect 41555 15348 41567 15351
rect 41874 15348 41880 15360
rect 41555 15320 41880 15348
rect 41555 15317 41567 15320
rect 41509 15311 41567 15317
rect 41874 15308 41880 15320
rect 41932 15308 41938 15360
rect 41969 15351 42027 15357
rect 41969 15317 41981 15351
rect 42015 15348 42027 15351
rect 42334 15348 42340 15360
rect 42015 15320 42340 15348
rect 42015 15317 42027 15320
rect 41969 15311 42027 15317
rect 42334 15308 42340 15320
rect 42392 15308 42398 15360
rect 57882 15308 57888 15360
rect 57940 15348 57946 15360
rect 58069 15351 58127 15357
rect 58069 15348 58081 15351
rect 57940 15320 58081 15348
rect 57940 15308 57946 15320
rect 58069 15317 58081 15320
rect 58115 15317 58127 15351
rect 58069 15311 58127 15317
rect 1104 15258 58880 15280
rect 1104 15206 20214 15258
rect 20266 15206 20278 15258
rect 20330 15206 20342 15258
rect 20394 15206 20406 15258
rect 20458 15206 20470 15258
rect 20522 15206 39478 15258
rect 39530 15206 39542 15258
rect 39594 15206 39606 15258
rect 39658 15206 39670 15258
rect 39722 15206 39734 15258
rect 39786 15206 58880 15258
rect 1104 15184 58880 15206
rect 39298 15144 39304 15156
rect 39259 15116 39304 15144
rect 39298 15104 39304 15116
rect 39356 15104 39362 15156
rect 57422 15076 57428 15088
rect 45526 15048 57428 15076
rect 39393 15011 39451 15017
rect 39393 14977 39405 15011
rect 39439 15008 39451 15011
rect 39758 15008 39764 15020
rect 39439 14980 39764 15008
rect 39439 14977 39451 14980
rect 39393 14971 39451 14977
rect 39758 14968 39764 14980
rect 39816 14968 39822 15020
rect 41325 15011 41383 15017
rect 41325 14977 41337 15011
rect 41371 15008 41383 15011
rect 42705 15011 42763 15017
rect 41371 14980 42656 15008
rect 41371 14977 41383 14980
rect 41325 14971 41383 14977
rect 39577 14943 39635 14949
rect 39577 14909 39589 14943
rect 39623 14909 39635 14943
rect 39577 14903 39635 14909
rect 41049 14943 41107 14949
rect 41049 14909 41061 14943
rect 41095 14940 41107 14943
rect 41138 14940 41144 14952
rect 41095 14912 41144 14940
rect 41095 14909 41107 14912
rect 41049 14903 41107 14909
rect 38102 14832 38108 14884
rect 38160 14872 38166 14884
rect 39592 14872 39620 14903
rect 41138 14900 41144 14912
rect 41196 14900 41202 14952
rect 41874 14900 41880 14952
rect 41932 14940 41938 14952
rect 42429 14943 42487 14949
rect 42429 14940 42441 14943
rect 41932 14912 42441 14940
rect 41932 14900 41938 14912
rect 42429 14909 42441 14912
rect 42475 14909 42487 14943
rect 42628 14940 42656 14980
rect 42705 14977 42717 15011
rect 42751 15008 42763 15011
rect 45526 15008 45554 15048
rect 57422 15036 57428 15048
rect 57480 15036 57486 15088
rect 42751 14980 45554 15008
rect 42751 14977 42763 14980
rect 42705 14971 42763 14977
rect 50246 14968 50252 15020
rect 50304 15008 50310 15020
rect 57885 15011 57943 15017
rect 57885 15008 57897 15011
rect 50304 14980 57897 15008
rect 50304 14968 50310 14980
rect 57885 14977 57897 14980
rect 57931 14977 57943 15011
rect 57885 14971 57943 14977
rect 56594 14940 56600 14952
rect 42628 14912 56600 14940
rect 42429 14903 42487 14909
rect 56594 14900 56600 14912
rect 56652 14900 56658 14952
rect 42058 14872 42064 14884
rect 38160 14844 42064 14872
rect 38160 14832 38166 14844
rect 42058 14832 42064 14844
rect 42116 14832 42122 14884
rect 38933 14807 38991 14813
rect 38933 14773 38945 14807
rect 38979 14804 38991 14807
rect 39850 14804 39856 14816
rect 38979 14776 39856 14804
rect 38979 14773 38991 14776
rect 38933 14767 38991 14773
rect 39850 14764 39856 14776
rect 39908 14764 39914 14816
rect 58066 14804 58072 14816
rect 58027 14776 58072 14804
rect 58066 14764 58072 14776
rect 58124 14764 58130 14816
rect 1104 14714 58880 14736
rect 1104 14662 10582 14714
rect 10634 14662 10646 14714
rect 10698 14662 10710 14714
rect 10762 14662 10774 14714
rect 10826 14662 10838 14714
rect 10890 14662 29846 14714
rect 29898 14662 29910 14714
rect 29962 14662 29974 14714
rect 30026 14662 30038 14714
rect 30090 14662 30102 14714
rect 30154 14662 49110 14714
rect 49162 14662 49174 14714
rect 49226 14662 49238 14714
rect 49290 14662 49302 14714
rect 49354 14662 49366 14714
rect 49418 14662 58880 14714
rect 1104 14640 58880 14662
rect 41138 14600 41144 14612
rect 41099 14572 41144 14600
rect 41138 14560 41144 14572
rect 41196 14560 41202 14612
rect 38102 14464 38108 14476
rect 38063 14436 38108 14464
rect 38102 14424 38108 14436
rect 38160 14424 38166 14476
rect 39850 14464 39856 14476
rect 39811 14436 39856 14464
rect 39850 14424 39856 14436
rect 39908 14424 39914 14476
rect 41785 14467 41843 14473
rect 41785 14433 41797 14467
rect 41831 14464 41843 14467
rect 42058 14464 42064 14476
rect 41831 14436 42064 14464
rect 41831 14433 41843 14436
rect 41785 14427 41843 14433
rect 42058 14424 42064 14436
rect 42116 14424 42122 14476
rect 37826 14396 37832 14408
rect 37787 14368 37832 14396
rect 37826 14356 37832 14368
rect 37884 14356 37890 14408
rect 40129 14399 40187 14405
rect 40129 14365 40141 14399
rect 40175 14396 40187 14399
rect 50246 14396 50252 14408
rect 40175 14368 50252 14396
rect 40175 14365 40187 14368
rect 40129 14359 40187 14365
rect 50246 14356 50252 14368
rect 50304 14356 50310 14408
rect 50338 14356 50344 14408
rect 50396 14396 50402 14408
rect 57885 14399 57943 14405
rect 57885 14396 57897 14399
rect 50396 14368 57897 14396
rect 50396 14356 50402 14368
rect 57885 14365 57897 14368
rect 57931 14365 57943 14399
rect 57885 14359 57943 14365
rect 41506 14328 41512 14340
rect 41467 14300 41512 14328
rect 41506 14288 41512 14300
rect 41564 14288 41570 14340
rect 37458 14260 37464 14272
rect 37419 14232 37464 14260
rect 37458 14220 37464 14232
rect 37516 14220 37522 14272
rect 37734 14220 37740 14272
rect 37792 14260 37798 14272
rect 37921 14263 37979 14269
rect 37921 14260 37933 14263
rect 37792 14232 37933 14260
rect 37792 14220 37798 14232
rect 37921 14229 37933 14232
rect 37967 14229 37979 14263
rect 37921 14223 37979 14229
rect 41598 14220 41604 14272
rect 41656 14260 41662 14272
rect 58066 14260 58072 14272
rect 41656 14232 41701 14260
rect 58027 14232 58072 14260
rect 41656 14220 41662 14232
rect 58066 14220 58072 14232
rect 58124 14220 58130 14272
rect 1104 14170 58880 14192
rect 1104 14118 20214 14170
rect 20266 14118 20278 14170
rect 20330 14118 20342 14170
rect 20394 14118 20406 14170
rect 20458 14118 20470 14170
rect 20522 14118 39478 14170
rect 39530 14118 39542 14170
rect 39594 14118 39606 14170
rect 39658 14118 39670 14170
rect 39722 14118 39734 14170
rect 39786 14118 58880 14170
rect 1104 14096 58880 14118
rect 57882 14016 57888 14068
rect 57940 14056 57946 14068
rect 58069 14059 58127 14065
rect 58069 14056 58081 14059
rect 57940 14028 58081 14056
rect 57940 14016 57946 14028
rect 58069 14025 58081 14028
rect 58115 14025 58127 14059
rect 58069 14019 58127 14025
rect 37458 13880 37464 13932
rect 37516 13920 37522 13932
rect 38197 13923 38255 13929
rect 38197 13920 38209 13923
rect 37516 13892 38209 13920
rect 37516 13880 37522 13892
rect 38197 13889 38209 13892
rect 38243 13889 38255 13923
rect 38197 13883 38255 13889
rect 52454 13880 52460 13932
rect 52512 13920 52518 13932
rect 57885 13923 57943 13929
rect 57885 13920 57897 13923
rect 52512 13892 57897 13920
rect 52512 13880 52518 13892
rect 57885 13889 57897 13892
rect 57931 13889 57943 13923
rect 57885 13883 57943 13889
rect 38473 13855 38531 13861
rect 38473 13821 38485 13855
rect 38519 13852 38531 13855
rect 50338 13852 50344 13864
rect 38519 13824 50344 13852
rect 38519 13821 38531 13824
rect 38473 13815 38531 13821
rect 50338 13812 50344 13824
rect 50396 13812 50402 13864
rect 1104 13626 58880 13648
rect 1104 13574 10582 13626
rect 10634 13574 10646 13626
rect 10698 13574 10710 13626
rect 10762 13574 10774 13626
rect 10826 13574 10838 13626
rect 10890 13574 29846 13626
rect 29898 13574 29910 13626
rect 29962 13574 29974 13626
rect 30026 13574 30038 13626
rect 30090 13574 30102 13626
rect 30154 13574 49110 13626
rect 49162 13574 49174 13626
rect 49226 13574 49238 13626
rect 49290 13574 49302 13626
rect 49354 13574 49366 13626
rect 49418 13574 58880 13626
rect 1104 13552 58880 13574
rect 36081 13447 36139 13453
rect 36081 13413 36093 13447
rect 36127 13444 36139 13447
rect 36127 13416 37320 13444
rect 36127 13413 36139 13416
rect 36081 13407 36139 13413
rect 37292 13385 37320 13416
rect 36725 13379 36783 13385
rect 36725 13345 36737 13379
rect 36771 13345 36783 13379
rect 36725 13339 36783 13345
rect 37277 13379 37335 13385
rect 37277 13345 37289 13379
rect 37323 13345 37335 13379
rect 37277 13339 37335 13345
rect 36446 13308 36452 13320
rect 36407 13280 36452 13308
rect 36446 13268 36452 13280
rect 36504 13268 36510 13320
rect 36740 13240 36768 13339
rect 37553 13311 37611 13317
rect 37553 13277 37565 13311
rect 37599 13308 37611 13311
rect 52454 13308 52460 13320
rect 37599 13280 52460 13308
rect 37599 13277 37611 13280
rect 37553 13271 37611 13277
rect 52454 13268 52460 13280
rect 52512 13268 52518 13320
rect 52546 13268 52552 13320
rect 52604 13308 52610 13320
rect 57885 13311 57943 13317
rect 57885 13308 57897 13311
rect 52604 13280 57897 13308
rect 52604 13268 52610 13280
rect 57885 13277 57897 13280
rect 57931 13277 57943 13311
rect 57885 13271 57943 13277
rect 38102 13240 38108 13252
rect 36740 13212 38108 13240
rect 38102 13200 38108 13212
rect 38160 13200 38166 13252
rect 36354 13132 36360 13184
rect 36412 13172 36418 13184
rect 36541 13175 36599 13181
rect 36541 13172 36553 13175
rect 36412 13144 36553 13172
rect 36412 13132 36418 13144
rect 36541 13141 36553 13144
rect 36587 13141 36599 13175
rect 58066 13172 58072 13184
rect 58027 13144 58072 13172
rect 36541 13135 36599 13141
rect 58066 13132 58072 13144
rect 58124 13132 58130 13184
rect 1104 13082 58880 13104
rect 1104 13030 20214 13082
rect 20266 13030 20278 13082
rect 20330 13030 20342 13082
rect 20394 13030 20406 13082
rect 20458 13030 20470 13082
rect 20522 13030 39478 13082
rect 39530 13030 39542 13082
rect 39594 13030 39606 13082
rect 39658 13030 39670 13082
rect 39722 13030 39734 13082
rect 39786 13030 58880 13082
rect 1104 13008 58880 13030
rect 38102 12928 38108 12980
rect 38160 12968 38166 12980
rect 38289 12971 38347 12977
rect 38289 12968 38301 12971
rect 38160 12940 38301 12968
rect 38160 12928 38166 12940
rect 38289 12937 38301 12940
rect 38335 12937 38347 12971
rect 38289 12931 38347 12937
rect 35158 12832 35164 12844
rect 35119 12804 35164 12832
rect 35158 12792 35164 12804
rect 35216 12792 35222 12844
rect 38197 12835 38255 12841
rect 38197 12801 38209 12835
rect 38243 12832 38255 12835
rect 38378 12832 38384 12844
rect 38243 12804 38384 12832
rect 38243 12801 38255 12804
rect 38197 12795 38255 12801
rect 38378 12792 38384 12804
rect 38436 12792 38442 12844
rect 57425 12835 57483 12841
rect 57425 12832 57437 12835
rect 45526 12804 57437 12832
rect 34238 12724 34244 12776
rect 34296 12764 34302 12776
rect 45526 12764 45554 12804
rect 57425 12801 57437 12804
rect 57471 12832 57483 12835
rect 57885 12835 57943 12841
rect 57885 12832 57897 12835
rect 57471 12804 57897 12832
rect 57471 12801 57483 12804
rect 57425 12795 57483 12801
rect 57885 12801 57897 12804
rect 57931 12801 57943 12835
rect 57885 12795 57943 12801
rect 34296 12736 45554 12764
rect 34296 12724 34302 12736
rect 35345 12699 35403 12705
rect 35345 12665 35357 12699
rect 35391 12696 35403 12699
rect 52546 12696 52552 12708
rect 35391 12668 52552 12696
rect 35391 12665 35403 12668
rect 35345 12659 35403 12665
rect 52546 12656 52552 12668
rect 52604 12656 52610 12708
rect 58066 12628 58072 12640
rect 58027 12600 58072 12628
rect 58066 12588 58072 12600
rect 58124 12588 58130 12640
rect 1104 12538 58880 12560
rect 1104 12486 10582 12538
rect 10634 12486 10646 12538
rect 10698 12486 10710 12538
rect 10762 12486 10774 12538
rect 10826 12486 10838 12538
rect 10890 12486 29846 12538
rect 29898 12486 29910 12538
rect 29962 12486 29974 12538
rect 30026 12486 30038 12538
rect 30090 12486 30102 12538
rect 30154 12486 49110 12538
rect 49162 12486 49174 12538
rect 49226 12486 49238 12538
rect 49290 12486 49302 12538
rect 49354 12486 49366 12538
rect 49418 12486 58880 12538
rect 1104 12464 58880 12486
rect 34701 12427 34759 12433
rect 34701 12393 34713 12427
rect 34747 12424 34759 12427
rect 35158 12424 35164 12436
rect 34747 12396 35164 12424
rect 34747 12393 34759 12396
rect 34701 12387 34759 12393
rect 35158 12384 35164 12396
rect 35216 12384 35222 12436
rect 31389 12359 31447 12365
rect 31389 12325 31401 12359
rect 31435 12356 31447 12359
rect 31435 12328 35894 12356
rect 31435 12325 31447 12328
rect 31389 12319 31447 12325
rect 32766 12248 32772 12300
rect 32824 12288 32830 12300
rect 33965 12291 34023 12297
rect 33965 12288 33977 12291
rect 32824 12260 33977 12288
rect 32824 12248 32830 12260
rect 33965 12257 33977 12260
rect 34011 12288 34023 12291
rect 35253 12291 35311 12297
rect 35253 12288 35265 12291
rect 34011 12260 35265 12288
rect 34011 12257 34023 12260
rect 33965 12251 34023 12257
rect 35253 12257 35265 12260
rect 35299 12257 35311 12291
rect 35866 12288 35894 12328
rect 50338 12288 50344 12300
rect 35866 12260 50344 12288
rect 35253 12251 35311 12257
rect 50338 12248 50344 12260
rect 50396 12248 50402 12300
rect 33686 12220 33692 12232
rect 33647 12192 33692 12220
rect 33686 12180 33692 12192
rect 33744 12180 33750 12232
rect 35066 12220 35072 12232
rect 35027 12192 35072 12220
rect 35066 12180 35072 12192
rect 35124 12180 35130 12232
rect 38654 12220 38660 12232
rect 38615 12192 38660 12220
rect 38654 12180 38660 12192
rect 38712 12180 38718 12232
rect 57885 12223 57943 12229
rect 57885 12220 57897 12223
rect 45526 12192 57897 12220
rect 30650 12112 30656 12164
rect 30708 12152 30714 12164
rect 31205 12155 31263 12161
rect 31205 12152 31217 12155
rect 30708 12124 31217 12152
rect 30708 12112 30714 12124
rect 31205 12121 31217 12124
rect 31251 12121 31263 12155
rect 31205 12115 31263 12121
rect 32122 12112 32128 12164
rect 32180 12152 32186 12164
rect 32585 12155 32643 12161
rect 32585 12152 32597 12155
rect 32180 12124 32597 12152
rect 32180 12112 32186 12124
rect 32585 12121 32597 12124
rect 32631 12121 32643 12155
rect 32585 12115 32643 12121
rect 32769 12155 32827 12161
rect 32769 12121 32781 12155
rect 32815 12152 32827 12155
rect 45526 12152 45554 12192
rect 57885 12189 57897 12192
rect 57931 12189 57943 12223
rect 57885 12183 57943 12189
rect 32815 12124 45554 12152
rect 32815 12121 32827 12124
rect 32769 12115 32827 12121
rect 33318 12084 33324 12096
rect 33279 12056 33324 12084
rect 33318 12044 33324 12056
rect 33376 12044 33382 12096
rect 33594 12044 33600 12096
rect 33652 12084 33658 12096
rect 33781 12087 33839 12093
rect 33781 12084 33793 12087
rect 33652 12056 33793 12084
rect 33652 12044 33658 12056
rect 33781 12053 33793 12056
rect 33827 12053 33839 12087
rect 33781 12047 33839 12053
rect 34974 12044 34980 12096
rect 35032 12084 35038 12096
rect 35161 12087 35219 12093
rect 35161 12084 35173 12087
rect 35032 12056 35173 12084
rect 35032 12044 35038 12056
rect 35161 12053 35173 12056
rect 35207 12053 35219 12087
rect 35161 12047 35219 12053
rect 38378 12044 38384 12096
rect 38436 12084 38442 12096
rect 38841 12087 38899 12093
rect 38841 12084 38853 12087
rect 38436 12056 38853 12084
rect 38436 12044 38442 12056
rect 38841 12053 38853 12056
rect 38887 12053 38899 12087
rect 58066 12084 58072 12096
rect 58027 12056 58072 12084
rect 38841 12047 38899 12053
rect 58066 12044 58072 12056
rect 58124 12044 58130 12096
rect 1104 11994 58880 12016
rect 1104 11942 20214 11994
rect 20266 11942 20278 11994
rect 20330 11942 20342 11994
rect 20394 11942 20406 11994
rect 20458 11942 20470 11994
rect 20522 11942 39478 11994
rect 39530 11942 39542 11994
rect 39594 11942 39606 11994
rect 39658 11942 39670 11994
rect 39722 11942 39734 11994
rect 39786 11942 58880 11994
rect 1104 11920 58880 11942
rect 29638 11840 29644 11892
rect 29696 11880 29702 11892
rect 29825 11883 29883 11889
rect 29825 11880 29837 11883
rect 29696 11852 29837 11880
rect 29696 11840 29702 11852
rect 29825 11849 29837 11852
rect 29871 11849 29883 11883
rect 30650 11880 30656 11892
rect 30611 11852 30656 11880
rect 29825 11843 29883 11849
rect 30650 11840 30656 11852
rect 30708 11840 30714 11892
rect 31018 11880 31024 11892
rect 30979 11852 31024 11880
rect 31018 11840 31024 11852
rect 31076 11840 31082 11892
rect 32122 11880 32128 11892
rect 32083 11852 32128 11880
rect 32122 11840 32128 11852
rect 32180 11840 32186 11892
rect 32490 11880 32496 11892
rect 32451 11852 32496 11880
rect 32490 11840 32496 11852
rect 32548 11840 32554 11892
rect 33318 11772 33324 11824
rect 33376 11812 33382 11824
rect 34057 11815 34115 11821
rect 34057 11812 34069 11815
rect 33376 11784 34069 11812
rect 33376 11772 33382 11784
rect 34057 11781 34069 11784
rect 34103 11781 34115 11815
rect 34238 11812 34244 11824
rect 34199 11784 34244 11812
rect 34057 11775 34115 11781
rect 34238 11772 34244 11784
rect 34296 11772 34302 11824
rect 31018 11744 31024 11756
rect 30116 11716 31024 11744
rect 29546 11636 29552 11688
rect 29604 11676 29610 11688
rect 30116 11685 30144 11716
rect 31018 11704 31024 11716
rect 31076 11744 31082 11756
rect 31076 11716 31248 11744
rect 31076 11704 31082 11716
rect 29917 11679 29975 11685
rect 29917 11676 29929 11679
rect 29604 11648 29929 11676
rect 29604 11636 29610 11648
rect 29917 11645 29929 11648
rect 29963 11645 29975 11679
rect 29917 11639 29975 11645
rect 30101 11679 30159 11685
rect 30101 11645 30113 11679
rect 30147 11645 30159 11679
rect 30101 11639 30159 11645
rect 30742 11636 30748 11688
rect 30800 11676 30806 11688
rect 31220 11685 31248 11716
rect 50338 11704 50344 11756
rect 50396 11744 50402 11756
rect 57885 11747 57943 11753
rect 57885 11744 57897 11747
rect 50396 11716 57897 11744
rect 50396 11704 50402 11716
rect 57885 11713 57897 11716
rect 57931 11713 57943 11747
rect 57885 11707 57943 11713
rect 31113 11679 31171 11685
rect 31113 11676 31125 11679
rect 30800 11648 31125 11676
rect 30800 11636 30806 11648
rect 31113 11645 31125 11648
rect 31159 11645 31171 11679
rect 31113 11639 31171 11645
rect 31205 11679 31263 11685
rect 31205 11645 31217 11679
rect 31251 11676 31263 11679
rect 31251 11648 31754 11676
rect 31251 11645 31263 11648
rect 31205 11639 31263 11645
rect 31726 11608 31754 11648
rect 32122 11636 32128 11688
rect 32180 11676 32186 11688
rect 32585 11679 32643 11685
rect 32585 11676 32597 11679
rect 32180 11648 32597 11676
rect 32180 11636 32186 11648
rect 32585 11645 32597 11648
rect 32631 11645 32643 11679
rect 32766 11676 32772 11688
rect 32727 11648 32772 11676
rect 32585 11639 32643 11645
rect 32766 11636 32772 11648
rect 32824 11636 32830 11688
rect 32784 11608 32812 11636
rect 31726 11580 32812 11608
rect 29457 11543 29515 11549
rect 29457 11509 29469 11543
rect 29503 11540 29515 11543
rect 30190 11540 30196 11552
rect 29503 11512 30196 11540
rect 29503 11509 29515 11512
rect 29457 11503 29515 11509
rect 30190 11500 30196 11512
rect 30248 11500 30254 11552
rect 58066 11540 58072 11552
rect 58027 11512 58072 11540
rect 58066 11500 58072 11512
rect 58124 11500 58130 11552
rect 1104 11450 58880 11472
rect 1104 11398 10582 11450
rect 10634 11398 10646 11450
rect 10698 11398 10710 11450
rect 10762 11398 10774 11450
rect 10826 11398 10838 11450
rect 10890 11398 29846 11450
rect 29898 11398 29910 11450
rect 29962 11398 29974 11450
rect 30026 11398 30038 11450
rect 30090 11398 30102 11450
rect 30154 11398 49110 11450
rect 49162 11398 49174 11450
rect 49226 11398 49238 11450
rect 49290 11398 49302 11450
rect 49354 11398 49366 11450
rect 49418 11398 58880 11450
rect 1104 11376 58880 11398
rect 31018 11336 31024 11348
rect 30979 11308 31024 11336
rect 31018 11296 31024 11308
rect 31076 11296 31082 11348
rect 38654 11228 38660 11280
rect 38712 11268 38718 11280
rect 42978 11268 42984 11280
rect 38712 11240 42984 11268
rect 38712 11228 38718 11240
rect 30190 11132 30196 11144
rect 30151 11104 30196 11132
rect 30190 11092 30196 11104
rect 30248 11092 30254 11144
rect 39868 11141 39896 11240
rect 42978 11228 42984 11240
rect 43036 11228 43042 11280
rect 57882 11228 57888 11280
rect 57940 11268 57946 11280
rect 58069 11271 58127 11277
rect 58069 11268 58081 11271
rect 57940 11240 58081 11268
rect 57940 11228 57946 11240
rect 58069 11237 58081 11240
rect 58115 11237 58127 11271
rect 58069 11231 58127 11237
rect 40218 11160 40224 11212
rect 40276 11200 40282 11212
rect 56778 11200 56784 11212
rect 40276 11172 56784 11200
rect 40276 11160 40282 11172
rect 56778 11160 56784 11172
rect 56836 11160 56842 11212
rect 30377 11135 30435 11141
rect 30377 11101 30389 11135
rect 30423 11132 30435 11135
rect 39853 11135 39911 11141
rect 30423 11104 39804 11132
rect 30423 11101 30435 11104
rect 30377 11095 30435 11101
rect 26510 11024 26516 11076
rect 26568 11064 26574 11076
rect 30929 11067 30987 11073
rect 30929 11064 30941 11067
rect 26568 11036 30941 11064
rect 26568 11024 26574 11036
rect 30929 11033 30941 11036
rect 30975 11064 30987 11067
rect 38378 11064 38384 11076
rect 30975 11036 38384 11064
rect 30975 11033 30987 11036
rect 30929 11027 30987 11033
rect 38378 11024 38384 11036
rect 38436 11024 38442 11076
rect 39776 11064 39804 11104
rect 39853 11101 39865 11135
rect 39899 11101 39911 11135
rect 57885 11135 57943 11141
rect 57885 11132 57897 11135
rect 39853 11095 39911 11101
rect 40052 11104 57897 11132
rect 40052 11064 40080 11104
rect 57885 11101 57897 11104
rect 57931 11101 57943 11135
rect 57885 11095 57943 11101
rect 39776 11036 40080 11064
rect 40129 11067 40187 11073
rect 40129 11033 40141 11067
rect 40175 11064 40187 11067
rect 40218 11064 40224 11076
rect 40175 11036 40224 11064
rect 40175 11033 40187 11036
rect 40129 11027 40187 11033
rect 40218 11024 40224 11036
rect 40276 11024 40282 11076
rect 1104 10906 58880 10928
rect 1104 10854 20214 10906
rect 20266 10854 20278 10906
rect 20330 10854 20342 10906
rect 20394 10854 20406 10906
rect 20458 10854 20470 10906
rect 20522 10854 39478 10906
rect 39530 10854 39542 10906
rect 39594 10854 39606 10906
rect 39658 10854 39670 10906
rect 39722 10854 39734 10906
rect 39786 10854 58880 10906
rect 1104 10832 58880 10854
rect 57054 10656 57060 10668
rect 57015 10628 57060 10656
rect 57054 10616 57060 10628
rect 57112 10616 57118 10668
rect 57146 10616 57152 10668
rect 57204 10656 57210 10668
rect 57885 10659 57943 10665
rect 57885 10656 57897 10659
rect 57204 10628 57897 10656
rect 57204 10616 57210 10628
rect 57885 10625 57897 10628
rect 57931 10625 57943 10659
rect 57885 10619 57943 10625
rect 57238 10452 57244 10464
rect 57199 10424 57244 10452
rect 57238 10412 57244 10424
rect 57296 10412 57302 10464
rect 58066 10452 58072 10464
rect 58027 10424 58072 10452
rect 58066 10412 58072 10424
rect 58124 10412 58130 10464
rect 1104 10362 58880 10384
rect 1104 10310 10582 10362
rect 10634 10310 10646 10362
rect 10698 10310 10710 10362
rect 10762 10310 10774 10362
rect 10826 10310 10838 10362
rect 10890 10310 29846 10362
rect 29898 10310 29910 10362
rect 29962 10310 29974 10362
rect 30026 10310 30038 10362
rect 30090 10310 30102 10362
rect 30154 10310 49110 10362
rect 49162 10310 49174 10362
rect 49226 10310 49238 10362
rect 49290 10310 49302 10362
rect 49354 10310 49366 10362
rect 49418 10310 58880 10362
rect 1104 10288 58880 10310
rect 28077 10251 28135 10257
rect 28077 10217 28089 10251
rect 28123 10248 28135 10251
rect 28123 10220 35894 10248
rect 28123 10217 28135 10220
rect 28077 10211 28135 10217
rect 27065 10047 27123 10053
rect 27065 10013 27077 10047
rect 27111 10044 27123 10047
rect 35866 10044 35894 10220
rect 57054 10044 57060 10056
rect 27111 10016 31754 10044
rect 35866 10016 57060 10044
rect 27111 10013 27123 10016
rect 27065 10007 27123 10013
rect 26878 9976 26884 9988
rect 26839 9948 26884 9976
rect 26878 9936 26884 9948
rect 26936 9936 26942 9988
rect 27982 9976 27988 9988
rect 27943 9948 27988 9976
rect 27982 9936 27988 9948
rect 28040 9936 28046 9988
rect 31726 9976 31754 10016
rect 57054 10004 57060 10016
rect 57112 10004 57118 10056
rect 57885 10047 57943 10053
rect 57885 10044 57897 10047
rect 57532 10016 57897 10044
rect 57146 9976 57152 9988
rect 31726 9948 57152 9976
rect 57146 9936 57152 9948
rect 57204 9936 57210 9988
rect 26050 9868 26056 9920
rect 26108 9908 26114 9920
rect 57532 9917 57560 10016
rect 57885 10013 57897 10016
rect 57931 10013 57943 10047
rect 57885 10007 57943 10013
rect 57517 9911 57575 9917
rect 57517 9908 57529 9911
rect 26108 9880 57529 9908
rect 26108 9868 26114 9880
rect 57517 9877 57529 9880
rect 57563 9877 57575 9911
rect 57517 9871 57575 9877
rect 57882 9868 57888 9920
rect 57940 9908 57946 9920
rect 58069 9911 58127 9917
rect 58069 9908 58081 9911
rect 57940 9880 58081 9908
rect 57940 9868 57946 9880
rect 58069 9877 58081 9880
rect 58115 9877 58127 9911
rect 58069 9871 58127 9877
rect 1104 9818 58880 9840
rect 1104 9766 20214 9818
rect 20266 9766 20278 9818
rect 20330 9766 20342 9818
rect 20394 9766 20406 9818
rect 20458 9766 20470 9818
rect 20522 9766 39478 9818
rect 39530 9766 39542 9818
rect 39594 9766 39606 9818
rect 39658 9766 39670 9818
rect 39722 9766 39734 9818
rect 39786 9766 58880 9818
rect 1104 9744 58880 9766
rect 26878 9664 26884 9716
rect 26936 9704 26942 9716
rect 26973 9707 27031 9713
rect 26973 9704 26985 9707
rect 26936 9676 26985 9704
rect 26936 9664 26942 9676
rect 26973 9673 26985 9676
rect 27019 9673 27031 9707
rect 26973 9667 27031 9673
rect 24946 9636 24952 9648
rect 24907 9608 24952 9636
rect 24946 9596 24952 9608
rect 25004 9596 25010 9648
rect 26050 9636 26056 9648
rect 26011 9608 26056 9636
rect 26050 9596 26056 9608
rect 26108 9596 26114 9648
rect 27338 9636 27344 9648
rect 27299 9608 27344 9636
rect 27338 9596 27344 9608
rect 27396 9596 27402 9648
rect 25869 9571 25927 9577
rect 25869 9568 25881 9571
rect 24596 9540 25881 9568
rect 24596 9441 24624 9540
rect 25869 9537 25881 9540
rect 25915 9537 25927 9571
rect 25869 9531 25927 9537
rect 50338 9528 50344 9580
rect 50396 9568 50402 9580
rect 57885 9571 57943 9577
rect 57885 9568 57897 9571
rect 50396 9540 57897 9568
rect 50396 9528 50402 9540
rect 57885 9537 57897 9540
rect 57931 9537 57943 9571
rect 57885 9531 57943 9537
rect 25038 9500 25044 9512
rect 24999 9472 25044 9500
rect 25038 9460 25044 9472
rect 25096 9460 25102 9512
rect 25133 9503 25191 9509
rect 25133 9469 25145 9503
rect 25179 9469 25191 9503
rect 27430 9500 27436 9512
rect 27391 9472 27436 9500
rect 25133 9463 25191 9469
rect 24581 9435 24639 9441
rect 24581 9401 24593 9435
rect 24627 9401 24639 9435
rect 25148 9432 25176 9463
rect 27430 9460 27436 9472
rect 27488 9460 27494 9512
rect 27525 9503 27583 9509
rect 27525 9469 27537 9503
rect 27571 9469 27583 9503
rect 27525 9463 27583 9469
rect 24581 9395 24639 9401
rect 25056 9404 25176 9432
rect 23750 9324 23756 9376
rect 23808 9364 23814 9376
rect 25056 9364 25084 9404
rect 27338 9392 27344 9444
rect 27396 9432 27402 9444
rect 27540 9432 27568 9463
rect 27396 9404 27568 9432
rect 27396 9392 27402 9404
rect 58066 9364 58072 9376
rect 23808 9336 25084 9364
rect 58027 9336 58072 9364
rect 23808 9324 23814 9336
rect 58066 9324 58072 9336
rect 58124 9324 58130 9376
rect 1104 9274 58880 9296
rect 1104 9222 10582 9274
rect 10634 9222 10646 9274
rect 10698 9222 10710 9274
rect 10762 9222 10774 9274
rect 10826 9222 10838 9274
rect 10890 9222 29846 9274
rect 29898 9222 29910 9274
rect 29962 9222 29974 9274
rect 30026 9222 30038 9274
rect 30090 9222 30102 9274
rect 30154 9222 49110 9274
rect 49162 9222 49174 9274
rect 49226 9222 49238 9274
rect 49290 9222 49302 9274
rect 49354 9222 49366 9274
rect 49418 9222 58880 9274
rect 1104 9200 58880 9222
rect 10502 9120 10508 9172
rect 10560 9160 10566 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 10560 9132 10609 9160
rect 10560 9120 10566 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 12066 9160 12072 9172
rect 12027 9132 12072 9160
rect 10597 9123 10655 9129
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 14090 9160 14096 9172
rect 14051 9132 14096 9160
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 27157 9163 27215 9169
rect 27157 9129 27169 9163
rect 27203 9160 27215 9163
rect 27982 9160 27988 9172
rect 27203 9132 27988 9160
rect 27203 9129 27215 9132
rect 27157 9123 27215 9129
rect 27982 9120 27988 9132
rect 28040 9120 28046 9172
rect 24581 9095 24639 9101
rect 24581 9061 24593 9095
rect 24627 9092 24639 9095
rect 24627 9064 35894 9092
rect 24627 9061 24639 9064
rect 24581 9055 24639 9061
rect 1394 8984 1400 9036
rect 1452 9024 1458 9036
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 1452 8996 9413 9024
rect 1452 8984 1458 8996
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 22833 9027 22891 9033
rect 22833 8993 22845 9027
rect 22879 9024 22891 9027
rect 23750 9024 23756 9036
rect 22879 8996 23756 9024
rect 22879 8993 22891 8996
rect 22833 8987 22891 8993
rect 23750 8984 23756 8996
rect 23808 9024 23814 9036
rect 26697 9027 26755 9033
rect 26697 9024 26709 9027
rect 23808 8996 26709 9024
rect 23808 8984 23814 8996
rect 26697 8993 26709 8996
rect 26743 9024 26755 9027
rect 27338 9024 27344 9036
rect 26743 8996 27344 9024
rect 26743 8993 26755 8996
rect 26697 8987 26755 8993
rect 27338 8984 27344 8996
rect 27396 9024 27402 9036
rect 27709 9027 27767 9033
rect 27709 9024 27721 9027
rect 27396 8996 27721 9024
rect 27396 8984 27402 8996
rect 27709 8993 27721 8996
rect 27755 8993 27767 9027
rect 27709 8987 27767 8993
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8956 9183 8959
rect 9766 8956 9772 8968
rect 9171 8928 9772 8956
rect 9171 8925 9183 8928
rect 9125 8919 9183 8925
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8956 10839 8959
rect 10962 8956 10968 8968
rect 10827 8928 10968 8956
rect 10827 8925 10839 8928
rect 10781 8919 10839 8925
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 12253 8959 12311 8965
rect 12253 8925 12265 8959
rect 12299 8956 12311 8959
rect 12526 8956 12532 8968
rect 12299 8928 12532 8956
rect 12299 8925 12311 8928
rect 12253 8919 12311 8925
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 14274 8956 14280 8968
rect 14235 8928 14280 8956
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 22554 8956 22560 8968
rect 22515 8928 22560 8956
rect 22554 8916 22560 8928
rect 22612 8916 22618 8968
rect 23198 8916 23204 8968
rect 23256 8956 23262 8968
rect 24397 8959 24455 8965
rect 24397 8956 24409 8959
rect 23256 8928 24409 8956
rect 23256 8916 23262 8928
rect 24397 8925 24409 8928
rect 24443 8925 24455 8959
rect 24397 8919 24455 8925
rect 27525 8959 27583 8965
rect 27525 8925 27537 8959
rect 27571 8956 27583 8959
rect 27798 8956 27804 8968
rect 27571 8928 27804 8956
rect 27571 8925 27583 8928
rect 27525 8919 27583 8925
rect 27798 8916 27804 8928
rect 27856 8916 27862 8968
rect 35866 8956 35894 9064
rect 50338 8956 50344 8968
rect 35866 8928 50344 8956
rect 50338 8916 50344 8928
rect 50396 8916 50402 8968
rect 50430 8916 50436 8968
rect 50488 8956 50494 8968
rect 57885 8959 57943 8965
rect 57885 8956 57897 8959
rect 50488 8928 57897 8956
rect 50488 8916 50494 8928
rect 57885 8925 57897 8928
rect 57931 8925 57943 8959
rect 57885 8919 57943 8925
rect 26510 8888 26516 8900
rect 26471 8860 26516 8888
rect 26510 8848 26516 8860
rect 26568 8848 26574 8900
rect 22189 8823 22247 8829
rect 22189 8789 22201 8823
rect 22235 8820 22247 8823
rect 22462 8820 22468 8832
rect 22235 8792 22468 8820
rect 22235 8789 22247 8792
rect 22189 8783 22247 8789
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 22646 8820 22652 8832
rect 22607 8792 22652 8820
rect 22646 8780 22652 8792
rect 22704 8780 22710 8832
rect 27614 8780 27620 8832
rect 27672 8820 27678 8832
rect 58066 8820 58072 8832
rect 27672 8792 27717 8820
rect 58027 8792 58072 8820
rect 27672 8780 27678 8792
rect 58066 8780 58072 8792
rect 58124 8780 58130 8832
rect 1104 8730 58880 8752
rect 1104 8678 20214 8730
rect 20266 8678 20278 8730
rect 20330 8678 20342 8730
rect 20394 8678 20406 8730
rect 20458 8678 20470 8730
rect 20522 8678 39478 8730
rect 39530 8678 39542 8730
rect 39594 8678 39606 8730
rect 39658 8678 39670 8730
rect 39722 8678 39734 8730
rect 39786 8678 58880 8730
rect 1104 8656 58880 8678
rect 9398 8576 9404 8628
rect 9456 8616 9462 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9456 8588 9505 8616
rect 9456 8576 9462 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 23198 8616 23204 8628
rect 23159 8588 23204 8616
rect 9493 8579 9551 8585
rect 23198 8576 23204 8588
rect 23256 8576 23262 8628
rect 23566 8616 23572 8628
rect 23527 8588 23572 8616
rect 23566 8576 23572 8588
rect 23624 8576 23630 8628
rect 57425 8619 57483 8625
rect 57425 8616 57437 8619
rect 23768 8588 57437 8616
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8480 9735 8483
rect 9858 8480 9864 8492
rect 9723 8452 9864 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 15102 8480 15108 8492
rect 13679 8452 15108 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 15102 8440 15108 8452
rect 15160 8440 15166 8492
rect 22462 8480 22468 8492
rect 22423 8452 22468 8480
rect 22462 8440 22468 8452
rect 22520 8440 22526 8492
rect 23768 8480 23796 8588
rect 57425 8585 57437 8588
rect 57471 8585 57483 8619
rect 57425 8579 57483 8585
rect 50430 8548 50436 8560
rect 23492 8452 23796 8480
rect 31726 8520 50436 8548
rect 20990 8372 20996 8424
rect 21048 8412 21054 8424
rect 23492 8412 23520 8452
rect 23658 8412 23664 8424
rect 21048 8384 23520 8412
rect 23619 8384 23664 8412
rect 21048 8372 21054 8384
rect 23658 8372 23664 8384
rect 23716 8372 23722 8424
rect 23750 8372 23756 8424
rect 23808 8412 23814 8424
rect 23808 8384 23853 8412
rect 23808 8372 23814 8384
rect 22649 8347 22707 8353
rect 22649 8313 22661 8347
rect 22695 8344 22707 8347
rect 31726 8344 31754 8520
rect 50430 8508 50436 8520
rect 50488 8508 50494 8560
rect 57440 8480 57468 8579
rect 57885 8483 57943 8489
rect 57885 8480 57897 8483
rect 57440 8452 57897 8480
rect 57885 8449 57897 8452
rect 57931 8449 57943 8483
rect 57885 8443 57943 8449
rect 22695 8316 31754 8344
rect 22695 8313 22707 8316
rect 22649 8307 22707 8313
rect 57882 8304 57888 8356
rect 57940 8344 57946 8356
rect 58069 8347 58127 8353
rect 58069 8344 58081 8347
rect 57940 8316 58081 8344
rect 57940 8304 57946 8316
rect 58069 8313 58081 8316
rect 58115 8313 58127 8347
rect 58069 8307 58127 8313
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 13449 8279 13507 8285
rect 13449 8276 13461 8279
rect 13044 8248 13461 8276
rect 13044 8236 13050 8248
rect 13449 8245 13461 8248
rect 13495 8245 13507 8279
rect 13449 8239 13507 8245
rect 1104 8186 58880 8208
rect 1104 8134 10582 8186
rect 10634 8134 10646 8186
rect 10698 8134 10710 8186
rect 10762 8134 10774 8186
rect 10826 8134 10838 8186
rect 10890 8134 29846 8186
rect 29898 8134 29910 8186
rect 29962 8134 29974 8186
rect 30026 8134 30038 8186
rect 30090 8134 30102 8186
rect 30154 8134 49110 8186
rect 49162 8134 49174 8186
rect 49226 8134 49238 8186
rect 49290 8134 49302 8186
rect 49354 8134 49366 8186
rect 49418 8134 58880 8186
rect 1104 8112 58880 8134
rect 9858 8072 9864 8084
rect 9819 8044 9864 8072
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 10962 8072 10968 8084
rect 10923 8044 10968 8072
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 12526 8072 12532 8084
rect 12487 8044 12532 8072
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 13449 8075 13507 8081
rect 13449 8041 13461 8075
rect 13495 8072 13507 8075
rect 14274 8072 14280 8084
rect 13495 8044 14280 8072
rect 13495 8041 13507 8044
rect 13449 8035 13507 8041
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 20990 8072 20996 8084
rect 20951 8044 20996 8072
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 9769 8007 9827 8013
rect 9769 7973 9781 8007
rect 9815 7973 9827 8007
rect 9769 7967 9827 7973
rect 10229 8007 10287 8013
rect 10229 7973 10241 8007
rect 10275 8004 10287 8007
rect 10870 8004 10876 8016
rect 10275 7976 10876 8004
rect 10275 7973 10287 7976
rect 10229 7967 10287 7973
rect 9784 7936 9812 7967
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 12342 8004 12348 8016
rect 12303 7976 12348 8004
rect 12342 7964 12348 7976
rect 12400 7964 12406 8016
rect 13354 8004 13360 8016
rect 13315 7976 13360 8004
rect 13354 7964 13360 7976
rect 13412 7964 13418 8016
rect 9858 7936 9864 7948
rect 9784 7908 9864 7936
rect 9858 7896 9864 7908
rect 9916 7896 9922 7948
rect 10505 7939 10563 7945
rect 10505 7905 10517 7939
rect 10551 7936 10563 7939
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 10551 7908 12081 7936
rect 10551 7905 10563 7908
rect 10505 7899 10563 7905
rect 12069 7905 12081 7908
rect 12115 7936 12127 7939
rect 12986 7936 12992 7948
rect 12115 7908 12992 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 9398 7868 9404 7880
rect 9311 7840 9404 7868
rect 9398 7828 9404 7840
rect 9456 7868 9462 7880
rect 10520 7868 10548 7899
rect 12986 7896 12992 7908
rect 13044 7896 13050 7948
rect 20806 7868 20812 7880
rect 9456 7840 10548 7868
rect 20767 7840 20812 7868
rect 9456 7828 9462 7840
rect 20806 7828 20812 7840
rect 20864 7828 20870 7880
rect 57885 7871 57943 7877
rect 57885 7868 57897 7871
rect 57532 7840 57897 7868
rect 15102 7760 15108 7812
rect 15160 7800 15166 7812
rect 19889 7803 19947 7809
rect 19889 7800 19901 7803
rect 15160 7772 19901 7800
rect 15160 7760 15166 7772
rect 19889 7769 19901 7772
rect 19935 7800 19947 7803
rect 26510 7800 26516 7812
rect 19935 7772 26516 7800
rect 19935 7769 19947 7772
rect 19889 7763 19947 7769
rect 26510 7760 26516 7772
rect 26568 7760 26574 7812
rect 57532 7744 57560 7840
rect 57885 7837 57897 7840
rect 57931 7837 57943 7871
rect 57885 7831 57943 7837
rect 19978 7732 19984 7744
rect 19939 7704 19984 7732
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 57514 7732 57520 7744
rect 57475 7704 57520 7732
rect 57514 7692 57520 7704
rect 57572 7692 57578 7744
rect 58066 7732 58072 7744
rect 58027 7704 58072 7732
rect 58066 7692 58072 7704
rect 58124 7692 58130 7744
rect 1104 7642 58880 7664
rect 1104 7590 20214 7642
rect 20266 7590 20278 7642
rect 20330 7590 20342 7642
rect 20394 7590 20406 7642
rect 20458 7590 20470 7642
rect 20522 7590 39478 7642
rect 39530 7590 39542 7642
rect 39594 7590 39606 7642
rect 39658 7590 39670 7642
rect 39722 7590 39734 7642
rect 39786 7590 58880 7642
rect 1104 7568 58880 7590
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 9824 7500 9873 7528
rect 9824 7488 9830 7500
rect 9861 7497 9873 7500
rect 9907 7497 9919 7531
rect 9861 7491 9919 7497
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 57974 7528 57980 7540
rect 10928 7500 57980 7528
rect 10928 7488 10934 7500
rect 57974 7488 57980 7500
rect 58032 7488 58038 7540
rect 9398 7460 9404 7472
rect 9359 7432 9404 7460
rect 9398 7420 9404 7432
rect 9456 7420 9462 7472
rect 19242 7420 19248 7472
rect 19300 7460 19306 7472
rect 19337 7463 19395 7469
rect 19337 7460 19349 7463
rect 19300 7432 19349 7460
rect 19300 7420 19306 7432
rect 19337 7429 19349 7432
rect 19383 7429 19395 7463
rect 19337 7423 19395 7429
rect 20070 7420 20076 7472
rect 20128 7460 20134 7472
rect 20533 7463 20591 7469
rect 20533 7460 20545 7463
rect 20128 7432 20545 7460
rect 20128 7420 20134 7432
rect 20533 7429 20545 7432
rect 20579 7429 20591 7463
rect 20533 7423 20591 7429
rect 20625 7463 20683 7469
rect 20625 7429 20637 7463
rect 20671 7460 20683 7463
rect 20714 7460 20720 7472
rect 20671 7432 20720 7460
rect 20671 7429 20683 7432
rect 20625 7423 20683 7429
rect 20714 7420 20720 7432
rect 20772 7420 20778 7472
rect 57422 7352 57428 7404
rect 57480 7392 57486 7404
rect 57885 7395 57943 7401
rect 57885 7392 57897 7395
rect 57480 7364 57897 7392
rect 57480 7352 57486 7364
rect 57885 7361 57897 7364
rect 57931 7361 57943 7395
rect 57885 7355 57943 7361
rect 19242 7284 19248 7336
rect 19300 7324 19306 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 19300 7296 19441 7324
rect 19300 7284 19306 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 19521 7327 19579 7333
rect 19521 7293 19533 7327
rect 19567 7324 19579 7327
rect 19978 7324 19984 7336
rect 19567 7296 19984 7324
rect 19567 7293 19579 7296
rect 19521 7287 19579 7293
rect 9766 7256 9772 7268
rect 9727 7228 9772 7256
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 17770 7216 17776 7268
rect 17828 7256 17834 7268
rect 19536 7256 19564 7287
rect 19978 7284 19984 7296
rect 20036 7324 20042 7336
rect 20717 7327 20775 7333
rect 20717 7324 20729 7327
rect 20036 7296 20729 7324
rect 20036 7284 20042 7296
rect 20717 7293 20729 7296
rect 20763 7293 20775 7327
rect 20717 7287 20775 7293
rect 17828 7228 19564 7256
rect 20165 7259 20223 7265
rect 17828 7216 17834 7228
rect 20165 7225 20177 7259
rect 20211 7256 20223 7259
rect 20806 7256 20812 7268
rect 20211 7228 20812 7256
rect 20211 7225 20223 7228
rect 20165 7219 20223 7225
rect 20806 7216 20812 7228
rect 20864 7216 20870 7268
rect 18969 7191 19027 7197
rect 18969 7157 18981 7191
rect 19015 7188 19027 7191
rect 19610 7188 19616 7200
rect 19015 7160 19616 7188
rect 19015 7157 19027 7160
rect 18969 7151 19027 7157
rect 19610 7148 19616 7160
rect 19668 7148 19674 7200
rect 57422 7188 57428 7200
rect 57383 7160 57428 7188
rect 57422 7148 57428 7160
rect 57480 7148 57486 7200
rect 58066 7188 58072 7200
rect 58027 7160 58072 7188
rect 58066 7148 58072 7160
rect 58124 7148 58130 7200
rect 1104 7098 58880 7120
rect 1104 7046 10582 7098
rect 10634 7046 10646 7098
rect 10698 7046 10710 7098
rect 10762 7046 10774 7098
rect 10826 7046 10838 7098
rect 10890 7046 29846 7098
rect 29898 7046 29910 7098
rect 29962 7046 29974 7098
rect 30026 7046 30038 7098
rect 30090 7046 30102 7098
rect 30154 7046 49110 7098
rect 49162 7046 49174 7098
rect 49226 7046 49238 7098
rect 49290 7046 49302 7098
rect 49354 7046 49366 7098
rect 49418 7046 58880 7098
rect 1104 7024 58880 7046
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16632 6820 16681 6848
rect 16632 6808 16638 6820
rect 16669 6817 16681 6820
rect 16715 6848 16727 6851
rect 17770 6848 17776 6860
rect 16715 6820 17776 6848
rect 16715 6817 16727 6820
rect 16669 6811 16727 6817
rect 17770 6808 17776 6820
rect 17828 6848 17834 6860
rect 18049 6851 18107 6857
rect 18049 6848 18061 6851
rect 17828 6820 18061 6848
rect 17828 6808 17834 6820
rect 18049 6817 18061 6820
rect 18095 6817 18107 6851
rect 18049 6811 18107 6817
rect 16390 6780 16396 6792
rect 16351 6752 16396 6780
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 17862 6780 17868 6792
rect 17823 6752 17868 6780
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 19610 6780 19616 6792
rect 19571 6752 19616 6780
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 50338 6740 50344 6792
rect 50396 6780 50402 6792
rect 57885 6783 57943 6789
rect 57885 6780 57897 6783
rect 50396 6752 57897 6780
rect 50396 6740 50402 6752
rect 57885 6749 57897 6752
rect 57931 6749 57943 6783
rect 57885 6743 57943 6749
rect 16022 6644 16028 6656
rect 15983 6616 16028 6644
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6644 16543 6647
rect 16666 6644 16672 6656
rect 16531 6616 16672 6644
rect 16531 6613 16543 6616
rect 16485 6607 16543 6613
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 17494 6644 17500 6656
rect 17455 6616 17500 6644
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 17957 6647 18015 6653
rect 17957 6644 17969 6647
rect 17920 6616 17969 6644
rect 17920 6604 17926 6616
rect 17957 6613 17969 6616
rect 18003 6613 18015 6647
rect 17957 6607 18015 6613
rect 19797 6647 19855 6653
rect 19797 6613 19809 6647
rect 19843 6644 19855 6647
rect 57514 6644 57520 6656
rect 19843 6616 57520 6644
rect 19843 6613 19855 6616
rect 19797 6607 19855 6613
rect 57514 6604 57520 6616
rect 57572 6604 57578 6656
rect 58066 6644 58072 6656
rect 58027 6616 58072 6644
rect 58066 6604 58072 6616
rect 58124 6604 58130 6656
rect 1104 6554 58880 6576
rect 1104 6502 20214 6554
rect 20266 6502 20278 6554
rect 20330 6502 20342 6554
rect 20394 6502 20406 6554
rect 20458 6502 20470 6554
rect 20522 6502 39478 6554
rect 39530 6502 39542 6554
rect 39594 6502 39606 6554
rect 39658 6502 39670 6554
rect 39722 6502 39734 6554
rect 39786 6502 58880 6554
rect 1104 6480 58880 6502
rect 15010 6400 15016 6452
rect 15068 6440 15074 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15068 6412 15577 6440
rect 15068 6400 15074 6412
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 18417 6443 18475 6449
rect 18417 6409 18429 6443
rect 18463 6440 18475 6443
rect 18463 6412 31754 6440
rect 18463 6409 18475 6412
rect 18417 6403 18475 6409
rect 16022 6332 16028 6384
rect 16080 6372 16086 6384
rect 16080 6344 17448 6372
rect 16080 6332 16086 6344
rect 17420 6313 17448 6344
rect 16669 6307 16727 6313
rect 16669 6273 16681 6307
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 17405 6307 17463 6313
rect 17405 6273 17417 6307
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 15654 6236 15660 6248
rect 15615 6208 15660 6236
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16574 6236 16580 6248
rect 15887 6208 16580 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 15197 6171 15255 6177
rect 15197 6137 15209 6171
rect 15243 6168 15255 6171
rect 16684 6168 16712 6267
rect 17494 6264 17500 6316
rect 17552 6304 17558 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 17552 6276 18245 6304
rect 17552 6264 17558 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 31726 6236 31754 6412
rect 57885 6307 57943 6313
rect 57885 6273 57897 6307
rect 57931 6273 57943 6307
rect 57885 6267 57943 6273
rect 57422 6236 57428 6248
rect 16868 6208 26924 6236
rect 31726 6208 57428 6236
rect 16868 6177 16896 6208
rect 15243 6140 16712 6168
rect 16853 6171 16911 6177
rect 15243 6137 15255 6140
rect 15197 6131 15255 6137
rect 16853 6137 16865 6171
rect 16899 6137 16911 6171
rect 16853 6131 16911 6137
rect 17589 6171 17647 6177
rect 17589 6137 17601 6171
rect 17635 6168 17647 6171
rect 26896 6168 26924 6208
rect 57422 6196 57428 6208
rect 57480 6196 57486 6248
rect 57900 6168 57928 6267
rect 17635 6140 22048 6168
rect 26896 6140 57928 6168
rect 17635 6137 17647 6140
rect 17589 6131 17647 6137
rect 22020 6100 22048 6140
rect 50338 6100 50344 6112
rect 22020 6072 50344 6100
rect 50338 6060 50344 6072
rect 50396 6060 50402 6112
rect 58066 6100 58072 6112
rect 58027 6072 58072 6100
rect 58066 6060 58072 6072
rect 58124 6060 58130 6112
rect 1104 6010 58880 6032
rect 1104 5958 10582 6010
rect 10634 5958 10646 6010
rect 10698 5958 10710 6010
rect 10762 5958 10774 6010
rect 10826 5958 10838 6010
rect 10890 5958 29846 6010
rect 29898 5958 29910 6010
rect 29962 5958 29974 6010
rect 30026 5958 30038 6010
rect 30090 5958 30102 6010
rect 30154 5958 49110 6010
rect 49162 5958 49174 6010
rect 49226 5958 49238 6010
rect 49290 5958 49302 6010
rect 49354 5958 49366 6010
rect 49418 5958 58880 6010
rect 1104 5936 58880 5958
rect 55766 5856 55772 5908
rect 55824 5896 55830 5908
rect 56965 5899 57023 5905
rect 56965 5896 56977 5899
rect 55824 5868 56977 5896
rect 55824 5856 55830 5868
rect 56965 5865 56977 5868
rect 57011 5865 57023 5899
rect 56965 5859 57023 5865
rect 57974 5828 57980 5840
rect 57935 5800 57980 5828
rect 57974 5788 57980 5800
rect 58032 5788 58038 5840
rect 56870 5624 56876 5636
rect 56831 5596 56876 5624
rect 56870 5584 56876 5596
rect 56928 5584 56934 5636
rect 57790 5624 57796 5636
rect 57751 5596 57796 5624
rect 57790 5584 57796 5596
rect 57848 5584 57854 5636
rect 1104 5466 58880 5488
rect 1104 5414 20214 5466
rect 20266 5414 20278 5466
rect 20330 5414 20342 5466
rect 20394 5414 20406 5466
rect 20458 5414 20470 5466
rect 20522 5414 39478 5466
rect 39530 5414 39542 5466
rect 39594 5414 39606 5466
rect 39658 5414 39670 5466
rect 39722 5414 39734 5466
rect 39786 5414 58880 5466
rect 1104 5392 58880 5414
rect 56502 5176 56508 5228
rect 56560 5216 56566 5228
rect 56965 5219 57023 5225
rect 56965 5216 56977 5219
rect 56560 5188 56977 5216
rect 56560 5176 56566 5188
rect 56965 5185 56977 5188
rect 57011 5185 57023 5219
rect 56965 5179 57023 5185
rect 56778 4972 56784 5024
rect 56836 5012 56842 5024
rect 57057 5015 57115 5021
rect 57057 5012 57069 5015
rect 56836 4984 57069 5012
rect 56836 4972 56842 4984
rect 57057 4981 57069 4984
rect 57103 4981 57115 5015
rect 57057 4975 57115 4981
rect 1104 4922 58880 4944
rect 1104 4870 10582 4922
rect 10634 4870 10646 4922
rect 10698 4870 10710 4922
rect 10762 4870 10774 4922
rect 10826 4870 10838 4922
rect 10890 4870 29846 4922
rect 29898 4870 29910 4922
rect 29962 4870 29974 4922
rect 30026 4870 30038 4922
rect 30090 4870 30102 4922
rect 30154 4870 49110 4922
rect 49162 4870 49174 4922
rect 49226 4870 49238 4922
rect 49290 4870 49302 4922
rect 49354 4870 49366 4922
rect 49418 4870 58880 4922
rect 1104 4848 58880 4870
rect 57606 4672 57612 4684
rect 57567 4644 57612 4672
rect 57606 4632 57612 4644
rect 57664 4632 57670 4684
rect 57333 4607 57391 4613
rect 57333 4573 57345 4607
rect 57379 4604 57391 4607
rect 59170 4604 59176 4616
rect 57379 4576 59176 4604
rect 57379 4573 57391 4576
rect 57333 4567 57391 4573
rect 59170 4564 59176 4576
rect 59228 4564 59234 4616
rect 56502 4536 56508 4548
rect 56463 4508 56508 4536
rect 56502 4496 56508 4508
rect 56560 4496 56566 4548
rect 56594 4468 56600 4480
rect 56555 4440 56600 4468
rect 56594 4428 56600 4440
rect 56652 4428 56658 4480
rect 1104 4378 58880 4400
rect 1104 4326 20214 4378
rect 20266 4326 20278 4378
rect 20330 4326 20342 4378
rect 20394 4326 20406 4378
rect 20458 4326 20470 4378
rect 20522 4326 39478 4378
rect 39530 4326 39542 4378
rect 39594 4326 39606 4378
rect 39658 4326 39670 4378
rect 39722 4326 39734 4378
rect 39786 4326 58880 4378
rect 1104 4304 58880 4326
rect 56042 4196 56048 4208
rect 56003 4168 56048 4196
rect 56042 4156 56048 4168
rect 56100 4156 56106 4208
rect 56965 4199 57023 4205
rect 56965 4165 56977 4199
rect 57011 4196 57023 4199
rect 57146 4196 57152 4208
rect 57011 4168 57152 4196
rect 57011 4165 57023 4168
rect 56965 4159 57023 4165
rect 57146 4156 57152 4168
rect 57204 4156 57210 4208
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 2188 4100 3249 4128
rect 2188 4088 2194 4100
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3786 4088 3792 4140
rect 3844 4128 3850 4140
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 3844 4100 4537 4128
rect 3844 4088 3850 4100
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 6641 4131 6699 4137
rect 6641 4128 6653 4131
rect 6604 4100 6653 4128
rect 6604 4088 6610 4100
rect 6641 4097 6653 4100
rect 6687 4097 6699 4131
rect 7926 4128 7932 4140
rect 7887 4100 7932 4128
rect 6641 4091 6699 4097
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 2958 4060 2964 4072
rect 2919 4032 2964 4060
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3970 4020 3976 4072
rect 4028 4060 4034 4072
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4028 4032 4261 4060
rect 4028 4020 4034 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 6365 4063 6423 4069
rect 6365 4029 6377 4063
rect 6411 4060 6423 4063
rect 6822 4060 6828 4072
rect 6411 4032 6828 4060
rect 6411 4029 6423 4032
rect 6365 4023 6423 4029
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 7282 4020 7288 4072
rect 7340 4060 7346 4072
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 7340 4032 7665 4060
rect 7340 4020 7346 4032
rect 7653 4029 7665 4032
rect 7699 4029 7711 4063
rect 7653 4023 7711 4029
rect 9858 3952 9864 4004
rect 9916 3992 9922 4004
rect 56229 3995 56287 4001
rect 56229 3992 56241 3995
rect 9916 3964 56241 3992
rect 9916 3952 9922 3964
rect 56229 3961 56241 3964
rect 56275 3961 56287 3995
rect 56229 3955 56287 3961
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 55674 3924 55680 3936
rect 6788 3896 55680 3924
rect 6788 3884 6794 3896
rect 55674 3884 55680 3896
rect 55732 3884 55738 3936
rect 57054 3924 57060 3936
rect 57015 3896 57060 3924
rect 57054 3884 57060 3896
rect 57112 3884 57118 3936
rect 1104 3834 58880 3856
rect 1104 3782 10582 3834
rect 10634 3782 10646 3834
rect 10698 3782 10710 3834
rect 10762 3782 10774 3834
rect 10826 3782 10838 3834
rect 10890 3782 29846 3834
rect 29898 3782 29910 3834
rect 29962 3782 29974 3834
rect 30026 3782 30038 3834
rect 30090 3782 30102 3834
rect 30154 3782 49110 3834
rect 49162 3782 49174 3834
rect 49226 3782 49238 3834
rect 49290 3782 49302 3834
rect 49354 3782 49366 3834
rect 49418 3782 58880 3834
rect 1104 3760 58880 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 4249 3723 4307 3729
rect 4249 3720 4261 3723
rect 3016 3692 4261 3720
rect 3016 3680 3022 3692
rect 4249 3689 4261 3692
rect 4295 3689 4307 3723
rect 56597 3723 56655 3729
rect 56597 3720 56609 3723
rect 4249 3683 4307 3689
rect 6886 3692 56609 3720
rect 4062 3652 4068 3664
rect 4023 3624 4068 3652
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 6886 3652 6914 3692
rect 56597 3689 56609 3692
rect 56643 3689 56655 3723
rect 56597 3683 56655 3689
rect 4172 3624 6914 3652
rect 7193 3655 7251 3661
rect 3878 3544 3884 3596
rect 3936 3584 3942 3596
rect 4172 3584 4200 3624
rect 7193 3621 7205 3655
rect 7239 3652 7251 3655
rect 7466 3652 7472 3664
rect 7239 3624 7472 3652
rect 7239 3621 7251 3624
rect 7193 3615 7251 3621
rect 7466 3612 7472 3624
rect 7524 3652 7530 3664
rect 55769 3655 55827 3661
rect 55769 3652 55781 3655
rect 7524 3624 55781 3652
rect 7524 3612 7530 3624
rect 55769 3621 55781 3624
rect 55815 3621 55827 3655
rect 55769 3615 55827 3621
rect 5074 3584 5080 3596
rect 3936 3556 4200 3584
rect 5035 3556 5080 3584
rect 3936 3544 3942 3556
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 57054 3584 57060 3596
rect 5408 3556 7144 3584
rect 5408 3544 5414 3556
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 4154 3516 4160 3528
rect 3283 3488 4160 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 4982 3516 4988 3528
rect 4847 3488 4988 3516
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3516 6423 3519
rect 7116 3516 7144 3556
rect 7300 3556 57060 3584
rect 7300 3516 7328 3556
rect 57054 3544 57060 3556
rect 57112 3544 57118 3596
rect 57333 3587 57391 3593
rect 57333 3553 57345 3587
rect 57379 3584 57391 3587
rect 57698 3584 57704 3596
rect 57379 3556 57704 3584
rect 57379 3553 57391 3556
rect 57333 3547 57391 3553
rect 57698 3544 57704 3556
rect 57756 3544 57762 3596
rect 6411 3488 6960 3516
rect 7116 3488 7328 3516
rect 6411 3485 6423 3488
rect 6365 3479 6423 3485
rect 3786 3448 3792 3460
rect 3747 3420 3792 3448
rect 3786 3408 3792 3420
rect 3844 3408 3850 3460
rect 6825 3451 6883 3457
rect 6825 3448 6837 3451
rect 6196 3420 6837 3448
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 6196 3389 6224 3420
rect 6825 3417 6837 3420
rect 6871 3417 6883 3451
rect 6932 3448 6960 3488
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 7929 3519 7987 3525
rect 7929 3516 7941 3519
rect 7708 3488 7941 3516
rect 7708 3476 7714 3488
rect 7929 3485 7941 3488
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9950 3516 9956 3528
rect 9355 3488 9956 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9950 3476 9956 3488
rect 10008 3476 10014 3528
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 8386 3448 8392 3460
rect 6932 3420 8392 3448
rect 6825 3411 6883 3417
rect 8386 3408 8392 3420
rect 8444 3448 8450 3460
rect 10888 3448 10916 3479
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 11517 3519 11575 3525
rect 11517 3516 11529 3519
rect 11020 3488 11529 3516
rect 11020 3476 11026 3488
rect 11517 3485 11529 3488
rect 11563 3485 11575 3519
rect 40126 3516 40132 3528
rect 11517 3479 11575 3485
rect 16546 3488 40132 3516
rect 16546 3448 16574 3488
rect 40126 3476 40132 3488
rect 40184 3476 40190 3528
rect 56962 3476 56968 3528
rect 57020 3516 57026 3528
rect 57609 3519 57667 3525
rect 57609 3516 57621 3519
rect 57020 3488 57621 3516
rect 57020 3476 57026 3488
rect 57609 3485 57621 3488
rect 57655 3485 57667 3519
rect 57609 3479 57667 3485
rect 8444 3420 16574 3448
rect 55585 3451 55643 3457
rect 8444 3408 8450 3420
rect 55585 3417 55597 3451
rect 55631 3448 55643 3451
rect 55766 3448 55772 3460
rect 55631 3420 55772 3448
rect 55631 3417 55643 3420
rect 55585 3411 55643 3417
rect 55766 3408 55772 3420
rect 55824 3408 55830 3460
rect 56502 3448 56508 3460
rect 56463 3420 56508 3448
rect 56502 3408 56508 3420
rect 56560 3408 56566 3460
rect 3053 3383 3111 3389
rect 3053 3380 3065 3383
rect 2832 3352 3065 3380
rect 2832 3340 2838 3352
rect 3053 3349 3065 3352
rect 3099 3349 3111 3383
rect 3053 3343 3111 3349
rect 6181 3383 6239 3389
rect 6181 3349 6193 3383
rect 6227 3380 6239 3383
rect 6362 3380 6368 3392
rect 6227 3352 6368 3380
rect 6227 3349 6239 3352
rect 6181 3343 6239 3349
rect 6362 3340 6368 3352
rect 6420 3340 6426 3392
rect 7282 3380 7288 3392
rect 7243 3352 7288 3380
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7745 3383 7803 3389
rect 7745 3349 7757 3383
rect 7791 3380 7803 3383
rect 7926 3380 7932 3392
rect 7791 3352 7932 3380
rect 7791 3349 7803 3352
rect 7745 3343 7803 3349
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 9122 3380 9128 3392
rect 9083 3352 9128 3380
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 10689 3383 10747 3389
rect 10689 3349 10701 3383
rect 10735 3380 10747 3383
rect 10778 3380 10784 3392
rect 10735 3352 10784 3380
rect 10735 3349 10747 3352
rect 10689 3343 10747 3349
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 11333 3383 11391 3389
rect 11333 3349 11345 3383
rect 11379 3380 11391 3383
rect 11514 3380 11520 3392
rect 11379 3352 11520 3380
rect 11379 3349 11391 3352
rect 11333 3343 11391 3349
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 48406 3340 48412 3392
rect 48464 3380 48470 3392
rect 56778 3380 56784 3392
rect 48464 3352 56784 3380
rect 48464 3340 48470 3352
rect 56778 3340 56784 3352
rect 56836 3340 56842 3392
rect 1104 3290 58880 3312
rect 1104 3238 20214 3290
rect 20266 3238 20278 3290
rect 20330 3238 20342 3290
rect 20394 3238 20406 3290
rect 20458 3238 20470 3290
rect 20522 3238 39478 3290
rect 39530 3238 39542 3290
rect 39594 3238 39606 3290
rect 39658 3238 39670 3290
rect 39722 3238 39734 3290
rect 39786 3238 58880 3290
rect 1104 3216 58880 3238
rect 3970 3176 3976 3188
rect 3931 3148 3976 3176
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 4982 3176 4988 3188
rect 4943 3148 4988 3176
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 6822 3176 6828 3188
rect 5224 3148 6500 3176
rect 6783 3148 6828 3176
rect 5224 3136 5230 3148
rect 3234 3108 3240 3120
rect 2332 3080 3240 3108
rect 2332 3049 2360 3080
rect 3234 3068 3240 3080
rect 3292 3068 3298 3120
rect 3513 3111 3571 3117
rect 3513 3077 3525 3111
rect 3559 3108 3571 3111
rect 3786 3108 3792 3120
rect 3559 3080 3792 3108
rect 3559 3077 3571 3080
rect 3513 3071 3571 3077
rect 3786 3068 3792 3080
rect 3844 3108 3850 3120
rect 4525 3111 4583 3117
rect 4525 3108 4537 3111
rect 3844 3080 4537 3108
rect 3844 3068 3850 3080
rect 4525 3077 4537 3080
rect 4571 3108 4583 3111
rect 6362 3108 6368 3120
rect 4571 3080 6368 3108
rect 4571 3077 4583 3080
rect 4525 3071 4583 3077
rect 6362 3068 6368 3080
rect 6420 3068 6426 3120
rect 6472 3108 6500 3148
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7650 3176 7656 3188
rect 7611 3148 7656 3176
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 10873 3179 10931 3185
rect 10873 3145 10885 3179
rect 10919 3176 10931 3179
rect 10962 3176 10968 3188
rect 10919 3148 10968 3176
rect 10919 3145 10931 3148
rect 10873 3139 10931 3145
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 13412 3148 13553 3176
rect 13412 3136 13418 3148
rect 13541 3145 13553 3148
rect 13587 3176 13599 3179
rect 48406 3176 48412 3188
rect 13587 3148 48412 3176
rect 13587 3145 13599 3148
rect 13541 3139 13599 3145
rect 48406 3136 48412 3148
rect 48464 3136 48470 3188
rect 55674 3176 55680 3188
rect 55635 3148 55680 3176
rect 55674 3136 55680 3148
rect 55732 3136 55738 3188
rect 9122 3108 9128 3120
rect 6472 3080 9128 3108
rect 9122 3068 9128 3080
rect 9180 3068 9186 3120
rect 10045 3111 10103 3117
rect 10045 3108 10057 3111
rect 9232 3080 10057 3108
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 5626 3040 5632 3052
rect 5587 3012 5632 3040
rect 2777 3003 2835 3009
rect 2792 2972 2820 3003
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 7466 3040 7472 3052
rect 7427 3012 7472 3040
rect 7466 3000 7472 3012
rect 7524 3000 7530 3052
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 8386 3040 8392 3052
rect 8343 3012 8392 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 9232 3049 9260 3080
rect 10045 3077 10057 3080
rect 10091 3077 10103 3111
rect 13372 3108 13400 3136
rect 56594 3108 56600 3120
rect 10045 3071 10103 3077
rect 13096 3080 13400 3108
rect 16546 3080 56600 3108
rect 9217 3043 9275 3049
rect 9217 3009 9229 3043
rect 9263 3009 9275 3043
rect 9858 3040 9864 3052
rect 9819 3012 9864 3040
rect 9217 3003 9275 3009
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3040 10747 3043
rect 10870 3040 10876 3052
rect 10735 3012 10876 3040
rect 10735 3009 10747 3012
rect 10689 3003 10747 3009
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3040 11851 3043
rect 12253 3043 12311 3049
rect 12253 3040 12265 3043
rect 11839 3012 12265 3040
rect 11839 3009 11851 3012
rect 11793 3003 11851 3009
rect 12253 3009 12265 3012
rect 12299 3040 12311 3043
rect 12342 3040 12348 3052
rect 12299 3012 12348 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 12342 3000 12348 3012
rect 12400 3040 12406 3052
rect 13096 3049 13124 3080
rect 13081 3043 13139 3049
rect 12400 3012 13032 3040
rect 12400 3000 12406 3012
rect 2148 2944 2820 2972
rect 2148 2913 2176 2944
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 7156 2944 7297 2972
rect 7156 2932 7162 2944
rect 7285 2941 7297 2944
rect 7331 2972 7343 2975
rect 9674 2972 9680 2984
rect 7331 2944 8156 2972
rect 9587 2944 9680 2972
rect 7331 2941 7343 2944
rect 7285 2935 7343 2941
rect 2133 2907 2191 2913
rect 2133 2873 2145 2907
rect 2179 2873 2191 2907
rect 3878 2904 3884 2916
rect 3839 2876 3884 2904
rect 2133 2867 2191 2873
rect 3878 2864 3884 2876
rect 3936 2864 3942 2916
rect 4890 2904 4896 2916
rect 4803 2876 4896 2904
rect 4890 2864 4896 2876
rect 4948 2904 4954 2916
rect 5350 2904 5356 2916
rect 4948 2876 5356 2904
rect 4948 2864 4954 2876
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 6730 2904 6736 2916
rect 6691 2876 6736 2904
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 8128 2913 8156 2944
rect 9674 2932 9680 2944
rect 9732 2972 9738 2984
rect 10505 2975 10563 2981
rect 10505 2972 10517 2975
rect 9732 2944 10517 2972
rect 9732 2932 9738 2944
rect 10505 2941 10517 2944
rect 10551 2972 10563 2975
rect 10778 2972 10784 2984
rect 10551 2944 10784 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 10778 2932 10784 2944
rect 10836 2972 10842 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 10836 2944 12081 2972
rect 10836 2932 10842 2944
rect 12069 2941 12081 2944
rect 12115 2972 12127 2975
rect 12897 2975 12955 2981
rect 12897 2972 12909 2975
rect 12115 2944 12909 2972
rect 12115 2941 12127 2944
rect 12069 2935 12127 2941
rect 12897 2941 12909 2944
rect 12943 2941 12955 2975
rect 13004 2972 13032 3012
rect 13081 3009 13093 3043
rect 13127 3009 13139 3043
rect 13081 3003 13139 3009
rect 13265 3043 13323 3049
rect 13265 3009 13277 3043
rect 13311 3040 13323 3043
rect 13909 3043 13967 3049
rect 13909 3040 13921 3043
rect 13311 3012 13921 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 13909 3009 13921 3012
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 16546 2972 16574 3080
rect 56594 3068 56600 3080
rect 56652 3068 56658 3120
rect 49510 3040 49516 3052
rect 49471 3012 49516 3040
rect 49510 3000 49516 3012
rect 49568 3000 49574 3052
rect 53834 3040 53840 3052
rect 53795 3012 53840 3040
rect 53834 3000 53840 3012
rect 53892 3000 53898 3052
rect 55582 3040 55588 3052
rect 55543 3012 55588 3040
rect 55582 3000 55588 3012
rect 55640 3000 55646 3052
rect 56686 3040 56692 3052
rect 56647 3012 56692 3040
rect 56686 3000 56692 3012
rect 56744 3000 56750 3052
rect 13004 2944 16574 2972
rect 12897 2935 12955 2941
rect 48958 2932 48964 2984
rect 49016 2972 49022 2984
rect 49237 2975 49295 2981
rect 49237 2972 49249 2975
rect 49016 2944 49249 2972
rect 49016 2932 49022 2944
rect 49237 2941 49249 2944
rect 49283 2941 49295 2975
rect 49237 2935 49295 2941
rect 53466 2932 53472 2984
rect 53524 2972 53530 2984
rect 53561 2975 53619 2981
rect 53561 2972 53573 2975
rect 53524 2944 53573 2972
rect 53524 2932 53530 2944
rect 53561 2941 53573 2944
rect 53607 2941 53619 2975
rect 53561 2935 53619 2941
rect 56318 2932 56324 2984
rect 56376 2972 56382 2984
rect 56413 2975 56471 2981
rect 56413 2972 56425 2975
rect 56376 2944 56425 2972
rect 56376 2932 56382 2944
rect 56413 2941 56425 2944
rect 56459 2941 56471 2975
rect 56413 2935 56471 2941
rect 8113 2907 8171 2913
rect 8113 2873 8125 2907
rect 8159 2873 8171 2907
rect 8113 2867 8171 2873
rect 2961 2839 3019 2845
rect 2961 2805 2973 2839
rect 3007 2836 3019 2839
rect 3510 2836 3516 2848
rect 3007 2808 3516 2836
rect 3007 2805 3019 2808
rect 2961 2799 3019 2805
rect 3510 2796 3516 2808
rect 3568 2796 3574 2848
rect 5445 2839 5503 2845
rect 5445 2805 5457 2839
rect 5491 2836 5503 2839
rect 5534 2836 5540 2848
rect 5491 2808 5540 2836
rect 5491 2805 5503 2808
rect 5445 2799 5503 2805
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2836 9091 2839
rect 10410 2836 10416 2848
rect 9079 2808 10416 2836
rect 9079 2805 9091 2808
rect 9033 2799 9091 2805
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 12437 2839 12495 2845
rect 12437 2805 12449 2839
rect 12483 2836 12495 2839
rect 13170 2836 13176 2848
rect 12483 2808 13176 2836
rect 12483 2805 12495 2808
rect 12437 2799 12495 2805
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13725 2839 13783 2845
rect 13725 2805 13737 2839
rect 13771 2836 13783 2839
rect 14090 2836 14096 2848
rect 13771 2808 14096 2836
rect 13771 2805 13783 2808
rect 13725 2799 13783 2805
rect 14090 2796 14096 2808
rect 14148 2796 14154 2848
rect 1104 2746 58880 2768
rect 1104 2694 10582 2746
rect 10634 2694 10646 2746
rect 10698 2694 10710 2746
rect 10762 2694 10774 2746
rect 10826 2694 10838 2746
rect 10890 2694 29846 2746
rect 29898 2694 29910 2746
rect 29962 2694 29974 2746
rect 30026 2694 30038 2746
rect 30090 2694 30102 2746
rect 30154 2694 49110 2746
rect 49162 2694 49174 2746
rect 49226 2694 49238 2746
rect 49290 2694 49302 2746
rect 49354 2694 49366 2746
rect 49418 2694 58880 2746
rect 1104 2672 58880 2694
rect 3234 2632 3240 2644
rect 3195 2604 3240 2632
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 4154 2632 4160 2644
rect 4115 2604 4160 2632
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 5077 2635 5135 2641
rect 5077 2601 5089 2635
rect 5123 2632 5135 2635
rect 5626 2632 5632 2644
rect 5123 2604 5632 2632
rect 5123 2601 5135 2604
rect 5077 2595 5135 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 16666 2632 16672 2644
rect 5736 2604 16574 2632
rect 16627 2604 16672 2632
rect 5166 2564 5172 2576
rect 1412 2536 5172 2564
rect 1412 2437 1440 2536
rect 5166 2524 5172 2536
rect 5224 2524 5230 2576
rect 4062 2496 4068 2508
rect 3975 2468 4068 2496
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2774 2428 2780 2440
rect 2179 2400 2780 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2397 3019 2431
rect 2961 2391 3019 2397
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2428 3111 2431
rect 3786 2428 3792 2440
rect 3099 2400 3792 2428
rect 3099 2397 3111 2400
rect 3053 2391 3111 2397
rect 2976 2360 3004 2391
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 3988 2437 4016 2468
rect 4062 2456 4068 2468
rect 4120 2496 4126 2508
rect 5736 2496 5764 2604
rect 6362 2524 6368 2576
rect 6420 2564 6426 2576
rect 7377 2567 7435 2573
rect 7377 2564 7389 2567
rect 6420 2536 7389 2564
rect 6420 2524 6426 2536
rect 7377 2533 7389 2536
rect 7423 2533 7435 2567
rect 7377 2527 7435 2533
rect 9214 2524 9220 2576
rect 9272 2564 9278 2576
rect 10597 2567 10655 2573
rect 10597 2564 10609 2567
rect 9272 2536 10609 2564
rect 9272 2524 9278 2536
rect 10597 2533 10609 2536
rect 10643 2533 10655 2567
rect 10597 2527 10655 2533
rect 12989 2567 13047 2573
rect 12989 2533 13001 2567
rect 13035 2533 13047 2567
rect 12989 2527 13047 2533
rect 15013 2567 15071 2573
rect 15013 2533 15025 2567
rect 15059 2564 15071 2567
rect 15654 2564 15660 2576
rect 15059 2536 15660 2564
rect 15059 2533 15071 2536
rect 15013 2527 15071 2533
rect 4120 2468 5764 2496
rect 6733 2499 6791 2505
rect 4120 2456 4126 2468
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 9585 2499 9643 2505
rect 6779 2468 9168 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2397 3939 2431
rect 3881 2391 3939 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 3896 2360 3924 2391
rect 4816 2360 4844 2391
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 5534 2428 5540 2440
rect 4948 2400 4993 2428
rect 5495 2400 5540 2428
rect 4948 2388 4954 2400
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2397 6515 2431
rect 6457 2391 6515 2397
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2428 6607 2431
rect 6638 2428 6644 2440
rect 6595 2400 6644 2428
rect 6595 2397 6607 2400
rect 6549 2391 6607 2397
rect 6472 2360 6500 2391
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7926 2428 7932 2440
rect 7887 2400 7932 2428
rect 7193 2391 7251 2397
rect 7098 2360 7104 2372
rect 2976 2332 7104 2360
rect 7098 2320 7104 2332
rect 7156 2320 7162 2372
rect 7208 2360 7236 2391
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 9140 2437 9168 2468
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 9674 2496 9680 2508
rect 9631 2468 9680 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 9950 2496 9956 2508
rect 9911 2468 9956 2496
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2397 9183 2431
rect 9766 2428 9772 2440
rect 9679 2400 9772 2428
rect 9125 2391 9183 2397
rect 9766 2388 9772 2400
rect 9824 2388 9830 2440
rect 10410 2428 10416 2440
rect 10371 2400 10416 2428
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 11514 2428 11520 2440
rect 11475 2400 11520 2428
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2428 12311 2431
rect 13004 2428 13032 2527
rect 15654 2524 15660 2536
rect 15712 2524 15718 2576
rect 16546 2564 16574 2604
rect 16666 2592 16672 2604
rect 16724 2592 16730 2644
rect 17862 2632 17868 2644
rect 17823 2604 17868 2632
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 19242 2632 19248 2644
rect 19203 2604 19248 2632
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 20714 2632 20720 2644
rect 20675 2604 20720 2632
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 22097 2635 22155 2641
rect 22097 2601 22109 2635
rect 22143 2632 22155 2635
rect 22646 2632 22652 2644
rect 22143 2604 22652 2632
rect 22143 2601 22155 2604
rect 22097 2595 22155 2601
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 23569 2635 23627 2641
rect 23569 2601 23581 2635
rect 23615 2632 23627 2635
rect 23658 2632 23664 2644
rect 23615 2604 23664 2632
rect 23615 2601 23627 2604
rect 23569 2595 23627 2601
rect 23658 2592 23664 2604
rect 23716 2592 23722 2644
rect 24949 2635 25007 2641
rect 24949 2601 24961 2635
rect 24995 2632 25007 2635
rect 25038 2632 25044 2644
rect 24995 2604 25044 2632
rect 24995 2601 25007 2604
rect 24949 2595 25007 2601
rect 25038 2592 25044 2604
rect 25096 2592 25102 2644
rect 26973 2635 27031 2641
rect 26973 2601 26985 2635
rect 27019 2632 27031 2635
rect 27430 2632 27436 2644
rect 27019 2604 27436 2632
rect 27019 2601 27031 2604
rect 26973 2595 27031 2601
rect 27430 2592 27436 2604
rect 27488 2592 27494 2644
rect 27614 2592 27620 2644
rect 27672 2632 27678 2644
rect 27801 2635 27859 2641
rect 27801 2632 27813 2635
rect 27672 2604 27813 2632
rect 27672 2592 27678 2604
rect 27801 2601 27813 2604
rect 27847 2601 27859 2635
rect 29546 2632 29552 2644
rect 29507 2604 29552 2632
rect 27801 2595 27859 2601
rect 29546 2592 29552 2604
rect 29604 2592 29610 2644
rect 30742 2632 30748 2644
rect 30703 2604 30748 2632
rect 30742 2592 30748 2604
rect 30800 2592 30806 2644
rect 32122 2632 32128 2644
rect 32083 2604 32128 2632
rect 32122 2592 32128 2604
rect 32180 2592 32186 2644
rect 33594 2632 33600 2644
rect 33555 2604 33600 2632
rect 33594 2592 33600 2604
rect 33652 2592 33658 2644
rect 34974 2632 34980 2644
rect 34935 2604 34980 2632
rect 34974 2592 34980 2604
rect 35032 2592 35038 2644
rect 36354 2592 36360 2644
rect 36412 2632 36418 2644
rect 36449 2635 36507 2641
rect 36449 2632 36461 2635
rect 36412 2604 36461 2632
rect 36412 2592 36418 2604
rect 36449 2601 36461 2604
rect 36495 2601 36507 2635
rect 36449 2595 36507 2601
rect 37734 2592 37740 2644
rect 37792 2632 37798 2644
rect 37829 2635 37887 2641
rect 37829 2632 37841 2635
rect 37792 2604 37841 2632
rect 37792 2592 37798 2604
rect 37829 2601 37841 2604
rect 37875 2601 37887 2635
rect 39850 2632 39856 2644
rect 39811 2604 39856 2632
rect 37829 2595 37887 2601
rect 39850 2592 39856 2604
rect 39908 2592 39914 2644
rect 40681 2635 40739 2641
rect 40681 2601 40693 2635
rect 40727 2632 40739 2635
rect 41598 2632 41604 2644
rect 40727 2604 41604 2632
rect 40727 2601 40739 2604
rect 40681 2595 40739 2601
rect 41598 2592 41604 2604
rect 41656 2592 41662 2644
rect 42334 2592 42340 2644
rect 42392 2632 42398 2644
rect 42429 2635 42487 2641
rect 42429 2632 42441 2635
rect 42392 2604 42441 2632
rect 42392 2592 42398 2604
rect 42429 2601 42441 2604
rect 42475 2601 42487 2635
rect 43530 2632 43536 2644
rect 43491 2604 43536 2632
rect 42429 2595 42487 2601
rect 43530 2592 43536 2604
rect 43588 2592 43594 2644
rect 45002 2632 45008 2644
rect 44963 2604 45008 2632
rect 45002 2592 45008 2604
rect 45060 2592 45066 2644
rect 46290 2592 46296 2644
rect 46348 2632 46354 2644
rect 46385 2635 46443 2641
rect 46385 2632 46397 2635
rect 46348 2604 46397 2632
rect 46348 2592 46354 2604
rect 46385 2601 46397 2604
rect 46431 2601 46443 2635
rect 57057 2635 57115 2641
rect 57057 2632 57069 2635
rect 46385 2595 46443 2601
rect 55186 2604 57069 2632
rect 55186 2564 55214 2604
rect 57057 2601 57069 2604
rect 57103 2601 57115 2635
rect 57057 2595 57115 2601
rect 16546 2536 55214 2564
rect 13280 2468 45554 2496
rect 13170 2428 13176 2440
rect 12299 2400 13032 2428
rect 13131 2400 13176 2428
rect 12299 2397 12311 2400
rect 12253 2391 12311 2397
rect 13170 2388 13176 2400
rect 13228 2388 13234 2440
rect 9784 2360 9812 2388
rect 13280 2360 13308 2468
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15197 2431 15255 2437
rect 15197 2428 15209 2431
rect 14976 2400 15209 2428
rect 14976 2388 14982 2400
rect 15197 2397 15209 2400
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 16298 2388 16304 2440
rect 16356 2428 16362 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16356 2400 16865 2428
rect 16356 2388 16362 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17770 2388 17776 2440
rect 17828 2428 17834 2440
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 17828 2400 18061 2428
rect 17828 2388 17834 2400
rect 18049 2397 18061 2400
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 19150 2388 19156 2440
rect 19208 2428 19214 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19208 2400 19441 2428
rect 19208 2388 19214 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 20622 2388 20628 2440
rect 20680 2428 20686 2440
rect 20901 2431 20959 2437
rect 20901 2428 20913 2431
rect 20680 2400 20913 2428
rect 20680 2388 20686 2400
rect 20901 2397 20913 2400
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22281 2431 22339 2437
rect 22281 2428 22293 2431
rect 22060 2400 22293 2428
rect 22060 2388 22066 2400
rect 22281 2397 22293 2400
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 23753 2431 23811 2437
rect 23753 2428 23765 2431
rect 23532 2400 23765 2428
rect 23532 2388 23538 2400
rect 23753 2397 23765 2400
rect 23799 2397 23811 2431
rect 23753 2391 23811 2397
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25133 2431 25191 2437
rect 25133 2428 25145 2431
rect 24912 2400 25145 2428
rect 24912 2388 24918 2400
rect 25133 2397 25145 2400
rect 25179 2397 25191 2431
rect 25133 2391 25191 2397
rect 26326 2388 26332 2440
rect 26384 2428 26390 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26384 2400 27169 2428
rect 26384 2388 26390 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 27985 2431 28043 2437
rect 27985 2428 27997 2431
rect 27764 2400 27997 2428
rect 27764 2388 27770 2400
rect 27985 2397 27997 2400
rect 28031 2397 28043 2431
rect 27985 2391 28043 2397
rect 29178 2388 29184 2440
rect 29236 2428 29242 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29236 2400 29745 2428
rect 29236 2388 29242 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 29733 2391 29791 2397
rect 30650 2388 30656 2440
rect 30708 2428 30714 2440
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 30708 2400 30941 2428
rect 30708 2388 30714 2400
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 32030 2388 32036 2440
rect 32088 2428 32094 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32088 2400 32321 2428
rect 32088 2388 32094 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 33781 2431 33839 2437
rect 33781 2428 33793 2431
rect 33560 2400 33793 2428
rect 33560 2388 33566 2400
rect 33781 2397 33793 2400
rect 33827 2397 33839 2431
rect 33781 2391 33839 2397
rect 34882 2388 34888 2440
rect 34940 2428 34946 2440
rect 35161 2431 35219 2437
rect 35161 2428 35173 2431
rect 34940 2400 35173 2428
rect 34940 2388 34946 2400
rect 35161 2397 35173 2400
rect 35207 2397 35219 2431
rect 35161 2391 35219 2397
rect 36354 2388 36360 2440
rect 36412 2428 36418 2440
rect 36633 2431 36691 2437
rect 36633 2428 36645 2431
rect 36412 2400 36645 2428
rect 36412 2388 36418 2400
rect 36633 2397 36645 2400
rect 36679 2397 36691 2431
rect 36633 2391 36691 2397
rect 37734 2388 37740 2440
rect 37792 2428 37798 2440
rect 38013 2431 38071 2437
rect 38013 2428 38025 2431
rect 37792 2400 38025 2428
rect 37792 2388 37798 2400
rect 38013 2397 38025 2400
rect 38059 2397 38071 2431
rect 38013 2391 38071 2397
rect 39206 2388 39212 2440
rect 39264 2428 39270 2440
rect 40037 2431 40095 2437
rect 40037 2428 40049 2431
rect 39264 2400 40049 2428
rect 39264 2388 39270 2400
rect 40037 2397 40049 2400
rect 40083 2397 40095 2431
rect 40037 2391 40095 2397
rect 40586 2388 40592 2440
rect 40644 2428 40650 2440
rect 40865 2431 40923 2437
rect 40865 2428 40877 2431
rect 40644 2400 40877 2428
rect 40644 2388 40650 2400
rect 40865 2397 40877 2400
rect 40911 2397 40923 2431
rect 40865 2391 40923 2397
rect 42058 2388 42064 2440
rect 42116 2428 42122 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 42116 2400 42625 2428
rect 42116 2388 42122 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 43438 2388 43444 2440
rect 43496 2428 43502 2440
rect 43717 2431 43775 2437
rect 43717 2428 43729 2431
rect 43496 2400 43729 2428
rect 43496 2388 43502 2400
rect 43717 2397 43729 2400
rect 43763 2397 43775 2431
rect 43717 2391 43775 2397
rect 44910 2388 44916 2440
rect 44968 2428 44974 2440
rect 45189 2431 45247 2437
rect 45189 2428 45201 2431
rect 44968 2400 45201 2428
rect 44968 2388 44974 2400
rect 45189 2397 45201 2400
rect 45235 2397 45247 2431
rect 45189 2391 45247 2397
rect 7208 2332 8984 2360
rect 9784 2332 13308 2360
rect 658 2252 664 2304
rect 716 2292 722 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 716 2264 1593 2292
rect 716 2252 722 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 2317 2295 2375 2301
rect 2317 2292 2329 2295
rect 2096 2264 2329 2292
rect 2096 2252 2102 2264
rect 2317 2261 2329 2264
rect 2363 2261 2375 2295
rect 2317 2255 2375 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5721 2295 5779 2301
rect 5721 2292 5733 2295
rect 5224 2264 5733 2292
rect 5224 2252 5230 2264
rect 5721 2261 5733 2264
rect 5767 2261 5779 2295
rect 5721 2255 5779 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8956 2301 8984 2332
rect 8113 2295 8171 2301
rect 8113 2292 8125 2295
rect 7800 2264 8125 2292
rect 7800 2252 7806 2264
rect 8113 2261 8125 2264
rect 8159 2261 8171 2295
rect 8113 2255 8171 2261
rect 8941 2295 8999 2301
rect 8941 2261 8953 2295
rect 8987 2261 8999 2295
rect 8941 2255 8999 2261
rect 10686 2252 10692 2304
rect 10744 2292 10750 2304
rect 11701 2295 11759 2301
rect 11701 2292 11713 2295
rect 10744 2264 11713 2292
rect 10744 2252 10750 2264
rect 11701 2261 11713 2264
rect 11747 2261 11759 2295
rect 11701 2255 11759 2261
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12124 2264 12449 2292
rect 12124 2252 12130 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 13446 2252 13452 2304
rect 13504 2292 13510 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13504 2264 14289 2292
rect 13504 2252 13510 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 45526 2292 45554 2468
rect 48038 2456 48044 2508
rect 48096 2496 48102 2508
rect 48133 2499 48191 2505
rect 48133 2496 48145 2499
rect 48096 2468 48145 2496
rect 48096 2456 48102 2468
rect 48133 2465 48145 2468
rect 48179 2465 48191 2499
rect 50982 2496 50988 2508
rect 50943 2468 50988 2496
rect 48133 2459 48191 2465
rect 50982 2456 50988 2468
rect 51040 2456 51046 2508
rect 52362 2456 52368 2508
rect 52420 2496 52426 2508
rect 53009 2499 53067 2505
rect 53009 2496 53021 2499
rect 52420 2468 53021 2496
rect 52420 2456 52426 2468
rect 53009 2465 53021 2468
rect 53055 2465 53067 2499
rect 53009 2459 53067 2465
rect 55490 2456 55496 2508
rect 55548 2496 55554 2508
rect 55585 2499 55643 2505
rect 55585 2496 55597 2499
rect 55548 2468 55597 2496
rect 55548 2456 55554 2468
rect 55585 2465 55597 2468
rect 55631 2465 55643 2499
rect 55585 2459 55643 2465
rect 46290 2388 46296 2440
rect 46348 2428 46354 2440
rect 46569 2431 46627 2437
rect 46569 2428 46581 2431
rect 46348 2400 46581 2428
rect 46348 2388 46354 2400
rect 46569 2397 46581 2400
rect 46615 2397 46627 2431
rect 46569 2391 46627 2397
rect 47762 2388 47768 2440
rect 47820 2428 47826 2440
rect 47857 2431 47915 2437
rect 47857 2428 47869 2431
rect 47820 2400 47869 2428
rect 47820 2388 47826 2400
rect 47857 2397 47869 2400
rect 47903 2397 47915 2431
rect 47857 2391 47915 2397
rect 50614 2388 50620 2440
rect 50672 2428 50678 2440
rect 50709 2431 50767 2437
rect 50709 2428 50721 2431
rect 50672 2400 50721 2428
rect 50672 2388 50678 2400
rect 50709 2397 50721 2400
rect 50755 2397 50767 2431
rect 50709 2391 50767 2397
rect 51994 2388 52000 2440
rect 52052 2428 52058 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52052 2400 52745 2428
rect 52052 2388 52058 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 54846 2388 54852 2440
rect 54904 2428 54910 2440
rect 55309 2431 55367 2437
rect 55309 2428 55321 2431
rect 54904 2400 55321 2428
rect 54904 2388 54910 2400
rect 55309 2397 55321 2400
rect 55355 2397 55367 2431
rect 55309 2391 55367 2397
rect 54389 2363 54447 2369
rect 54389 2329 54401 2363
rect 54435 2360 54447 2363
rect 55122 2360 55128 2372
rect 54435 2332 55128 2360
rect 54435 2329 54447 2332
rect 54389 2323 54447 2329
rect 55122 2320 55128 2332
rect 55180 2320 55186 2372
rect 56962 2360 56968 2372
rect 56923 2332 56968 2360
rect 56962 2320 56968 2332
rect 57020 2320 57026 2372
rect 54481 2295 54539 2301
rect 54481 2292 54493 2295
rect 45526 2264 54493 2292
rect 14277 2255 14335 2261
rect 54481 2261 54493 2264
rect 54527 2261 54539 2295
rect 54481 2255 54539 2261
rect 1104 2202 58880 2224
rect 1104 2150 20214 2202
rect 20266 2150 20278 2202
rect 20330 2150 20342 2202
rect 20394 2150 20406 2202
rect 20458 2150 20470 2202
rect 20522 2150 39478 2202
rect 39530 2150 39542 2202
rect 39594 2150 39606 2202
rect 39658 2150 39670 2202
rect 39722 2150 39734 2202
rect 39786 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 53012 19796 53064 19848
rect 57152 19796 57204 19848
rect 53380 19728 53432 19780
rect 56968 19728 57020 19780
rect 53932 19660 53984 19712
rect 57060 19660 57112 19712
rect 20214 19558 20266 19610
rect 20278 19558 20330 19610
rect 20342 19558 20394 19610
rect 20406 19558 20458 19610
rect 20470 19558 20522 19610
rect 39478 19558 39530 19610
rect 39542 19558 39594 19610
rect 39606 19558 39658 19610
rect 39670 19558 39722 19610
rect 39734 19558 39786 19610
rect 1032 19456 1084 19508
rect 2320 19499 2372 19508
rect 2320 19465 2329 19499
rect 2329 19465 2363 19499
rect 2363 19465 2372 19499
rect 2320 19456 2372 19465
rect 3516 19456 3568 19508
rect 5172 19499 5224 19508
rect 5172 19465 5181 19499
rect 5181 19465 5215 19499
rect 5215 19465 5224 19499
rect 5172 19456 5224 19465
rect 6644 19499 6696 19508
rect 6644 19465 6653 19499
rect 6653 19465 6687 19499
rect 6687 19465 6696 19499
rect 6644 19456 6696 19465
rect 8024 19499 8076 19508
rect 8024 19465 8033 19499
rect 8033 19465 8067 19499
rect 8067 19465 8076 19499
rect 8024 19456 8076 19465
rect 9496 19499 9548 19508
rect 9496 19465 9505 19499
rect 9505 19465 9539 19499
rect 9539 19465 9548 19499
rect 9496 19456 9548 19465
rect 10876 19499 10928 19508
rect 10876 19465 10885 19499
rect 10885 19465 10919 19499
rect 10919 19465 10928 19499
rect 10876 19456 10928 19465
rect 12348 19499 12400 19508
rect 12348 19465 12357 19499
rect 12357 19465 12391 19499
rect 12391 19465 12400 19499
rect 12348 19456 12400 19465
rect 13452 19456 13504 19508
rect 16396 19456 16448 19508
rect 20076 19456 20128 19508
rect 22560 19456 22612 19508
rect 27344 19456 27396 19508
rect 29644 19456 29696 19508
rect 31024 19456 31076 19508
rect 32496 19456 32548 19508
rect 33692 19456 33744 19508
rect 35072 19456 35124 19508
rect 39304 19456 39356 19508
rect 41512 19456 41564 19508
rect 41880 19456 41932 19508
rect 43996 19456 44048 19508
rect 45376 19456 45428 19508
rect 48964 19456 49016 19508
rect 51172 19456 51224 19508
rect 56232 19456 56284 19508
rect 56508 19499 56560 19508
rect 56508 19465 56517 19499
rect 56517 19465 56551 19499
rect 56551 19465 56560 19499
rect 56508 19456 56560 19465
rect 57888 19456 57940 19508
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2136 19363 2188 19372
rect 2136 19329 2145 19363
rect 2145 19329 2179 19363
rect 2179 19329 2188 19363
rect 2136 19320 2188 19329
rect 3792 19363 3844 19372
rect 3792 19329 3801 19363
rect 3801 19329 3835 19363
rect 3835 19329 3844 19363
rect 3792 19320 3844 19329
rect 5080 19320 5132 19372
rect 6552 19320 6604 19372
rect 7932 19320 7984 19372
rect 9404 19320 9456 19372
rect 10508 19320 10560 19372
rect 12072 19320 12124 19372
rect 14096 19363 14148 19372
rect 14096 19329 14105 19363
rect 14105 19329 14139 19363
rect 14139 19329 14148 19363
rect 14096 19320 14148 19329
rect 14924 19320 14976 19372
rect 16304 19320 16356 19372
rect 17776 19320 17828 19372
rect 19156 19320 19208 19372
rect 20628 19320 20680 19372
rect 22008 19320 22060 19372
rect 23756 19363 23808 19372
rect 23756 19329 23765 19363
rect 23765 19329 23799 19363
rect 23799 19329 23808 19363
rect 23756 19320 23808 19329
rect 25136 19363 25188 19372
rect 25136 19329 25145 19363
rect 25145 19329 25179 19363
rect 25179 19329 25188 19363
rect 25136 19320 25188 19329
rect 26332 19320 26384 19372
rect 27988 19363 28040 19372
rect 27988 19329 27997 19363
rect 27997 19329 28031 19363
rect 28031 19329 28040 19363
rect 27988 19320 28040 19329
rect 29184 19320 29236 19372
rect 30932 19363 30984 19372
rect 30932 19329 30941 19363
rect 30941 19329 30975 19363
rect 30975 19329 30984 19363
rect 30932 19320 30984 19329
rect 32312 19363 32364 19372
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 33784 19363 33836 19372
rect 33784 19329 33793 19363
rect 33793 19329 33827 19363
rect 33827 19329 33836 19363
rect 33784 19320 33836 19329
rect 35164 19363 35216 19372
rect 35164 19329 35173 19363
rect 35173 19329 35207 19363
rect 35207 19329 35216 19363
rect 35164 19320 35216 19329
rect 36636 19363 36688 19372
rect 36636 19329 36645 19363
rect 36645 19329 36679 19363
rect 36679 19329 36688 19363
rect 36636 19320 36688 19329
rect 38016 19363 38068 19372
rect 38016 19329 38025 19363
rect 38025 19329 38059 19363
rect 38059 19329 38068 19363
rect 38016 19320 38068 19329
rect 39212 19320 39264 19372
rect 40868 19363 40920 19372
rect 40868 19329 40877 19363
rect 40877 19329 40911 19363
rect 40911 19329 40920 19363
rect 40868 19320 40920 19329
rect 42064 19320 42116 19372
rect 43720 19363 43772 19372
rect 43720 19329 43729 19363
rect 43729 19329 43763 19363
rect 43763 19329 43772 19363
rect 43720 19320 43772 19329
rect 44916 19320 44968 19372
rect 46572 19363 46624 19372
rect 46572 19329 46581 19363
rect 46581 19329 46615 19363
rect 46615 19329 46624 19363
rect 46572 19320 46624 19329
rect 48044 19363 48096 19372
rect 48044 19329 48053 19363
rect 48053 19329 48087 19363
rect 48087 19329 48096 19363
rect 48044 19320 48096 19329
rect 49424 19363 49476 19372
rect 49424 19329 49433 19363
rect 49433 19329 49467 19363
rect 49467 19329 49476 19363
rect 49424 19320 49476 19329
rect 50896 19363 50948 19372
rect 50896 19329 50905 19363
rect 50905 19329 50939 19363
rect 50939 19329 50948 19363
rect 50896 19320 50948 19329
rect 52184 19363 52236 19372
rect 52184 19329 52193 19363
rect 52193 19329 52227 19363
rect 52227 19329 52236 19363
rect 52184 19320 52236 19329
rect 53380 19363 53432 19372
rect 53380 19329 53389 19363
rect 53389 19329 53423 19363
rect 53423 19329 53432 19363
rect 53380 19320 53432 19329
rect 54024 19363 54076 19372
rect 54024 19329 54033 19363
rect 54033 19329 54067 19363
rect 54067 19329 54076 19363
rect 54024 19320 54076 19329
rect 55588 19363 55640 19372
rect 55588 19329 55597 19363
rect 55597 19329 55631 19363
rect 55631 19329 55640 19363
rect 55588 19320 55640 19329
rect 55772 19320 55824 19372
rect 57060 19363 57112 19372
rect 57060 19329 57069 19363
rect 57069 19329 57103 19363
rect 57103 19329 57112 19363
rect 57060 19320 57112 19329
rect 57152 19320 57204 19372
rect 15016 19159 15068 19168
rect 15016 19125 15025 19159
rect 15025 19125 15059 19159
rect 15059 19125 15068 19159
rect 15016 19116 15068 19125
rect 17868 19159 17920 19168
rect 17868 19125 17877 19159
rect 17877 19125 17911 19159
rect 17911 19125 17920 19159
rect 17868 19116 17920 19125
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 23572 19159 23624 19168
rect 23572 19125 23581 19159
rect 23581 19125 23615 19159
rect 23615 19125 23624 19159
rect 23572 19116 23624 19125
rect 24952 19159 25004 19168
rect 24952 19125 24961 19159
rect 24961 19125 24995 19159
rect 24995 19125 25004 19159
rect 24952 19116 25004 19125
rect 27804 19159 27856 19168
rect 27804 19125 27813 19159
rect 27813 19125 27847 19159
rect 27847 19125 27856 19159
rect 27804 19116 27856 19125
rect 36452 19159 36504 19168
rect 36452 19125 36461 19159
rect 36461 19125 36495 19159
rect 36495 19125 36504 19159
rect 36452 19116 36504 19125
rect 37832 19159 37884 19168
rect 37832 19125 37841 19159
rect 37841 19125 37875 19159
rect 37875 19125 37884 19159
rect 37832 19116 37884 19125
rect 46388 19159 46440 19168
rect 46388 19125 46397 19159
rect 46397 19125 46431 19159
rect 46431 19125 46440 19159
rect 46388 19116 46440 19125
rect 47860 19159 47912 19168
rect 47860 19125 47869 19159
rect 47869 19125 47903 19159
rect 47903 19125 47912 19159
rect 47860 19116 47912 19125
rect 52276 19116 52328 19168
rect 57244 19159 57296 19168
rect 57244 19125 57253 19159
rect 57253 19125 57287 19159
rect 57287 19125 57296 19159
rect 57244 19116 57296 19125
rect 10582 19014 10634 19066
rect 10646 19014 10698 19066
rect 10710 19014 10762 19066
rect 10774 19014 10826 19066
rect 10838 19014 10890 19066
rect 29846 19014 29898 19066
rect 29910 19014 29962 19066
rect 29974 19014 30026 19066
rect 30038 19014 30090 19066
rect 30102 19014 30154 19066
rect 49110 19014 49162 19066
rect 49174 19014 49226 19066
rect 49238 19014 49290 19066
rect 49302 19014 49354 19066
rect 49366 19014 49418 19066
rect 54024 18912 54076 18964
rect 55588 18912 55640 18964
rect 51080 18844 51132 18896
rect 55864 18776 55916 18828
rect 51172 18751 51224 18760
rect 51172 18717 51181 18751
rect 51181 18717 51215 18751
rect 51215 18717 51224 18751
rect 51172 18708 51224 18717
rect 52368 18708 52420 18760
rect 50804 18615 50856 18624
rect 50804 18581 50813 18615
rect 50813 18581 50847 18615
rect 50847 18581 50856 18615
rect 50804 18572 50856 18581
rect 50988 18572 51040 18624
rect 52000 18615 52052 18624
rect 52000 18581 52009 18615
rect 52009 18581 52043 18615
rect 52043 18581 52052 18615
rect 52000 18572 52052 18581
rect 52276 18572 52328 18624
rect 53564 18615 53616 18624
rect 53564 18581 53573 18615
rect 53573 18581 53607 18615
rect 53607 18581 53616 18615
rect 53564 18572 53616 18581
rect 53840 18572 53892 18624
rect 55496 18640 55548 18692
rect 56692 18640 56744 18692
rect 55680 18615 55732 18624
rect 55680 18581 55689 18615
rect 55689 18581 55723 18615
rect 55723 18581 55732 18615
rect 55680 18572 55732 18581
rect 56508 18615 56560 18624
rect 56508 18581 56517 18615
rect 56517 18581 56551 18615
rect 56551 18581 56560 18615
rect 56508 18572 56560 18581
rect 56876 18615 56928 18624
rect 56876 18581 56885 18615
rect 56885 18581 56919 18615
rect 56919 18581 56928 18615
rect 56876 18572 56928 18581
rect 58072 18615 58124 18624
rect 58072 18581 58081 18615
rect 58081 18581 58115 18615
rect 58115 18581 58124 18615
rect 58072 18572 58124 18581
rect 20214 18470 20266 18522
rect 20278 18470 20330 18522
rect 20342 18470 20394 18522
rect 20406 18470 20458 18522
rect 20470 18470 20522 18522
rect 39478 18470 39530 18522
rect 39542 18470 39594 18522
rect 39606 18470 39658 18522
rect 39670 18470 39722 18522
rect 39734 18470 39786 18522
rect 53012 18368 53064 18420
rect 53564 18411 53616 18420
rect 53564 18377 53573 18411
rect 53573 18377 53607 18411
rect 53607 18377 53616 18411
rect 53564 18368 53616 18377
rect 55680 18368 55732 18420
rect 56048 18411 56100 18420
rect 56048 18377 56057 18411
rect 56057 18377 56091 18411
rect 56091 18377 56100 18411
rect 56048 18368 56100 18377
rect 50804 18232 50856 18284
rect 52000 18232 52052 18284
rect 53748 18275 53800 18284
rect 53748 18241 53757 18275
rect 53757 18241 53791 18275
rect 53791 18241 53800 18275
rect 53748 18232 53800 18241
rect 54760 18275 54812 18284
rect 54760 18241 54769 18275
rect 54769 18241 54803 18275
rect 54803 18241 54812 18275
rect 54760 18232 54812 18241
rect 56508 18300 56560 18352
rect 57704 18300 57756 18352
rect 56600 18232 56652 18284
rect 57244 18232 57296 18284
rect 53932 18096 53984 18148
rect 56784 18164 56836 18216
rect 57428 18028 57480 18080
rect 57888 18028 57940 18080
rect 10582 17926 10634 17978
rect 10646 17926 10698 17978
rect 10710 17926 10762 17978
rect 10774 17926 10826 17978
rect 10838 17926 10890 17978
rect 29846 17926 29898 17978
rect 29910 17926 29962 17978
rect 29974 17926 30026 17978
rect 30038 17926 30090 17978
rect 30102 17926 30154 17978
rect 49110 17926 49162 17978
rect 49174 17926 49226 17978
rect 49238 17926 49290 17978
rect 49302 17926 49354 17978
rect 49366 17926 49418 17978
rect 55864 17867 55916 17876
rect 48228 17688 48280 17740
rect 46020 17620 46072 17672
rect 47584 17620 47636 17672
rect 48964 17663 49016 17672
rect 48964 17629 48973 17663
rect 48973 17629 49007 17663
rect 49007 17629 49016 17663
rect 48964 17620 49016 17629
rect 55864 17833 55873 17867
rect 55873 17833 55907 17867
rect 55907 17833 55916 17867
rect 55864 17824 55916 17833
rect 55956 17824 56008 17876
rect 56968 17824 57020 17876
rect 56784 17756 56836 17808
rect 57244 17688 57296 17740
rect 57152 17620 57204 17672
rect 55772 17595 55824 17604
rect 55772 17561 55781 17595
rect 55781 17561 55815 17595
rect 55815 17561 55824 17595
rect 55772 17552 55824 17561
rect 56968 17552 57020 17604
rect 46756 17527 46808 17536
rect 46756 17493 46765 17527
rect 46765 17493 46799 17527
rect 46799 17493 46808 17527
rect 46756 17484 46808 17493
rect 49516 17484 49568 17536
rect 51080 17484 51132 17536
rect 57520 17527 57572 17536
rect 57520 17493 57529 17527
rect 57529 17493 57563 17527
rect 57563 17493 57572 17527
rect 57520 17484 57572 17493
rect 20214 17382 20266 17434
rect 20278 17382 20330 17434
rect 20342 17382 20394 17434
rect 20406 17382 20458 17434
rect 20470 17382 20522 17434
rect 39478 17382 39530 17434
rect 39542 17382 39594 17434
rect 39606 17382 39658 17434
rect 39670 17382 39722 17434
rect 39734 17382 39786 17434
rect 46020 17323 46072 17332
rect 46020 17289 46029 17323
rect 46029 17289 46063 17323
rect 46063 17289 46072 17323
rect 46020 17280 46072 17289
rect 46388 17323 46440 17332
rect 46388 17289 46397 17323
rect 46397 17289 46431 17323
rect 46431 17289 46440 17323
rect 46388 17280 46440 17289
rect 47584 17323 47636 17332
rect 47584 17289 47593 17323
rect 47593 17289 47627 17323
rect 47627 17289 47636 17323
rect 47584 17280 47636 17289
rect 47860 17280 47912 17332
rect 46756 17212 46808 17264
rect 42984 17144 43036 17196
rect 46296 17076 46348 17128
rect 45008 16983 45060 16992
rect 45008 16949 45017 16983
rect 45017 16949 45051 16983
rect 45051 16949 45060 16983
rect 56324 17144 56376 17196
rect 57612 17144 57664 17196
rect 48044 17119 48096 17128
rect 48044 17085 48053 17119
rect 48053 17085 48087 17119
rect 48087 17085 48096 17119
rect 48044 17076 48096 17085
rect 48228 17119 48280 17128
rect 48228 17085 48237 17119
rect 48237 17085 48271 17119
rect 48271 17085 48280 17119
rect 48228 17076 48280 17085
rect 55772 17008 55824 17060
rect 56876 17008 56928 17060
rect 57244 17051 57296 17060
rect 57244 17017 57253 17051
rect 57253 17017 57287 17051
rect 57287 17017 57296 17051
rect 57244 17008 57296 17017
rect 45008 16940 45060 16949
rect 48228 16940 48280 16992
rect 58072 16983 58124 16992
rect 58072 16949 58081 16983
rect 58081 16949 58115 16983
rect 58115 16949 58124 16983
rect 58072 16940 58124 16949
rect 10582 16838 10634 16890
rect 10646 16838 10698 16890
rect 10710 16838 10762 16890
rect 10774 16838 10826 16890
rect 10838 16838 10890 16890
rect 29846 16838 29898 16890
rect 29910 16838 29962 16890
rect 29974 16838 30026 16890
rect 30038 16838 30090 16890
rect 30102 16838 30154 16890
rect 49110 16838 49162 16890
rect 49174 16838 49226 16890
rect 49238 16838 49290 16890
rect 49302 16838 49354 16890
rect 49366 16838 49418 16890
rect 45008 16736 45060 16788
rect 57152 16736 57204 16788
rect 43536 16600 43588 16652
rect 45008 16600 45060 16652
rect 57060 16668 57112 16720
rect 59176 16668 59228 16720
rect 43996 16575 44048 16584
rect 43996 16541 44005 16575
rect 44005 16541 44039 16575
rect 44039 16541 44048 16575
rect 43996 16532 44048 16541
rect 45376 16575 45428 16584
rect 45376 16541 45385 16575
rect 45385 16541 45419 16575
rect 45419 16541 45428 16575
rect 45376 16532 45428 16541
rect 57060 16532 57112 16584
rect 57428 16575 57480 16584
rect 57428 16541 57437 16575
rect 57437 16541 57471 16575
rect 57471 16541 57480 16575
rect 57428 16532 57480 16541
rect 57888 16575 57940 16584
rect 57888 16541 57897 16575
rect 57897 16541 57931 16575
rect 57931 16541 57940 16575
rect 57888 16532 57940 16541
rect 43628 16439 43680 16448
rect 43628 16405 43637 16439
rect 43637 16405 43671 16439
rect 43671 16405 43680 16439
rect 43628 16396 43680 16405
rect 57612 16464 57664 16516
rect 56600 16439 56652 16448
rect 56600 16405 56609 16439
rect 56609 16405 56643 16439
rect 56643 16405 56652 16439
rect 56600 16396 56652 16405
rect 58072 16439 58124 16448
rect 58072 16405 58081 16439
rect 58081 16405 58115 16439
rect 58115 16405 58124 16439
rect 58072 16396 58124 16405
rect 20214 16294 20266 16346
rect 20278 16294 20330 16346
rect 20342 16294 20394 16346
rect 20406 16294 20458 16346
rect 20470 16294 20522 16346
rect 39478 16294 39530 16346
rect 39542 16294 39594 16346
rect 39606 16294 39658 16346
rect 39670 16294 39722 16346
rect 39734 16294 39786 16346
rect 57520 16192 57572 16244
rect 43628 16056 43680 16108
rect 57336 16099 57388 16108
rect 57336 16065 57345 16099
rect 57345 16065 57379 16099
rect 57379 16065 57388 16099
rect 57336 16056 57388 16065
rect 57428 16056 57480 16108
rect 57888 15852 57940 15904
rect 58072 15895 58124 15904
rect 58072 15861 58081 15895
rect 58081 15861 58115 15895
rect 58115 15861 58124 15895
rect 58072 15852 58124 15861
rect 10582 15750 10634 15802
rect 10646 15750 10698 15802
rect 10710 15750 10762 15802
rect 10774 15750 10826 15802
rect 10838 15750 10890 15802
rect 29846 15750 29898 15802
rect 29910 15750 29962 15802
rect 29974 15750 30026 15802
rect 30038 15750 30090 15802
rect 30102 15750 30154 15802
rect 49110 15750 49162 15802
rect 49174 15750 49226 15802
rect 49238 15750 49290 15802
rect 49302 15750 49354 15802
rect 49366 15750 49418 15802
rect 42064 15555 42116 15564
rect 42064 15521 42073 15555
rect 42073 15521 42107 15555
rect 42107 15521 42116 15555
rect 42064 15512 42116 15521
rect 41880 15487 41932 15496
rect 41880 15453 41889 15487
rect 41889 15453 41923 15487
rect 41923 15453 41932 15487
rect 41880 15444 41932 15453
rect 56600 15444 56652 15496
rect 41880 15308 41932 15360
rect 42340 15308 42392 15360
rect 57888 15308 57940 15360
rect 20214 15206 20266 15258
rect 20278 15206 20330 15258
rect 20342 15206 20394 15258
rect 20406 15206 20458 15258
rect 20470 15206 20522 15258
rect 39478 15206 39530 15258
rect 39542 15206 39594 15258
rect 39606 15206 39658 15258
rect 39670 15206 39722 15258
rect 39734 15206 39786 15258
rect 39304 15147 39356 15156
rect 39304 15113 39313 15147
rect 39313 15113 39347 15147
rect 39347 15113 39356 15147
rect 39304 15104 39356 15113
rect 39764 14968 39816 15020
rect 38108 14832 38160 14884
rect 41144 14900 41196 14952
rect 41880 14900 41932 14952
rect 57428 15036 57480 15088
rect 50252 14968 50304 15020
rect 56600 14900 56652 14952
rect 42064 14832 42116 14884
rect 39856 14764 39908 14816
rect 58072 14807 58124 14816
rect 58072 14773 58081 14807
rect 58081 14773 58115 14807
rect 58115 14773 58124 14807
rect 58072 14764 58124 14773
rect 10582 14662 10634 14714
rect 10646 14662 10698 14714
rect 10710 14662 10762 14714
rect 10774 14662 10826 14714
rect 10838 14662 10890 14714
rect 29846 14662 29898 14714
rect 29910 14662 29962 14714
rect 29974 14662 30026 14714
rect 30038 14662 30090 14714
rect 30102 14662 30154 14714
rect 49110 14662 49162 14714
rect 49174 14662 49226 14714
rect 49238 14662 49290 14714
rect 49302 14662 49354 14714
rect 49366 14662 49418 14714
rect 41144 14603 41196 14612
rect 41144 14569 41153 14603
rect 41153 14569 41187 14603
rect 41187 14569 41196 14603
rect 41144 14560 41196 14569
rect 38108 14467 38160 14476
rect 38108 14433 38117 14467
rect 38117 14433 38151 14467
rect 38151 14433 38160 14467
rect 38108 14424 38160 14433
rect 39856 14467 39908 14476
rect 39856 14433 39865 14467
rect 39865 14433 39899 14467
rect 39899 14433 39908 14467
rect 39856 14424 39908 14433
rect 42064 14424 42116 14476
rect 37832 14399 37884 14408
rect 37832 14365 37841 14399
rect 37841 14365 37875 14399
rect 37875 14365 37884 14399
rect 37832 14356 37884 14365
rect 50252 14356 50304 14408
rect 50344 14356 50396 14408
rect 41512 14331 41564 14340
rect 41512 14297 41521 14331
rect 41521 14297 41555 14331
rect 41555 14297 41564 14331
rect 41512 14288 41564 14297
rect 37464 14263 37516 14272
rect 37464 14229 37473 14263
rect 37473 14229 37507 14263
rect 37507 14229 37516 14263
rect 37464 14220 37516 14229
rect 37740 14220 37792 14272
rect 41604 14263 41656 14272
rect 41604 14229 41613 14263
rect 41613 14229 41647 14263
rect 41647 14229 41656 14263
rect 58072 14263 58124 14272
rect 41604 14220 41656 14229
rect 58072 14229 58081 14263
rect 58081 14229 58115 14263
rect 58115 14229 58124 14263
rect 58072 14220 58124 14229
rect 20214 14118 20266 14170
rect 20278 14118 20330 14170
rect 20342 14118 20394 14170
rect 20406 14118 20458 14170
rect 20470 14118 20522 14170
rect 39478 14118 39530 14170
rect 39542 14118 39594 14170
rect 39606 14118 39658 14170
rect 39670 14118 39722 14170
rect 39734 14118 39786 14170
rect 57888 14016 57940 14068
rect 37464 13880 37516 13932
rect 52460 13880 52512 13932
rect 50344 13812 50396 13864
rect 10582 13574 10634 13626
rect 10646 13574 10698 13626
rect 10710 13574 10762 13626
rect 10774 13574 10826 13626
rect 10838 13574 10890 13626
rect 29846 13574 29898 13626
rect 29910 13574 29962 13626
rect 29974 13574 30026 13626
rect 30038 13574 30090 13626
rect 30102 13574 30154 13626
rect 49110 13574 49162 13626
rect 49174 13574 49226 13626
rect 49238 13574 49290 13626
rect 49302 13574 49354 13626
rect 49366 13574 49418 13626
rect 36452 13311 36504 13320
rect 36452 13277 36461 13311
rect 36461 13277 36495 13311
rect 36495 13277 36504 13311
rect 36452 13268 36504 13277
rect 52460 13268 52512 13320
rect 52552 13268 52604 13320
rect 38108 13200 38160 13252
rect 36360 13132 36412 13184
rect 58072 13175 58124 13184
rect 58072 13141 58081 13175
rect 58081 13141 58115 13175
rect 58115 13141 58124 13175
rect 58072 13132 58124 13141
rect 20214 13030 20266 13082
rect 20278 13030 20330 13082
rect 20342 13030 20394 13082
rect 20406 13030 20458 13082
rect 20470 13030 20522 13082
rect 39478 13030 39530 13082
rect 39542 13030 39594 13082
rect 39606 13030 39658 13082
rect 39670 13030 39722 13082
rect 39734 13030 39786 13082
rect 38108 12928 38160 12980
rect 35164 12835 35216 12844
rect 35164 12801 35173 12835
rect 35173 12801 35207 12835
rect 35207 12801 35216 12835
rect 35164 12792 35216 12801
rect 38384 12792 38436 12844
rect 34244 12724 34296 12776
rect 52552 12656 52604 12708
rect 58072 12631 58124 12640
rect 58072 12597 58081 12631
rect 58081 12597 58115 12631
rect 58115 12597 58124 12631
rect 58072 12588 58124 12597
rect 10582 12486 10634 12538
rect 10646 12486 10698 12538
rect 10710 12486 10762 12538
rect 10774 12486 10826 12538
rect 10838 12486 10890 12538
rect 29846 12486 29898 12538
rect 29910 12486 29962 12538
rect 29974 12486 30026 12538
rect 30038 12486 30090 12538
rect 30102 12486 30154 12538
rect 49110 12486 49162 12538
rect 49174 12486 49226 12538
rect 49238 12486 49290 12538
rect 49302 12486 49354 12538
rect 49366 12486 49418 12538
rect 35164 12384 35216 12436
rect 32772 12248 32824 12300
rect 50344 12248 50396 12300
rect 33692 12223 33744 12232
rect 33692 12189 33701 12223
rect 33701 12189 33735 12223
rect 33735 12189 33744 12223
rect 33692 12180 33744 12189
rect 35072 12223 35124 12232
rect 35072 12189 35081 12223
rect 35081 12189 35115 12223
rect 35115 12189 35124 12223
rect 35072 12180 35124 12189
rect 38660 12223 38712 12232
rect 38660 12189 38669 12223
rect 38669 12189 38703 12223
rect 38703 12189 38712 12223
rect 38660 12180 38712 12189
rect 30656 12112 30708 12164
rect 32128 12112 32180 12164
rect 33324 12087 33376 12096
rect 33324 12053 33333 12087
rect 33333 12053 33367 12087
rect 33367 12053 33376 12087
rect 33324 12044 33376 12053
rect 33600 12044 33652 12096
rect 34980 12044 35032 12096
rect 38384 12044 38436 12096
rect 58072 12087 58124 12096
rect 58072 12053 58081 12087
rect 58081 12053 58115 12087
rect 58115 12053 58124 12087
rect 58072 12044 58124 12053
rect 20214 11942 20266 11994
rect 20278 11942 20330 11994
rect 20342 11942 20394 11994
rect 20406 11942 20458 11994
rect 20470 11942 20522 11994
rect 39478 11942 39530 11994
rect 39542 11942 39594 11994
rect 39606 11942 39658 11994
rect 39670 11942 39722 11994
rect 39734 11942 39786 11994
rect 29644 11840 29696 11892
rect 30656 11883 30708 11892
rect 30656 11849 30665 11883
rect 30665 11849 30699 11883
rect 30699 11849 30708 11883
rect 30656 11840 30708 11849
rect 31024 11883 31076 11892
rect 31024 11849 31033 11883
rect 31033 11849 31067 11883
rect 31067 11849 31076 11883
rect 31024 11840 31076 11849
rect 32128 11883 32180 11892
rect 32128 11849 32137 11883
rect 32137 11849 32171 11883
rect 32171 11849 32180 11883
rect 32128 11840 32180 11849
rect 32496 11883 32548 11892
rect 32496 11849 32505 11883
rect 32505 11849 32539 11883
rect 32539 11849 32548 11883
rect 32496 11840 32548 11849
rect 33324 11772 33376 11824
rect 34244 11815 34296 11824
rect 34244 11781 34253 11815
rect 34253 11781 34287 11815
rect 34287 11781 34296 11815
rect 34244 11772 34296 11781
rect 29552 11636 29604 11688
rect 31024 11704 31076 11756
rect 30748 11636 30800 11688
rect 50344 11704 50396 11756
rect 32128 11636 32180 11688
rect 32772 11679 32824 11688
rect 32772 11645 32781 11679
rect 32781 11645 32815 11679
rect 32815 11645 32824 11679
rect 32772 11636 32824 11645
rect 30196 11500 30248 11552
rect 58072 11543 58124 11552
rect 58072 11509 58081 11543
rect 58081 11509 58115 11543
rect 58115 11509 58124 11543
rect 58072 11500 58124 11509
rect 10582 11398 10634 11450
rect 10646 11398 10698 11450
rect 10710 11398 10762 11450
rect 10774 11398 10826 11450
rect 10838 11398 10890 11450
rect 29846 11398 29898 11450
rect 29910 11398 29962 11450
rect 29974 11398 30026 11450
rect 30038 11398 30090 11450
rect 30102 11398 30154 11450
rect 49110 11398 49162 11450
rect 49174 11398 49226 11450
rect 49238 11398 49290 11450
rect 49302 11398 49354 11450
rect 49366 11398 49418 11450
rect 31024 11339 31076 11348
rect 31024 11305 31033 11339
rect 31033 11305 31067 11339
rect 31067 11305 31076 11339
rect 31024 11296 31076 11305
rect 38660 11228 38712 11280
rect 30196 11135 30248 11144
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 42984 11228 43036 11280
rect 57888 11228 57940 11280
rect 40224 11160 40276 11212
rect 56784 11160 56836 11212
rect 26516 11024 26568 11076
rect 38384 11024 38436 11076
rect 40224 11024 40276 11076
rect 20214 10854 20266 10906
rect 20278 10854 20330 10906
rect 20342 10854 20394 10906
rect 20406 10854 20458 10906
rect 20470 10854 20522 10906
rect 39478 10854 39530 10906
rect 39542 10854 39594 10906
rect 39606 10854 39658 10906
rect 39670 10854 39722 10906
rect 39734 10854 39786 10906
rect 57060 10659 57112 10668
rect 57060 10625 57069 10659
rect 57069 10625 57103 10659
rect 57103 10625 57112 10659
rect 57060 10616 57112 10625
rect 57152 10616 57204 10668
rect 57244 10455 57296 10464
rect 57244 10421 57253 10455
rect 57253 10421 57287 10455
rect 57287 10421 57296 10455
rect 57244 10412 57296 10421
rect 58072 10455 58124 10464
rect 58072 10421 58081 10455
rect 58081 10421 58115 10455
rect 58115 10421 58124 10455
rect 58072 10412 58124 10421
rect 10582 10310 10634 10362
rect 10646 10310 10698 10362
rect 10710 10310 10762 10362
rect 10774 10310 10826 10362
rect 10838 10310 10890 10362
rect 29846 10310 29898 10362
rect 29910 10310 29962 10362
rect 29974 10310 30026 10362
rect 30038 10310 30090 10362
rect 30102 10310 30154 10362
rect 49110 10310 49162 10362
rect 49174 10310 49226 10362
rect 49238 10310 49290 10362
rect 49302 10310 49354 10362
rect 49366 10310 49418 10362
rect 26884 9979 26936 9988
rect 26884 9945 26893 9979
rect 26893 9945 26927 9979
rect 26927 9945 26936 9979
rect 26884 9936 26936 9945
rect 27988 9979 28040 9988
rect 27988 9945 27997 9979
rect 27997 9945 28031 9979
rect 28031 9945 28040 9979
rect 27988 9936 28040 9945
rect 57060 10004 57112 10056
rect 57152 9936 57204 9988
rect 26056 9868 26108 9920
rect 57888 9868 57940 9920
rect 20214 9766 20266 9818
rect 20278 9766 20330 9818
rect 20342 9766 20394 9818
rect 20406 9766 20458 9818
rect 20470 9766 20522 9818
rect 39478 9766 39530 9818
rect 39542 9766 39594 9818
rect 39606 9766 39658 9818
rect 39670 9766 39722 9818
rect 39734 9766 39786 9818
rect 26884 9664 26936 9716
rect 24952 9639 25004 9648
rect 24952 9605 24961 9639
rect 24961 9605 24995 9639
rect 24995 9605 25004 9639
rect 24952 9596 25004 9605
rect 26056 9639 26108 9648
rect 26056 9605 26065 9639
rect 26065 9605 26099 9639
rect 26099 9605 26108 9639
rect 26056 9596 26108 9605
rect 27344 9639 27396 9648
rect 27344 9605 27353 9639
rect 27353 9605 27387 9639
rect 27387 9605 27396 9639
rect 27344 9596 27396 9605
rect 50344 9528 50396 9580
rect 25044 9503 25096 9512
rect 25044 9469 25053 9503
rect 25053 9469 25087 9503
rect 25087 9469 25096 9503
rect 25044 9460 25096 9469
rect 27436 9503 27488 9512
rect 27436 9469 27445 9503
rect 27445 9469 27479 9503
rect 27479 9469 27488 9503
rect 27436 9460 27488 9469
rect 23756 9324 23808 9376
rect 27344 9392 27396 9444
rect 58072 9367 58124 9376
rect 58072 9333 58081 9367
rect 58081 9333 58115 9367
rect 58115 9333 58124 9367
rect 58072 9324 58124 9333
rect 10582 9222 10634 9274
rect 10646 9222 10698 9274
rect 10710 9222 10762 9274
rect 10774 9222 10826 9274
rect 10838 9222 10890 9274
rect 29846 9222 29898 9274
rect 29910 9222 29962 9274
rect 29974 9222 30026 9274
rect 30038 9222 30090 9274
rect 30102 9222 30154 9274
rect 49110 9222 49162 9274
rect 49174 9222 49226 9274
rect 49238 9222 49290 9274
rect 49302 9222 49354 9274
rect 49366 9222 49418 9274
rect 10508 9120 10560 9172
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 27988 9120 28040 9172
rect 1400 8984 1452 9036
rect 23756 8984 23808 9036
rect 27344 8984 27396 9036
rect 9772 8916 9824 8968
rect 10968 8916 11020 8968
rect 12532 8916 12584 8968
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 22560 8959 22612 8968
rect 22560 8925 22569 8959
rect 22569 8925 22603 8959
rect 22603 8925 22612 8959
rect 22560 8916 22612 8925
rect 23204 8916 23256 8968
rect 27804 8916 27856 8968
rect 50344 8916 50396 8968
rect 50436 8916 50488 8968
rect 26516 8891 26568 8900
rect 26516 8857 26525 8891
rect 26525 8857 26559 8891
rect 26559 8857 26568 8891
rect 26516 8848 26568 8857
rect 22468 8780 22520 8832
rect 22652 8823 22704 8832
rect 22652 8789 22661 8823
rect 22661 8789 22695 8823
rect 22695 8789 22704 8823
rect 22652 8780 22704 8789
rect 27620 8823 27672 8832
rect 27620 8789 27629 8823
rect 27629 8789 27663 8823
rect 27663 8789 27672 8823
rect 58072 8823 58124 8832
rect 27620 8780 27672 8789
rect 58072 8789 58081 8823
rect 58081 8789 58115 8823
rect 58115 8789 58124 8823
rect 58072 8780 58124 8789
rect 20214 8678 20266 8730
rect 20278 8678 20330 8730
rect 20342 8678 20394 8730
rect 20406 8678 20458 8730
rect 20470 8678 20522 8730
rect 39478 8678 39530 8730
rect 39542 8678 39594 8730
rect 39606 8678 39658 8730
rect 39670 8678 39722 8730
rect 39734 8678 39786 8730
rect 9404 8576 9456 8628
rect 23204 8619 23256 8628
rect 23204 8585 23213 8619
rect 23213 8585 23247 8619
rect 23247 8585 23256 8619
rect 23204 8576 23256 8585
rect 23572 8619 23624 8628
rect 23572 8585 23581 8619
rect 23581 8585 23615 8619
rect 23615 8585 23624 8619
rect 23572 8576 23624 8585
rect 9864 8440 9916 8492
rect 15108 8440 15160 8492
rect 22468 8483 22520 8492
rect 22468 8449 22477 8483
rect 22477 8449 22511 8483
rect 22511 8449 22520 8483
rect 22468 8440 22520 8449
rect 20996 8372 21048 8424
rect 23664 8415 23716 8424
rect 23664 8381 23673 8415
rect 23673 8381 23707 8415
rect 23707 8381 23716 8415
rect 23664 8372 23716 8381
rect 23756 8415 23808 8424
rect 23756 8381 23765 8415
rect 23765 8381 23799 8415
rect 23799 8381 23808 8415
rect 23756 8372 23808 8381
rect 50436 8508 50488 8560
rect 57888 8304 57940 8356
rect 12992 8236 13044 8288
rect 10582 8134 10634 8186
rect 10646 8134 10698 8186
rect 10710 8134 10762 8186
rect 10774 8134 10826 8186
rect 10838 8134 10890 8186
rect 29846 8134 29898 8186
rect 29910 8134 29962 8186
rect 29974 8134 30026 8186
rect 30038 8134 30090 8186
rect 30102 8134 30154 8186
rect 49110 8134 49162 8186
rect 49174 8134 49226 8186
rect 49238 8134 49290 8186
rect 49302 8134 49354 8186
rect 49366 8134 49418 8186
rect 9864 8075 9916 8084
rect 9864 8041 9873 8075
rect 9873 8041 9907 8075
rect 9907 8041 9916 8075
rect 9864 8032 9916 8041
rect 10968 8075 11020 8084
rect 10968 8041 10977 8075
rect 10977 8041 11011 8075
rect 11011 8041 11020 8075
rect 10968 8032 11020 8041
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 14280 8032 14332 8084
rect 20996 8075 21048 8084
rect 20996 8041 21005 8075
rect 21005 8041 21039 8075
rect 21039 8041 21048 8075
rect 20996 8032 21048 8041
rect 10876 8007 10928 8016
rect 10876 7973 10885 8007
rect 10885 7973 10919 8007
rect 10919 7973 10928 8007
rect 10876 7964 10928 7973
rect 12348 8007 12400 8016
rect 12348 7973 12357 8007
rect 12357 7973 12391 8007
rect 12391 7973 12400 8007
rect 12348 7964 12400 7973
rect 13360 8007 13412 8016
rect 13360 7973 13369 8007
rect 13369 7973 13403 8007
rect 13403 7973 13412 8007
rect 13360 7964 13412 7973
rect 9864 7896 9916 7948
rect 12992 7939 13044 7948
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 12992 7905 13001 7939
rect 13001 7905 13035 7939
rect 13035 7905 13044 7939
rect 12992 7896 13044 7905
rect 20812 7871 20864 7880
rect 9404 7828 9456 7837
rect 20812 7837 20821 7871
rect 20821 7837 20855 7871
rect 20855 7837 20864 7871
rect 20812 7828 20864 7837
rect 15108 7760 15160 7812
rect 26516 7760 26568 7812
rect 19984 7735 20036 7744
rect 19984 7701 19993 7735
rect 19993 7701 20027 7735
rect 20027 7701 20036 7735
rect 19984 7692 20036 7701
rect 57520 7735 57572 7744
rect 57520 7701 57529 7735
rect 57529 7701 57563 7735
rect 57563 7701 57572 7735
rect 57520 7692 57572 7701
rect 58072 7735 58124 7744
rect 58072 7701 58081 7735
rect 58081 7701 58115 7735
rect 58115 7701 58124 7735
rect 58072 7692 58124 7701
rect 20214 7590 20266 7642
rect 20278 7590 20330 7642
rect 20342 7590 20394 7642
rect 20406 7590 20458 7642
rect 20470 7590 20522 7642
rect 39478 7590 39530 7642
rect 39542 7590 39594 7642
rect 39606 7590 39658 7642
rect 39670 7590 39722 7642
rect 39734 7590 39786 7642
rect 9772 7488 9824 7540
rect 10876 7488 10928 7540
rect 57980 7488 58032 7540
rect 9404 7463 9456 7472
rect 9404 7429 9413 7463
rect 9413 7429 9447 7463
rect 9447 7429 9456 7463
rect 9404 7420 9456 7429
rect 19248 7420 19300 7472
rect 20076 7420 20128 7472
rect 20720 7420 20772 7472
rect 57428 7352 57480 7404
rect 19248 7284 19300 7336
rect 9772 7259 9824 7268
rect 9772 7225 9781 7259
rect 9781 7225 9815 7259
rect 9815 7225 9824 7259
rect 9772 7216 9824 7225
rect 17776 7216 17828 7268
rect 19984 7284 20036 7336
rect 20812 7216 20864 7268
rect 19616 7148 19668 7200
rect 57428 7191 57480 7200
rect 57428 7157 57437 7191
rect 57437 7157 57471 7191
rect 57471 7157 57480 7191
rect 57428 7148 57480 7157
rect 58072 7191 58124 7200
rect 58072 7157 58081 7191
rect 58081 7157 58115 7191
rect 58115 7157 58124 7191
rect 58072 7148 58124 7157
rect 10582 7046 10634 7098
rect 10646 7046 10698 7098
rect 10710 7046 10762 7098
rect 10774 7046 10826 7098
rect 10838 7046 10890 7098
rect 29846 7046 29898 7098
rect 29910 7046 29962 7098
rect 29974 7046 30026 7098
rect 30038 7046 30090 7098
rect 30102 7046 30154 7098
rect 49110 7046 49162 7098
rect 49174 7046 49226 7098
rect 49238 7046 49290 7098
rect 49302 7046 49354 7098
rect 49366 7046 49418 7098
rect 16580 6808 16632 6860
rect 17776 6808 17828 6860
rect 16396 6783 16448 6792
rect 16396 6749 16405 6783
rect 16405 6749 16439 6783
rect 16439 6749 16448 6783
rect 16396 6740 16448 6749
rect 17868 6783 17920 6792
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 50344 6740 50396 6792
rect 16028 6647 16080 6656
rect 16028 6613 16037 6647
rect 16037 6613 16071 6647
rect 16071 6613 16080 6647
rect 16028 6604 16080 6613
rect 16672 6604 16724 6656
rect 17500 6647 17552 6656
rect 17500 6613 17509 6647
rect 17509 6613 17543 6647
rect 17543 6613 17552 6647
rect 17500 6604 17552 6613
rect 17868 6604 17920 6656
rect 57520 6604 57572 6656
rect 58072 6647 58124 6656
rect 58072 6613 58081 6647
rect 58081 6613 58115 6647
rect 58115 6613 58124 6647
rect 58072 6604 58124 6613
rect 20214 6502 20266 6554
rect 20278 6502 20330 6554
rect 20342 6502 20394 6554
rect 20406 6502 20458 6554
rect 20470 6502 20522 6554
rect 39478 6502 39530 6554
rect 39542 6502 39594 6554
rect 39606 6502 39658 6554
rect 39670 6502 39722 6554
rect 39734 6502 39786 6554
rect 15016 6400 15068 6452
rect 16028 6332 16080 6384
rect 15660 6239 15712 6248
rect 15660 6205 15669 6239
rect 15669 6205 15703 6239
rect 15703 6205 15712 6239
rect 15660 6196 15712 6205
rect 16580 6196 16632 6248
rect 17500 6264 17552 6316
rect 57428 6196 57480 6248
rect 50344 6060 50396 6112
rect 58072 6103 58124 6112
rect 58072 6069 58081 6103
rect 58081 6069 58115 6103
rect 58115 6069 58124 6103
rect 58072 6060 58124 6069
rect 10582 5958 10634 6010
rect 10646 5958 10698 6010
rect 10710 5958 10762 6010
rect 10774 5958 10826 6010
rect 10838 5958 10890 6010
rect 29846 5958 29898 6010
rect 29910 5958 29962 6010
rect 29974 5958 30026 6010
rect 30038 5958 30090 6010
rect 30102 5958 30154 6010
rect 49110 5958 49162 6010
rect 49174 5958 49226 6010
rect 49238 5958 49290 6010
rect 49302 5958 49354 6010
rect 49366 5958 49418 6010
rect 55772 5856 55824 5908
rect 57980 5831 58032 5840
rect 57980 5797 57989 5831
rect 57989 5797 58023 5831
rect 58023 5797 58032 5831
rect 57980 5788 58032 5797
rect 56876 5627 56928 5636
rect 56876 5593 56885 5627
rect 56885 5593 56919 5627
rect 56919 5593 56928 5627
rect 56876 5584 56928 5593
rect 57796 5627 57848 5636
rect 57796 5593 57805 5627
rect 57805 5593 57839 5627
rect 57839 5593 57848 5627
rect 57796 5584 57848 5593
rect 20214 5414 20266 5466
rect 20278 5414 20330 5466
rect 20342 5414 20394 5466
rect 20406 5414 20458 5466
rect 20470 5414 20522 5466
rect 39478 5414 39530 5466
rect 39542 5414 39594 5466
rect 39606 5414 39658 5466
rect 39670 5414 39722 5466
rect 39734 5414 39786 5466
rect 56508 5176 56560 5228
rect 56784 4972 56836 5024
rect 10582 4870 10634 4922
rect 10646 4870 10698 4922
rect 10710 4870 10762 4922
rect 10774 4870 10826 4922
rect 10838 4870 10890 4922
rect 29846 4870 29898 4922
rect 29910 4870 29962 4922
rect 29974 4870 30026 4922
rect 30038 4870 30090 4922
rect 30102 4870 30154 4922
rect 49110 4870 49162 4922
rect 49174 4870 49226 4922
rect 49238 4870 49290 4922
rect 49302 4870 49354 4922
rect 49366 4870 49418 4922
rect 57612 4675 57664 4684
rect 57612 4641 57621 4675
rect 57621 4641 57655 4675
rect 57655 4641 57664 4675
rect 57612 4632 57664 4641
rect 59176 4564 59228 4616
rect 56508 4539 56560 4548
rect 56508 4505 56517 4539
rect 56517 4505 56551 4539
rect 56551 4505 56560 4539
rect 56508 4496 56560 4505
rect 56600 4471 56652 4480
rect 56600 4437 56609 4471
rect 56609 4437 56643 4471
rect 56643 4437 56652 4471
rect 56600 4428 56652 4437
rect 20214 4326 20266 4378
rect 20278 4326 20330 4378
rect 20342 4326 20394 4378
rect 20406 4326 20458 4378
rect 20470 4326 20522 4378
rect 39478 4326 39530 4378
rect 39542 4326 39594 4378
rect 39606 4326 39658 4378
rect 39670 4326 39722 4378
rect 39734 4326 39786 4378
rect 56048 4199 56100 4208
rect 56048 4165 56057 4199
rect 56057 4165 56091 4199
rect 56091 4165 56100 4199
rect 56048 4156 56100 4165
rect 57152 4156 57204 4208
rect 2136 4088 2188 4140
rect 3792 4088 3844 4140
rect 6552 4088 6604 4140
rect 7932 4131 7984 4140
rect 7932 4097 7941 4131
rect 7941 4097 7975 4131
rect 7975 4097 7984 4131
rect 7932 4088 7984 4097
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 3976 4020 4028 4072
rect 6828 4020 6880 4072
rect 7288 4020 7340 4072
rect 9864 3952 9916 4004
rect 6736 3884 6788 3936
rect 55680 3884 55732 3936
rect 57060 3927 57112 3936
rect 57060 3893 57069 3927
rect 57069 3893 57103 3927
rect 57103 3893 57112 3927
rect 57060 3884 57112 3893
rect 10582 3782 10634 3834
rect 10646 3782 10698 3834
rect 10710 3782 10762 3834
rect 10774 3782 10826 3834
rect 10838 3782 10890 3834
rect 29846 3782 29898 3834
rect 29910 3782 29962 3834
rect 29974 3782 30026 3834
rect 30038 3782 30090 3834
rect 30102 3782 30154 3834
rect 49110 3782 49162 3834
rect 49174 3782 49226 3834
rect 49238 3782 49290 3834
rect 49302 3782 49354 3834
rect 49366 3782 49418 3834
rect 2964 3680 3016 3732
rect 4068 3655 4120 3664
rect 4068 3621 4077 3655
rect 4077 3621 4111 3655
rect 4111 3621 4120 3655
rect 4068 3612 4120 3621
rect 3884 3544 3936 3596
rect 7472 3612 7524 3664
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 5356 3544 5408 3596
rect 4160 3476 4212 3528
rect 4988 3476 5040 3528
rect 57060 3544 57112 3596
rect 57704 3544 57756 3596
rect 3792 3451 3844 3460
rect 3792 3417 3801 3451
rect 3801 3417 3835 3451
rect 3835 3417 3844 3451
rect 3792 3408 3844 3417
rect 2780 3340 2832 3392
rect 7656 3476 7708 3528
rect 9956 3476 10008 3528
rect 8392 3408 8444 3460
rect 10968 3476 11020 3528
rect 40132 3476 40184 3528
rect 56968 3476 57020 3528
rect 55772 3408 55824 3460
rect 56508 3451 56560 3460
rect 56508 3417 56517 3451
rect 56517 3417 56551 3451
rect 56551 3417 56560 3451
rect 56508 3408 56560 3417
rect 6368 3340 6420 3392
rect 7288 3383 7340 3392
rect 7288 3349 7297 3383
rect 7297 3349 7331 3383
rect 7331 3349 7340 3383
rect 7288 3340 7340 3349
rect 7932 3340 7984 3392
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 10784 3340 10836 3392
rect 11520 3340 11572 3392
rect 48412 3340 48464 3392
rect 56784 3340 56836 3392
rect 20214 3238 20266 3290
rect 20278 3238 20330 3290
rect 20342 3238 20394 3290
rect 20406 3238 20458 3290
rect 20470 3238 20522 3290
rect 39478 3238 39530 3290
rect 39542 3238 39594 3290
rect 39606 3238 39658 3290
rect 39670 3238 39722 3290
rect 39734 3238 39786 3290
rect 3976 3179 4028 3188
rect 3976 3145 3985 3179
rect 3985 3145 4019 3179
rect 4019 3145 4028 3179
rect 3976 3136 4028 3145
rect 4988 3179 5040 3188
rect 4988 3145 4997 3179
rect 4997 3145 5031 3179
rect 5031 3145 5040 3179
rect 4988 3136 5040 3145
rect 5172 3136 5224 3188
rect 6828 3179 6880 3188
rect 3240 3068 3292 3120
rect 3792 3068 3844 3120
rect 6368 3111 6420 3120
rect 6368 3077 6377 3111
rect 6377 3077 6411 3111
rect 6411 3077 6420 3111
rect 6368 3068 6420 3077
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 7656 3179 7708 3188
rect 7656 3145 7665 3179
rect 7665 3145 7699 3179
rect 7699 3145 7708 3179
rect 7656 3136 7708 3145
rect 10968 3136 11020 3188
rect 13360 3136 13412 3188
rect 48412 3136 48464 3188
rect 55680 3179 55732 3188
rect 55680 3145 55689 3179
rect 55689 3145 55723 3179
rect 55723 3145 55732 3179
rect 55680 3136 55732 3145
rect 9128 3068 9180 3120
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 5632 3000 5684 3009
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 8392 3000 8444 3052
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 10876 3000 10928 3052
rect 12348 3000 12400 3052
rect 7104 2932 7156 2984
rect 9680 2975 9732 2984
rect 3884 2907 3936 2916
rect 3884 2873 3893 2907
rect 3893 2873 3927 2907
rect 3927 2873 3936 2907
rect 3884 2864 3936 2873
rect 4896 2907 4948 2916
rect 4896 2873 4905 2907
rect 4905 2873 4939 2907
rect 4939 2873 4948 2907
rect 4896 2864 4948 2873
rect 5356 2864 5408 2916
rect 6736 2907 6788 2916
rect 6736 2873 6745 2907
rect 6745 2873 6779 2907
rect 6779 2873 6788 2907
rect 6736 2864 6788 2873
rect 9680 2941 9689 2975
rect 9689 2941 9723 2975
rect 9723 2941 9732 2975
rect 9680 2932 9732 2941
rect 10784 2932 10836 2984
rect 56600 3068 56652 3120
rect 49516 3043 49568 3052
rect 49516 3009 49525 3043
rect 49525 3009 49559 3043
rect 49559 3009 49568 3043
rect 49516 3000 49568 3009
rect 53840 3043 53892 3052
rect 53840 3009 53849 3043
rect 53849 3009 53883 3043
rect 53883 3009 53892 3043
rect 53840 3000 53892 3009
rect 55588 3043 55640 3052
rect 55588 3009 55597 3043
rect 55597 3009 55631 3043
rect 55631 3009 55640 3043
rect 55588 3000 55640 3009
rect 56692 3043 56744 3052
rect 56692 3009 56701 3043
rect 56701 3009 56735 3043
rect 56735 3009 56744 3043
rect 56692 3000 56744 3009
rect 48964 2932 49016 2984
rect 53472 2932 53524 2984
rect 56324 2932 56376 2984
rect 3516 2796 3568 2848
rect 5540 2796 5592 2848
rect 10416 2796 10468 2848
rect 13176 2796 13228 2848
rect 14096 2796 14148 2848
rect 10582 2694 10634 2746
rect 10646 2694 10698 2746
rect 10710 2694 10762 2746
rect 10774 2694 10826 2746
rect 10838 2694 10890 2746
rect 29846 2694 29898 2746
rect 29910 2694 29962 2746
rect 29974 2694 30026 2746
rect 30038 2694 30090 2746
rect 30102 2694 30154 2746
rect 49110 2694 49162 2746
rect 49174 2694 49226 2746
rect 49238 2694 49290 2746
rect 49302 2694 49354 2746
rect 49366 2694 49418 2746
rect 3240 2635 3292 2644
rect 3240 2601 3249 2635
rect 3249 2601 3283 2635
rect 3283 2601 3292 2635
rect 3240 2592 3292 2601
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 5632 2592 5684 2644
rect 16672 2635 16724 2644
rect 5172 2524 5224 2576
rect 2780 2388 2832 2440
rect 3792 2388 3844 2440
rect 4068 2456 4120 2508
rect 6368 2524 6420 2576
rect 9220 2524 9272 2576
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 5540 2431 5592 2440
rect 4896 2388 4948 2397
rect 5540 2397 5549 2431
rect 5549 2397 5583 2431
rect 5583 2397 5592 2431
rect 5540 2388 5592 2397
rect 6644 2388 6696 2440
rect 7932 2431 7984 2440
rect 7104 2320 7156 2372
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 9680 2456 9732 2508
rect 9956 2499 10008 2508
rect 9956 2465 9965 2499
rect 9965 2465 9999 2499
rect 9999 2465 10008 2499
rect 9956 2456 10008 2465
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 10416 2431 10468 2440
rect 10416 2397 10425 2431
rect 10425 2397 10459 2431
rect 10459 2397 10468 2431
rect 10416 2388 10468 2397
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 15660 2524 15712 2576
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 17868 2635 17920 2644
rect 17868 2601 17877 2635
rect 17877 2601 17911 2635
rect 17911 2601 17920 2635
rect 17868 2592 17920 2601
rect 19248 2635 19300 2644
rect 19248 2601 19257 2635
rect 19257 2601 19291 2635
rect 19291 2601 19300 2635
rect 19248 2592 19300 2601
rect 20720 2635 20772 2644
rect 20720 2601 20729 2635
rect 20729 2601 20763 2635
rect 20763 2601 20772 2635
rect 20720 2592 20772 2601
rect 22652 2592 22704 2644
rect 23664 2592 23716 2644
rect 25044 2592 25096 2644
rect 27436 2592 27488 2644
rect 27620 2592 27672 2644
rect 29552 2635 29604 2644
rect 29552 2601 29561 2635
rect 29561 2601 29595 2635
rect 29595 2601 29604 2635
rect 29552 2592 29604 2601
rect 30748 2635 30800 2644
rect 30748 2601 30757 2635
rect 30757 2601 30791 2635
rect 30791 2601 30800 2635
rect 30748 2592 30800 2601
rect 32128 2635 32180 2644
rect 32128 2601 32137 2635
rect 32137 2601 32171 2635
rect 32171 2601 32180 2635
rect 32128 2592 32180 2601
rect 33600 2635 33652 2644
rect 33600 2601 33609 2635
rect 33609 2601 33643 2635
rect 33643 2601 33652 2635
rect 33600 2592 33652 2601
rect 34980 2635 35032 2644
rect 34980 2601 34989 2635
rect 34989 2601 35023 2635
rect 35023 2601 35032 2635
rect 34980 2592 35032 2601
rect 36360 2592 36412 2644
rect 37740 2592 37792 2644
rect 39856 2635 39908 2644
rect 39856 2601 39865 2635
rect 39865 2601 39899 2635
rect 39899 2601 39908 2635
rect 39856 2592 39908 2601
rect 41604 2592 41656 2644
rect 42340 2592 42392 2644
rect 43536 2635 43588 2644
rect 43536 2601 43545 2635
rect 43545 2601 43579 2635
rect 43579 2601 43588 2635
rect 43536 2592 43588 2601
rect 45008 2635 45060 2644
rect 45008 2601 45017 2635
rect 45017 2601 45051 2635
rect 45051 2601 45060 2635
rect 45008 2592 45060 2601
rect 46296 2592 46348 2644
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 14924 2388 14976 2440
rect 16304 2388 16356 2440
rect 17776 2388 17828 2440
rect 19156 2388 19208 2440
rect 20628 2388 20680 2440
rect 22008 2388 22060 2440
rect 23480 2388 23532 2440
rect 24860 2388 24912 2440
rect 26332 2388 26384 2440
rect 27712 2388 27764 2440
rect 29184 2388 29236 2440
rect 30656 2388 30708 2440
rect 32036 2388 32088 2440
rect 33508 2388 33560 2440
rect 34888 2388 34940 2440
rect 36360 2388 36412 2440
rect 37740 2388 37792 2440
rect 39212 2388 39264 2440
rect 40592 2388 40644 2440
rect 42064 2388 42116 2440
rect 43444 2388 43496 2440
rect 44916 2388 44968 2440
rect 664 2252 716 2304
rect 2044 2252 2096 2304
rect 5172 2252 5224 2304
rect 7748 2252 7800 2304
rect 10692 2252 10744 2304
rect 12072 2252 12124 2304
rect 13452 2252 13504 2304
rect 48044 2456 48096 2508
rect 50988 2499 51040 2508
rect 50988 2465 50997 2499
rect 50997 2465 51031 2499
rect 51031 2465 51040 2499
rect 50988 2456 51040 2465
rect 52368 2456 52420 2508
rect 55496 2456 55548 2508
rect 46296 2388 46348 2440
rect 47768 2388 47820 2440
rect 50620 2388 50672 2440
rect 52000 2388 52052 2440
rect 54852 2388 54904 2440
rect 55128 2320 55180 2372
rect 56968 2363 57020 2372
rect 56968 2329 56977 2363
rect 56977 2329 57011 2363
rect 57011 2329 57020 2363
rect 56968 2320 57020 2329
rect 20214 2150 20266 2202
rect 20278 2150 20330 2202
rect 20342 2150 20394 2202
rect 20406 2150 20458 2202
rect 20470 2150 20522 2202
rect 39478 2150 39530 2202
rect 39542 2150 39594 2202
rect 39606 2150 39658 2202
rect 39670 2150 39722 2202
rect 39734 2150 39786 2202
<< metal2 >>
rect 662 21298 718 22000
rect 2042 21298 2098 22000
rect 662 21270 1072 21298
rect 662 21200 718 21270
rect 1044 19514 1072 21270
rect 2042 21270 2360 21298
rect 2042 21200 2098 21270
rect 2332 19514 2360 21270
rect 3514 21200 3570 22000
rect 4894 21298 4950 22000
rect 6366 21298 6422 22000
rect 7746 21298 7802 22000
rect 9218 21298 9274 22000
rect 10598 21298 10654 22000
rect 12070 21298 12126 22000
rect 4894 21270 5212 21298
rect 4894 21200 4950 21270
rect 3528 19514 3556 21200
rect 5184 19514 5212 21270
rect 6366 21270 6684 21298
rect 6366 21200 6422 21270
rect 6656 19514 6684 21270
rect 7746 21270 8064 21298
rect 7746 21200 7802 21270
rect 8036 19514 8064 21270
rect 9218 21270 9536 21298
rect 9218 21200 9274 21270
rect 9508 19514 9536 21270
rect 10598 21270 10916 21298
rect 10598 21200 10654 21270
rect 10888 19514 10916 21270
rect 12070 21270 12388 21298
rect 12070 21200 12126 21270
rect 12360 19514 12388 21270
rect 13450 21200 13506 22000
rect 14922 21200 14978 22000
rect 16302 21200 16358 22000
rect 17774 21200 17830 22000
rect 19154 21200 19210 22000
rect 20626 21200 20682 22000
rect 22006 21200 22062 22000
rect 23478 21298 23534 22000
rect 24858 21298 24914 22000
rect 23478 21270 23796 21298
rect 23478 21200 23534 21270
rect 13464 19514 13492 21200
rect 1032 19508 1084 19514
rect 1032 19450 1084 19456
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 14936 19378 14964 21200
rect 16316 19378 16344 21200
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 2136 19372 2188 19378
rect 2136 19314 2188 19320
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 16304 19372 16356 19378
rect 16304 19314 16356 19320
rect 1412 9042 1440 19314
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 2148 4146 2176 19314
rect 3804 4146 3832 19314
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 2976 3738 3004 4014
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2792 2446 2820 3334
rect 3804 3126 3832 3402
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3252 2650 3280 3062
rect 3896 2922 3924 3538
rect 3988 3194 4016 4014
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 664 2304 716 2310
rect 664 2246 716 2252
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 676 800 704 2246
rect 2056 800 2084 2246
rect 3528 800 3556 2790
rect 3896 2530 3924 2858
rect 3804 2502 3924 2530
rect 4080 2514 4108 3606
rect 5092 3602 5120 19314
rect 6564 4146 6592 19314
rect 7944 4146 7972 19314
rect 9416 8634 9444 19314
rect 10520 9178 10548 19314
rect 10582 19068 10890 19088
rect 10582 19066 10588 19068
rect 10644 19066 10668 19068
rect 10724 19066 10748 19068
rect 10804 19066 10828 19068
rect 10884 19066 10890 19068
rect 10644 19014 10646 19066
rect 10826 19014 10828 19066
rect 10582 19012 10588 19014
rect 10644 19012 10668 19014
rect 10724 19012 10748 19014
rect 10804 19012 10828 19014
rect 10884 19012 10890 19014
rect 10582 18992 10890 19012
rect 10582 17980 10890 18000
rect 10582 17978 10588 17980
rect 10644 17978 10668 17980
rect 10724 17978 10748 17980
rect 10804 17978 10828 17980
rect 10884 17978 10890 17980
rect 10644 17926 10646 17978
rect 10826 17926 10828 17978
rect 10582 17924 10588 17926
rect 10644 17924 10668 17926
rect 10724 17924 10748 17926
rect 10804 17924 10828 17926
rect 10884 17924 10890 17926
rect 10582 17904 10890 17924
rect 10582 16892 10890 16912
rect 10582 16890 10588 16892
rect 10644 16890 10668 16892
rect 10724 16890 10748 16892
rect 10804 16890 10828 16892
rect 10884 16890 10890 16892
rect 10644 16838 10646 16890
rect 10826 16838 10828 16890
rect 10582 16836 10588 16838
rect 10644 16836 10668 16838
rect 10724 16836 10748 16838
rect 10804 16836 10828 16838
rect 10884 16836 10890 16838
rect 10582 16816 10890 16836
rect 10582 15804 10890 15824
rect 10582 15802 10588 15804
rect 10644 15802 10668 15804
rect 10724 15802 10748 15804
rect 10804 15802 10828 15804
rect 10884 15802 10890 15804
rect 10644 15750 10646 15802
rect 10826 15750 10828 15802
rect 10582 15748 10588 15750
rect 10644 15748 10668 15750
rect 10724 15748 10748 15750
rect 10804 15748 10828 15750
rect 10884 15748 10890 15750
rect 10582 15728 10890 15748
rect 10582 14716 10890 14736
rect 10582 14714 10588 14716
rect 10644 14714 10668 14716
rect 10724 14714 10748 14716
rect 10804 14714 10828 14716
rect 10884 14714 10890 14716
rect 10644 14662 10646 14714
rect 10826 14662 10828 14714
rect 10582 14660 10588 14662
rect 10644 14660 10668 14662
rect 10724 14660 10748 14662
rect 10804 14660 10828 14662
rect 10884 14660 10890 14662
rect 10582 14640 10890 14660
rect 10582 13628 10890 13648
rect 10582 13626 10588 13628
rect 10644 13626 10668 13628
rect 10724 13626 10748 13628
rect 10804 13626 10828 13628
rect 10884 13626 10890 13628
rect 10644 13574 10646 13626
rect 10826 13574 10828 13626
rect 10582 13572 10588 13574
rect 10644 13572 10668 13574
rect 10724 13572 10748 13574
rect 10804 13572 10828 13574
rect 10884 13572 10890 13574
rect 10582 13552 10890 13572
rect 10582 12540 10890 12560
rect 10582 12538 10588 12540
rect 10644 12538 10668 12540
rect 10724 12538 10748 12540
rect 10804 12538 10828 12540
rect 10884 12538 10890 12540
rect 10644 12486 10646 12538
rect 10826 12486 10828 12538
rect 10582 12484 10588 12486
rect 10644 12484 10668 12486
rect 10724 12484 10748 12486
rect 10804 12484 10828 12486
rect 10884 12484 10890 12486
rect 10582 12464 10890 12484
rect 10582 11452 10890 11472
rect 10582 11450 10588 11452
rect 10644 11450 10668 11452
rect 10724 11450 10748 11452
rect 10804 11450 10828 11452
rect 10884 11450 10890 11452
rect 10644 11398 10646 11450
rect 10826 11398 10828 11450
rect 10582 11396 10588 11398
rect 10644 11396 10668 11398
rect 10724 11396 10748 11398
rect 10804 11396 10828 11398
rect 10884 11396 10890 11398
rect 10582 11376 10890 11396
rect 10582 10364 10890 10384
rect 10582 10362 10588 10364
rect 10644 10362 10668 10364
rect 10724 10362 10748 10364
rect 10804 10362 10828 10364
rect 10884 10362 10890 10364
rect 10644 10310 10646 10362
rect 10826 10310 10828 10362
rect 10582 10308 10588 10310
rect 10644 10308 10668 10310
rect 10724 10308 10748 10310
rect 10804 10308 10828 10310
rect 10884 10308 10890 10310
rect 10582 10288 10890 10308
rect 10582 9276 10890 9296
rect 10582 9274 10588 9276
rect 10644 9274 10668 9276
rect 10724 9274 10748 9276
rect 10804 9274 10828 9276
rect 10884 9274 10890 9276
rect 10644 9222 10646 9274
rect 10826 9222 10828 9274
rect 10582 9220 10588 9222
rect 10644 9220 10668 9222
rect 10724 9220 10748 9222
rect 10804 9220 10828 9222
rect 10884 9220 10890 9222
rect 10582 9200 10890 9220
rect 12084 9178 12112 19314
rect 14108 9178 14136 19314
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9416 7478 9444 7822
rect 9784 7546 9812 8910
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9876 8090 9904 8434
rect 10582 8188 10890 8208
rect 10582 8186 10588 8188
rect 10644 8186 10668 8188
rect 10724 8186 10748 8188
rect 10804 8186 10828 8188
rect 10884 8186 10890 8188
rect 10644 8134 10646 8186
rect 10826 8134 10828 8186
rect 10582 8132 10588 8134
rect 10644 8132 10668 8134
rect 10724 8132 10748 8134
rect 10804 8132 10828 8134
rect 10884 8132 10890 8134
rect 10582 8112 10890 8132
rect 10980 8090 11008 8910
rect 12544 8090 12572 8910
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4172 2650 4200 3470
rect 5000 3194 5028 3470
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4068 2508 4120 2514
rect 3804 2446 3832 2502
rect 4068 2450 4120 2456
rect 4908 2446 4936 2858
rect 5184 2582 5212 3130
rect 5368 2922 5396 3538
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6380 3126 6408 3334
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5172 2576 5224 2582
rect 5172 2518 5224 2524
rect 5552 2446 5580 2790
rect 5644 2650 5672 2994
rect 6748 2922 6776 3878
rect 6840 3194 6868 4014
rect 7300 3398 7328 4014
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7484 3058 7512 3606
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 3194 7696 3470
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 6368 2576 6420 2582
rect 6748 2530 6776 2858
rect 6368 2518 6420 2524
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 4908 870 5028 898
rect 4908 800 4936 870
rect 662 0 718 800
rect 2042 0 2098 800
rect 3514 0 3570 800
rect 4894 0 4950 800
rect 5000 762 5028 870
rect 5184 762 5212 2246
rect 6380 800 6408 2518
rect 6656 2502 6776 2530
rect 6656 2446 6684 2502
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 7116 2378 7144 2926
rect 7944 2446 7972 3334
rect 8404 3058 8432 3402
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9140 3126 9168 3334
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 800 7788 2246
rect 9232 800 9260 2518
rect 9692 2514 9720 2926
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9784 2446 9812 7210
rect 9876 4010 9904 7890
rect 10888 7546 10916 7958
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10888 7426 10916 7482
rect 10888 7398 11008 7426
rect 10582 7100 10890 7120
rect 10582 7098 10588 7100
rect 10644 7098 10668 7100
rect 10724 7098 10748 7100
rect 10804 7098 10828 7100
rect 10884 7098 10890 7100
rect 10644 7046 10646 7098
rect 10826 7046 10828 7098
rect 10582 7044 10588 7046
rect 10644 7044 10668 7046
rect 10724 7044 10748 7046
rect 10804 7044 10828 7046
rect 10884 7044 10890 7046
rect 10582 7024 10890 7044
rect 10582 6012 10890 6032
rect 10582 6010 10588 6012
rect 10644 6010 10668 6012
rect 10724 6010 10748 6012
rect 10804 6010 10828 6012
rect 10884 6010 10890 6012
rect 10644 5958 10646 6010
rect 10826 5958 10828 6010
rect 10582 5956 10588 5958
rect 10644 5956 10668 5958
rect 10724 5956 10748 5958
rect 10804 5956 10828 5958
rect 10884 5956 10890 5958
rect 10582 5936 10890 5956
rect 10582 4924 10890 4944
rect 10582 4922 10588 4924
rect 10644 4922 10668 4924
rect 10724 4922 10748 4924
rect 10804 4922 10828 4924
rect 10884 4922 10890 4924
rect 10644 4870 10646 4922
rect 10826 4870 10828 4922
rect 10582 4868 10588 4870
rect 10644 4868 10668 4870
rect 10724 4868 10748 4870
rect 10804 4868 10828 4870
rect 10884 4868 10890 4870
rect 10582 4848 10890 4868
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9876 3058 9904 3946
rect 10582 3836 10890 3856
rect 10582 3834 10588 3836
rect 10644 3834 10668 3836
rect 10724 3834 10748 3836
rect 10804 3834 10828 3836
rect 10884 3834 10890 3836
rect 10644 3782 10646 3834
rect 10826 3782 10828 3834
rect 10582 3780 10588 3782
rect 10644 3780 10668 3782
rect 10724 3780 10748 3782
rect 10804 3780 10828 3782
rect 10884 3780 10890 3782
rect 10582 3760 10890 3780
rect 10980 3618 11008 7398
rect 10888 3590 11008 3618
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9968 2514 9996 3470
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10796 2990 10824 3334
rect 10888 3058 10916 3590
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10980 3194 11008 3470
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 10428 2446 10456 2790
rect 10582 2748 10890 2768
rect 10582 2746 10588 2748
rect 10644 2746 10668 2748
rect 10724 2746 10748 2748
rect 10804 2746 10828 2748
rect 10884 2746 10890 2748
rect 10644 2694 10646 2746
rect 10826 2694 10828 2746
rect 10582 2692 10588 2694
rect 10644 2692 10668 2694
rect 10724 2692 10748 2694
rect 10804 2692 10828 2694
rect 10884 2692 10890 2694
rect 10582 2672 10890 2692
rect 11532 2446 11560 3334
rect 12360 3058 12388 7958
rect 13004 7954 13032 8230
rect 14292 8090 14320 8910
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 13360 8016 13412 8022
rect 13360 7958 13412 7964
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13372 3194 13400 7958
rect 15028 6458 15056 19110
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15120 7818 15148 8434
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 16408 6798 16436 19450
rect 17788 19378 17816 21200
rect 19168 19378 19196 21200
rect 20214 19612 20522 19632
rect 20214 19610 20220 19612
rect 20276 19610 20300 19612
rect 20356 19610 20380 19612
rect 20436 19610 20460 19612
rect 20516 19610 20522 19612
rect 20276 19558 20278 19610
rect 20458 19558 20460 19610
rect 20214 19556 20220 19558
rect 20276 19556 20300 19558
rect 20356 19556 20380 19558
rect 20436 19556 20460 19558
rect 20516 19556 20522 19558
rect 20214 19536 20522 19556
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17788 6866 17816 7210
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 16040 6390 16068 6598
rect 16028 6384 16080 6390
rect 16028 6326 16080 6332
rect 16592 6254 16620 6802
rect 17880 6798 17908 19110
rect 19260 7478 19288 19110
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19996 7342 20024 7686
rect 20088 7478 20116 19450
rect 20640 19378 20668 21200
rect 22020 19378 22048 21200
rect 22560 19508 22612 19514
rect 22560 19450 22612 19456
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 20214 18524 20522 18544
rect 20214 18522 20220 18524
rect 20276 18522 20300 18524
rect 20356 18522 20380 18524
rect 20436 18522 20460 18524
rect 20516 18522 20522 18524
rect 20276 18470 20278 18522
rect 20458 18470 20460 18522
rect 20214 18468 20220 18470
rect 20276 18468 20300 18470
rect 20356 18468 20380 18470
rect 20436 18468 20460 18470
rect 20516 18468 20522 18470
rect 20214 18448 20522 18468
rect 20214 17436 20522 17456
rect 20214 17434 20220 17436
rect 20276 17434 20300 17436
rect 20356 17434 20380 17436
rect 20436 17434 20460 17436
rect 20516 17434 20522 17436
rect 20276 17382 20278 17434
rect 20458 17382 20460 17434
rect 20214 17380 20220 17382
rect 20276 17380 20300 17382
rect 20356 17380 20380 17382
rect 20436 17380 20460 17382
rect 20516 17380 20522 17382
rect 20214 17360 20522 17380
rect 20214 16348 20522 16368
rect 20214 16346 20220 16348
rect 20276 16346 20300 16348
rect 20356 16346 20380 16348
rect 20436 16346 20460 16348
rect 20516 16346 20522 16348
rect 20276 16294 20278 16346
rect 20458 16294 20460 16346
rect 20214 16292 20220 16294
rect 20276 16292 20300 16294
rect 20356 16292 20380 16294
rect 20436 16292 20460 16294
rect 20516 16292 20522 16294
rect 20214 16272 20522 16292
rect 20214 15260 20522 15280
rect 20214 15258 20220 15260
rect 20276 15258 20300 15260
rect 20356 15258 20380 15260
rect 20436 15258 20460 15260
rect 20516 15258 20522 15260
rect 20276 15206 20278 15258
rect 20458 15206 20460 15258
rect 20214 15204 20220 15206
rect 20276 15204 20300 15206
rect 20356 15204 20380 15206
rect 20436 15204 20460 15206
rect 20516 15204 20522 15206
rect 20214 15184 20522 15204
rect 20214 14172 20522 14192
rect 20214 14170 20220 14172
rect 20276 14170 20300 14172
rect 20356 14170 20380 14172
rect 20436 14170 20460 14172
rect 20516 14170 20522 14172
rect 20276 14118 20278 14170
rect 20458 14118 20460 14170
rect 20214 14116 20220 14118
rect 20276 14116 20300 14118
rect 20356 14116 20380 14118
rect 20436 14116 20460 14118
rect 20516 14116 20522 14118
rect 20214 14096 20522 14116
rect 20214 13084 20522 13104
rect 20214 13082 20220 13084
rect 20276 13082 20300 13084
rect 20356 13082 20380 13084
rect 20436 13082 20460 13084
rect 20516 13082 20522 13084
rect 20276 13030 20278 13082
rect 20458 13030 20460 13082
rect 20214 13028 20220 13030
rect 20276 13028 20300 13030
rect 20356 13028 20380 13030
rect 20436 13028 20460 13030
rect 20516 13028 20522 13030
rect 20214 13008 20522 13028
rect 20214 11996 20522 12016
rect 20214 11994 20220 11996
rect 20276 11994 20300 11996
rect 20356 11994 20380 11996
rect 20436 11994 20460 11996
rect 20516 11994 20522 11996
rect 20276 11942 20278 11994
rect 20458 11942 20460 11994
rect 20214 11940 20220 11942
rect 20276 11940 20300 11942
rect 20356 11940 20380 11942
rect 20436 11940 20460 11942
rect 20516 11940 20522 11942
rect 20214 11920 20522 11940
rect 20214 10908 20522 10928
rect 20214 10906 20220 10908
rect 20276 10906 20300 10908
rect 20356 10906 20380 10908
rect 20436 10906 20460 10908
rect 20516 10906 20522 10908
rect 20276 10854 20278 10906
rect 20458 10854 20460 10906
rect 20214 10852 20220 10854
rect 20276 10852 20300 10854
rect 20356 10852 20380 10854
rect 20436 10852 20460 10854
rect 20516 10852 20522 10854
rect 20214 10832 20522 10852
rect 20214 9820 20522 9840
rect 20214 9818 20220 9820
rect 20276 9818 20300 9820
rect 20356 9818 20380 9820
rect 20436 9818 20460 9820
rect 20516 9818 20522 9820
rect 20276 9766 20278 9818
rect 20458 9766 20460 9818
rect 20214 9764 20220 9766
rect 20276 9764 20300 9766
rect 20356 9764 20380 9766
rect 20436 9764 20460 9766
rect 20516 9764 20522 9766
rect 20214 9744 20522 9764
rect 22572 8974 22600 19450
rect 23768 19378 23796 21270
rect 24858 21270 25176 21298
rect 24858 21200 24914 21270
rect 25148 19378 25176 21270
rect 26330 21200 26386 22000
rect 27710 21298 27766 22000
rect 27710 21270 28028 21298
rect 27710 21200 27766 21270
rect 26344 19378 26372 21200
rect 27344 19508 27396 19514
rect 27344 19450 27396 19456
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 25136 19372 25188 19378
rect 25136 19314 25188 19320
rect 26332 19372 26384 19378
rect 26332 19314 26384 19320
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 20214 8732 20522 8752
rect 20214 8730 20220 8732
rect 20276 8730 20300 8732
rect 20356 8730 20380 8732
rect 20436 8730 20460 8732
rect 20516 8730 20522 8732
rect 20276 8678 20278 8730
rect 20458 8678 20460 8730
rect 20214 8676 20220 8678
rect 20276 8676 20300 8678
rect 20356 8676 20380 8678
rect 20436 8676 20460 8678
rect 20516 8676 20522 8678
rect 20214 8656 20522 8676
rect 22480 8498 22508 8774
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 20996 8424 21048 8430
rect 20996 8366 21048 8372
rect 21008 8090 21036 8366
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 20214 7644 20522 7664
rect 20214 7642 20220 7644
rect 20276 7642 20300 7644
rect 20356 7642 20380 7644
rect 20436 7642 20460 7644
rect 20516 7642 20522 7644
rect 20276 7590 20278 7642
rect 20458 7590 20460 7642
rect 20214 7588 20220 7590
rect 20276 7588 20300 7590
rect 20356 7588 20380 7590
rect 20436 7588 20460 7590
rect 20516 7588 20522 7590
rect 20214 7568 20522 7588
rect 20076 7472 20128 7478
rect 20076 7414 20128 7420
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 13188 2446 13216 2790
rect 14108 2446 14136 2790
rect 15672 2582 15700 6190
rect 16684 2650 16712 6598
rect 17512 6322 17540 6598
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17880 2650 17908 6598
rect 19260 2650 19288 7278
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19628 6798 19656 7142
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 20214 6556 20522 6576
rect 20214 6554 20220 6556
rect 20276 6554 20300 6556
rect 20356 6554 20380 6556
rect 20436 6554 20460 6556
rect 20516 6554 20522 6556
rect 20276 6502 20278 6554
rect 20458 6502 20460 6554
rect 20214 6500 20220 6502
rect 20276 6500 20300 6502
rect 20356 6500 20380 6502
rect 20436 6500 20460 6502
rect 20516 6500 20522 6502
rect 20214 6480 20522 6500
rect 20214 5468 20522 5488
rect 20214 5466 20220 5468
rect 20276 5466 20300 5468
rect 20356 5466 20380 5468
rect 20436 5466 20460 5468
rect 20516 5466 20522 5468
rect 20276 5414 20278 5466
rect 20458 5414 20460 5466
rect 20214 5412 20220 5414
rect 20276 5412 20300 5414
rect 20356 5412 20380 5414
rect 20436 5412 20460 5414
rect 20516 5412 20522 5414
rect 20214 5392 20522 5412
rect 20214 4380 20522 4400
rect 20214 4378 20220 4380
rect 20276 4378 20300 4380
rect 20356 4378 20380 4380
rect 20436 4378 20460 4380
rect 20516 4378 20522 4380
rect 20276 4326 20278 4378
rect 20458 4326 20460 4378
rect 20214 4324 20220 4326
rect 20276 4324 20300 4326
rect 20356 4324 20380 4326
rect 20436 4324 20460 4326
rect 20516 4324 20522 4326
rect 20214 4304 20522 4324
rect 20214 3292 20522 3312
rect 20214 3290 20220 3292
rect 20276 3290 20300 3292
rect 20356 3290 20380 3292
rect 20436 3290 20460 3292
rect 20516 3290 20522 3292
rect 20276 3238 20278 3290
rect 20458 3238 20460 3290
rect 20214 3236 20220 3238
rect 20276 3236 20300 3238
rect 20356 3236 20380 3238
rect 20436 3236 20460 3238
rect 20516 3236 20522 3238
rect 20214 3216 20522 3236
rect 20732 2650 20760 7414
rect 20824 7274 20852 7822
rect 20812 7268 20864 7274
rect 20812 7210 20864 7216
rect 22664 2650 22692 8774
rect 23216 8634 23244 8910
rect 23584 8634 23612 19110
rect 24964 9654 24992 19110
rect 26516 11076 26568 11082
rect 26516 11018 26568 11024
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 26068 9654 26096 9862
rect 24952 9648 25004 9654
rect 24952 9590 25004 9596
rect 26056 9648 26108 9654
rect 26056 9590 26108 9596
rect 25044 9512 25096 9518
rect 25044 9454 25096 9460
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23768 9042 23796 9318
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23768 8430 23796 8978
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23676 2650 23704 8366
rect 25056 2650 25084 9454
rect 26528 8906 26556 11018
rect 26884 9988 26936 9994
rect 26884 9930 26936 9936
rect 26896 9722 26924 9930
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 27356 9654 27384 19450
rect 28000 19378 28028 21270
rect 29182 21200 29238 22000
rect 30654 21298 30710 22000
rect 32034 21298 32090 22000
rect 33506 21298 33562 22000
rect 34886 21298 34942 22000
rect 36358 21298 36414 22000
rect 37738 21298 37794 22000
rect 30654 21270 30972 21298
rect 30654 21200 30710 21270
rect 29196 19378 29224 21200
rect 29644 19508 29696 19514
rect 29644 19450 29696 19456
rect 27988 19372 28040 19378
rect 27988 19314 28040 19320
rect 29184 19372 29236 19378
rect 29184 19314 29236 19320
rect 27804 19168 27856 19174
rect 27804 19110 27856 19116
rect 27344 9648 27396 9654
rect 27344 9590 27396 9596
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 27356 9042 27384 9386
rect 27344 9036 27396 9042
rect 27344 8978 27396 8984
rect 26516 8900 26568 8906
rect 26516 8842 26568 8848
rect 26528 7818 26556 8842
rect 26516 7812 26568 7818
rect 26516 7754 26568 7760
rect 27448 2650 27476 9454
rect 27816 8974 27844 19110
rect 29656 11898 29684 19450
rect 30944 19378 30972 21270
rect 32034 21270 32352 21298
rect 32034 21200 32090 21270
rect 31024 19508 31076 19514
rect 31024 19450 31076 19456
rect 30932 19372 30984 19378
rect 30932 19314 30984 19320
rect 29846 19068 30154 19088
rect 29846 19066 29852 19068
rect 29908 19066 29932 19068
rect 29988 19066 30012 19068
rect 30068 19066 30092 19068
rect 30148 19066 30154 19068
rect 29908 19014 29910 19066
rect 30090 19014 30092 19066
rect 29846 19012 29852 19014
rect 29908 19012 29932 19014
rect 29988 19012 30012 19014
rect 30068 19012 30092 19014
rect 30148 19012 30154 19014
rect 29846 18992 30154 19012
rect 29846 17980 30154 18000
rect 29846 17978 29852 17980
rect 29908 17978 29932 17980
rect 29988 17978 30012 17980
rect 30068 17978 30092 17980
rect 30148 17978 30154 17980
rect 29908 17926 29910 17978
rect 30090 17926 30092 17978
rect 29846 17924 29852 17926
rect 29908 17924 29932 17926
rect 29988 17924 30012 17926
rect 30068 17924 30092 17926
rect 30148 17924 30154 17926
rect 29846 17904 30154 17924
rect 29846 16892 30154 16912
rect 29846 16890 29852 16892
rect 29908 16890 29932 16892
rect 29988 16890 30012 16892
rect 30068 16890 30092 16892
rect 30148 16890 30154 16892
rect 29908 16838 29910 16890
rect 30090 16838 30092 16890
rect 29846 16836 29852 16838
rect 29908 16836 29932 16838
rect 29988 16836 30012 16838
rect 30068 16836 30092 16838
rect 30148 16836 30154 16838
rect 29846 16816 30154 16836
rect 29846 15804 30154 15824
rect 29846 15802 29852 15804
rect 29908 15802 29932 15804
rect 29988 15802 30012 15804
rect 30068 15802 30092 15804
rect 30148 15802 30154 15804
rect 29908 15750 29910 15802
rect 30090 15750 30092 15802
rect 29846 15748 29852 15750
rect 29908 15748 29932 15750
rect 29988 15748 30012 15750
rect 30068 15748 30092 15750
rect 30148 15748 30154 15750
rect 29846 15728 30154 15748
rect 29846 14716 30154 14736
rect 29846 14714 29852 14716
rect 29908 14714 29932 14716
rect 29988 14714 30012 14716
rect 30068 14714 30092 14716
rect 30148 14714 30154 14716
rect 29908 14662 29910 14714
rect 30090 14662 30092 14714
rect 29846 14660 29852 14662
rect 29908 14660 29932 14662
rect 29988 14660 30012 14662
rect 30068 14660 30092 14662
rect 30148 14660 30154 14662
rect 29846 14640 30154 14660
rect 29846 13628 30154 13648
rect 29846 13626 29852 13628
rect 29908 13626 29932 13628
rect 29988 13626 30012 13628
rect 30068 13626 30092 13628
rect 30148 13626 30154 13628
rect 29908 13574 29910 13626
rect 30090 13574 30092 13626
rect 29846 13572 29852 13574
rect 29908 13572 29932 13574
rect 29988 13572 30012 13574
rect 30068 13572 30092 13574
rect 30148 13572 30154 13574
rect 29846 13552 30154 13572
rect 29846 12540 30154 12560
rect 29846 12538 29852 12540
rect 29908 12538 29932 12540
rect 29988 12538 30012 12540
rect 30068 12538 30092 12540
rect 30148 12538 30154 12540
rect 29908 12486 29910 12538
rect 30090 12486 30092 12538
rect 29846 12484 29852 12486
rect 29908 12484 29932 12486
rect 29988 12484 30012 12486
rect 30068 12484 30092 12486
rect 30148 12484 30154 12486
rect 29846 12464 30154 12484
rect 30656 12164 30708 12170
rect 30656 12106 30708 12112
rect 30668 11898 30696 12106
rect 31036 11898 31064 19450
rect 32324 19378 32352 21270
rect 33506 21270 33824 21298
rect 33506 21200 33562 21270
rect 32496 19508 32548 19514
rect 32496 19450 32548 19456
rect 33692 19508 33744 19514
rect 33692 19450 33744 19456
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32128 12164 32180 12170
rect 32128 12106 32180 12112
rect 32140 11898 32168 12106
rect 32508 11898 32536 19450
rect 32772 12300 32824 12306
rect 32772 12242 32824 12248
rect 29644 11892 29696 11898
rect 29644 11834 29696 11840
rect 30656 11892 30708 11898
rect 30656 11834 30708 11840
rect 31024 11892 31076 11898
rect 31024 11834 31076 11840
rect 32128 11892 32180 11898
rect 32128 11834 32180 11840
rect 32496 11892 32548 11898
rect 32496 11834 32548 11840
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 29552 11688 29604 11694
rect 29552 11630 29604 11636
rect 30748 11688 30800 11694
rect 30748 11630 30800 11636
rect 27988 9988 28040 9994
rect 27988 9930 28040 9936
rect 28000 9178 28028 9930
rect 27988 9172 28040 9178
rect 27988 9114 28040 9120
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27632 2650 27660 8774
rect 29564 2650 29592 11630
rect 30196 11552 30248 11558
rect 30196 11494 30248 11500
rect 29846 11452 30154 11472
rect 29846 11450 29852 11452
rect 29908 11450 29932 11452
rect 29988 11450 30012 11452
rect 30068 11450 30092 11452
rect 30148 11450 30154 11452
rect 29908 11398 29910 11450
rect 30090 11398 30092 11450
rect 29846 11396 29852 11398
rect 29908 11396 29932 11398
rect 29988 11396 30012 11398
rect 30068 11396 30092 11398
rect 30148 11396 30154 11398
rect 29846 11376 30154 11396
rect 30208 11150 30236 11494
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 29846 10364 30154 10384
rect 29846 10362 29852 10364
rect 29908 10362 29932 10364
rect 29988 10362 30012 10364
rect 30068 10362 30092 10364
rect 30148 10362 30154 10364
rect 29908 10310 29910 10362
rect 30090 10310 30092 10362
rect 29846 10308 29852 10310
rect 29908 10308 29932 10310
rect 29988 10308 30012 10310
rect 30068 10308 30092 10310
rect 30148 10308 30154 10310
rect 29846 10288 30154 10308
rect 29846 9276 30154 9296
rect 29846 9274 29852 9276
rect 29908 9274 29932 9276
rect 29988 9274 30012 9276
rect 30068 9274 30092 9276
rect 30148 9274 30154 9276
rect 29908 9222 29910 9274
rect 30090 9222 30092 9274
rect 29846 9220 29852 9222
rect 29908 9220 29932 9222
rect 29988 9220 30012 9222
rect 30068 9220 30092 9222
rect 30148 9220 30154 9222
rect 29846 9200 30154 9220
rect 29846 8188 30154 8208
rect 29846 8186 29852 8188
rect 29908 8186 29932 8188
rect 29988 8186 30012 8188
rect 30068 8186 30092 8188
rect 30148 8186 30154 8188
rect 29908 8134 29910 8186
rect 30090 8134 30092 8186
rect 29846 8132 29852 8134
rect 29908 8132 29932 8134
rect 29988 8132 30012 8134
rect 30068 8132 30092 8134
rect 30148 8132 30154 8134
rect 29846 8112 30154 8132
rect 29846 7100 30154 7120
rect 29846 7098 29852 7100
rect 29908 7098 29932 7100
rect 29988 7098 30012 7100
rect 30068 7098 30092 7100
rect 30148 7098 30154 7100
rect 29908 7046 29910 7098
rect 30090 7046 30092 7098
rect 29846 7044 29852 7046
rect 29908 7044 29932 7046
rect 29988 7044 30012 7046
rect 30068 7044 30092 7046
rect 30148 7044 30154 7046
rect 29846 7024 30154 7044
rect 29846 6012 30154 6032
rect 29846 6010 29852 6012
rect 29908 6010 29932 6012
rect 29988 6010 30012 6012
rect 30068 6010 30092 6012
rect 30148 6010 30154 6012
rect 29908 5958 29910 6010
rect 30090 5958 30092 6010
rect 29846 5956 29852 5958
rect 29908 5956 29932 5958
rect 29988 5956 30012 5958
rect 30068 5956 30092 5958
rect 30148 5956 30154 5958
rect 29846 5936 30154 5956
rect 29846 4924 30154 4944
rect 29846 4922 29852 4924
rect 29908 4922 29932 4924
rect 29988 4922 30012 4924
rect 30068 4922 30092 4924
rect 30148 4922 30154 4924
rect 29908 4870 29910 4922
rect 30090 4870 30092 4922
rect 29846 4868 29852 4870
rect 29908 4868 29932 4870
rect 29988 4868 30012 4870
rect 30068 4868 30092 4870
rect 30148 4868 30154 4870
rect 29846 4848 30154 4868
rect 29846 3836 30154 3856
rect 29846 3834 29852 3836
rect 29908 3834 29932 3836
rect 29988 3834 30012 3836
rect 30068 3834 30092 3836
rect 30148 3834 30154 3836
rect 29908 3782 29910 3834
rect 30090 3782 30092 3834
rect 29846 3780 29852 3782
rect 29908 3780 29932 3782
rect 29988 3780 30012 3782
rect 30068 3780 30092 3782
rect 30148 3780 30154 3782
rect 29846 3760 30154 3780
rect 29846 2748 30154 2768
rect 29846 2746 29852 2748
rect 29908 2746 29932 2748
rect 29988 2746 30012 2748
rect 30068 2746 30092 2748
rect 30148 2746 30154 2748
rect 29908 2694 29910 2746
rect 30090 2694 30092 2746
rect 29846 2692 29852 2694
rect 29908 2692 29932 2694
rect 29988 2692 30012 2694
rect 30068 2692 30092 2694
rect 30148 2692 30154 2694
rect 29846 2672 30154 2692
rect 30760 2650 30788 11630
rect 31036 11354 31064 11698
rect 32784 11694 32812 12242
rect 33704 12238 33732 19450
rect 33796 19378 33824 21270
rect 34886 21270 35204 21298
rect 34886 21200 34942 21270
rect 35072 19508 35124 19514
rect 35072 19450 35124 19456
rect 33784 19372 33836 19378
rect 33784 19314 33836 19320
rect 34244 12776 34296 12782
rect 34244 12718 34296 12724
rect 33692 12232 33744 12238
rect 33692 12174 33744 12180
rect 33324 12096 33376 12102
rect 33324 12038 33376 12044
rect 33600 12096 33652 12102
rect 33600 12038 33652 12044
rect 33336 11830 33364 12038
rect 33324 11824 33376 11830
rect 33324 11766 33376 11772
rect 32128 11688 32180 11694
rect 32128 11630 32180 11636
rect 32772 11688 32824 11694
rect 32772 11630 32824 11636
rect 31024 11348 31076 11354
rect 31024 11290 31076 11296
rect 32140 2650 32168 11630
rect 33612 2650 33640 12038
rect 34256 11830 34284 12718
rect 35084 12238 35112 19450
rect 35176 19378 35204 21270
rect 36358 21270 36676 21298
rect 36358 21200 36414 21270
rect 36648 19378 36676 21270
rect 37738 21270 38056 21298
rect 37738 21200 37794 21270
rect 38028 19378 38056 21270
rect 39210 21200 39266 22000
rect 40590 21298 40646 22000
rect 40590 21270 40908 21298
rect 40590 21200 40646 21270
rect 39224 19378 39252 21200
rect 39478 19612 39786 19632
rect 39478 19610 39484 19612
rect 39540 19610 39564 19612
rect 39620 19610 39644 19612
rect 39700 19610 39724 19612
rect 39780 19610 39786 19612
rect 39540 19558 39542 19610
rect 39722 19558 39724 19610
rect 39478 19556 39484 19558
rect 39540 19556 39564 19558
rect 39620 19556 39644 19558
rect 39700 19556 39724 19558
rect 39780 19556 39786 19558
rect 39478 19536 39786 19556
rect 39304 19508 39356 19514
rect 39304 19450 39356 19456
rect 35164 19372 35216 19378
rect 35164 19314 35216 19320
rect 36636 19372 36688 19378
rect 36636 19314 36688 19320
rect 38016 19372 38068 19378
rect 38016 19314 38068 19320
rect 39212 19372 39264 19378
rect 39212 19314 39264 19320
rect 36452 19168 36504 19174
rect 36452 19110 36504 19116
rect 37832 19168 37884 19174
rect 37832 19110 37884 19116
rect 36464 13326 36492 19110
rect 37844 14414 37872 19110
rect 39316 15162 39344 19450
rect 40880 19378 40908 21270
rect 42062 21200 42118 22000
rect 43442 21298 43498 22000
rect 43442 21270 43760 21298
rect 43442 21200 43498 21270
rect 41512 19508 41564 19514
rect 41512 19450 41564 19456
rect 41880 19508 41932 19514
rect 41880 19450 41932 19456
rect 40868 19372 40920 19378
rect 40868 19314 40920 19320
rect 39478 18524 39786 18544
rect 39478 18522 39484 18524
rect 39540 18522 39564 18524
rect 39620 18522 39644 18524
rect 39700 18522 39724 18524
rect 39780 18522 39786 18524
rect 39540 18470 39542 18522
rect 39722 18470 39724 18522
rect 39478 18468 39484 18470
rect 39540 18468 39564 18470
rect 39620 18468 39644 18470
rect 39700 18468 39724 18470
rect 39780 18468 39786 18470
rect 39478 18448 39786 18468
rect 39478 17436 39786 17456
rect 39478 17434 39484 17436
rect 39540 17434 39564 17436
rect 39620 17434 39644 17436
rect 39700 17434 39724 17436
rect 39780 17434 39786 17436
rect 39540 17382 39542 17434
rect 39722 17382 39724 17434
rect 39478 17380 39484 17382
rect 39540 17380 39564 17382
rect 39620 17380 39644 17382
rect 39700 17380 39724 17382
rect 39780 17380 39786 17382
rect 39478 17360 39786 17380
rect 39478 16348 39786 16368
rect 39478 16346 39484 16348
rect 39540 16346 39564 16348
rect 39620 16346 39644 16348
rect 39700 16346 39724 16348
rect 39780 16346 39786 16348
rect 39540 16294 39542 16346
rect 39722 16294 39724 16346
rect 39478 16292 39484 16294
rect 39540 16292 39564 16294
rect 39620 16292 39644 16294
rect 39700 16292 39724 16294
rect 39780 16292 39786 16294
rect 39478 16272 39786 16292
rect 39478 15260 39786 15280
rect 39478 15258 39484 15260
rect 39540 15258 39564 15260
rect 39620 15258 39644 15260
rect 39700 15258 39724 15260
rect 39780 15258 39786 15260
rect 39540 15206 39542 15258
rect 39722 15206 39724 15258
rect 39478 15204 39484 15206
rect 39540 15204 39564 15206
rect 39620 15204 39644 15206
rect 39700 15204 39724 15206
rect 39780 15204 39786 15206
rect 39478 15184 39786 15204
rect 39304 15156 39356 15162
rect 39304 15098 39356 15104
rect 39764 15020 39816 15026
rect 39764 14962 39816 14968
rect 38108 14884 38160 14890
rect 38108 14826 38160 14832
rect 38120 14482 38148 14826
rect 38108 14476 38160 14482
rect 38108 14418 38160 14424
rect 37832 14408 37884 14414
rect 37832 14350 37884 14356
rect 37464 14272 37516 14278
rect 37464 14214 37516 14220
rect 37740 14272 37792 14278
rect 37740 14214 37792 14220
rect 37476 13938 37504 14214
rect 37464 13932 37516 13938
rect 37464 13874 37516 13880
rect 36452 13320 36504 13326
rect 36452 13262 36504 13268
rect 36360 13184 36412 13190
rect 36360 13126 36412 13132
rect 35164 12844 35216 12850
rect 35164 12786 35216 12792
rect 35176 12442 35204 12786
rect 35164 12436 35216 12442
rect 35164 12378 35216 12384
rect 35072 12232 35124 12238
rect 35072 12174 35124 12180
rect 34980 12096 35032 12102
rect 34980 12038 35032 12044
rect 34244 11824 34296 11830
rect 34244 11766 34296 11772
rect 34992 2650 35020 12038
rect 36372 2650 36400 13126
rect 37752 2650 37780 14214
rect 38120 13258 38148 14418
rect 39776 14362 39804 14962
rect 41144 14952 41196 14958
rect 41144 14894 41196 14900
rect 39856 14816 39908 14822
rect 39856 14758 39908 14764
rect 39868 14482 39896 14758
rect 41156 14618 41184 14894
rect 41144 14612 41196 14618
rect 41144 14554 41196 14560
rect 39856 14476 39908 14482
rect 39856 14418 39908 14424
rect 39776 14334 39896 14362
rect 41524 14346 41552 19450
rect 41892 15502 41920 19450
rect 42076 19378 42104 21200
rect 43732 19378 43760 21270
rect 44914 21200 44970 22000
rect 46294 21298 46350 22000
rect 47766 21298 47822 22000
rect 49146 21298 49202 22000
rect 50618 21298 50674 22000
rect 51998 21298 52054 22000
rect 53470 21298 53526 22000
rect 54850 21298 54906 22000
rect 55954 21720 56010 21729
rect 55954 21655 56010 21664
rect 46294 21270 46612 21298
rect 46294 21200 46350 21270
rect 43996 19508 44048 19514
rect 43996 19450 44048 19456
rect 42064 19372 42116 19378
rect 42064 19314 42116 19320
rect 43720 19372 43772 19378
rect 43720 19314 43772 19320
rect 42984 17196 43036 17202
rect 42984 17138 43036 17144
rect 42064 15564 42116 15570
rect 42064 15506 42116 15512
rect 41880 15496 41932 15502
rect 41880 15438 41932 15444
rect 41880 15360 41932 15366
rect 41880 15302 41932 15308
rect 41892 14958 41920 15302
rect 41880 14952 41932 14958
rect 41880 14894 41932 14900
rect 42076 14890 42104 15506
rect 42340 15360 42392 15366
rect 42340 15302 42392 15308
rect 42064 14884 42116 14890
rect 42064 14826 42116 14832
rect 42076 14482 42104 14826
rect 42064 14476 42116 14482
rect 42064 14418 42116 14424
rect 39478 14172 39786 14192
rect 39478 14170 39484 14172
rect 39540 14170 39564 14172
rect 39620 14170 39644 14172
rect 39700 14170 39724 14172
rect 39780 14170 39786 14172
rect 39540 14118 39542 14170
rect 39722 14118 39724 14170
rect 39478 14116 39484 14118
rect 39540 14116 39564 14118
rect 39620 14116 39644 14118
rect 39700 14116 39724 14118
rect 39780 14116 39786 14118
rect 39478 14096 39786 14116
rect 38108 13252 38160 13258
rect 38108 13194 38160 13200
rect 38120 12986 38148 13194
rect 39478 13084 39786 13104
rect 39478 13082 39484 13084
rect 39540 13082 39564 13084
rect 39620 13082 39644 13084
rect 39700 13082 39724 13084
rect 39780 13082 39786 13084
rect 39540 13030 39542 13082
rect 39722 13030 39724 13082
rect 39478 13028 39484 13030
rect 39540 13028 39564 13030
rect 39620 13028 39644 13030
rect 39700 13028 39724 13030
rect 39780 13028 39786 13030
rect 39478 13008 39786 13028
rect 38108 12980 38160 12986
rect 38108 12922 38160 12928
rect 38384 12844 38436 12850
rect 38384 12786 38436 12792
rect 38396 12102 38424 12786
rect 38660 12232 38712 12238
rect 38660 12174 38712 12180
rect 38384 12096 38436 12102
rect 38384 12038 38436 12044
rect 38396 11082 38424 12038
rect 38672 11286 38700 12174
rect 39478 11996 39786 12016
rect 39478 11994 39484 11996
rect 39540 11994 39564 11996
rect 39620 11994 39644 11996
rect 39700 11994 39724 11996
rect 39780 11994 39786 11996
rect 39540 11942 39542 11994
rect 39722 11942 39724 11994
rect 39478 11940 39484 11942
rect 39540 11940 39564 11942
rect 39620 11940 39644 11942
rect 39700 11940 39724 11942
rect 39780 11940 39786 11942
rect 39478 11920 39786 11940
rect 38660 11280 38712 11286
rect 38660 11222 38712 11228
rect 38384 11076 38436 11082
rect 38384 11018 38436 11024
rect 39478 10908 39786 10928
rect 39478 10906 39484 10908
rect 39540 10906 39564 10908
rect 39620 10906 39644 10908
rect 39700 10906 39724 10908
rect 39780 10906 39786 10908
rect 39540 10854 39542 10906
rect 39722 10854 39724 10906
rect 39478 10852 39484 10854
rect 39540 10852 39564 10854
rect 39620 10852 39644 10854
rect 39700 10852 39724 10854
rect 39780 10852 39786 10854
rect 39478 10832 39786 10852
rect 39478 9820 39786 9840
rect 39478 9818 39484 9820
rect 39540 9818 39564 9820
rect 39620 9818 39644 9820
rect 39700 9818 39724 9820
rect 39780 9818 39786 9820
rect 39540 9766 39542 9818
rect 39722 9766 39724 9818
rect 39478 9764 39484 9766
rect 39540 9764 39564 9766
rect 39620 9764 39644 9766
rect 39700 9764 39724 9766
rect 39780 9764 39786 9766
rect 39478 9744 39786 9764
rect 39478 8732 39786 8752
rect 39478 8730 39484 8732
rect 39540 8730 39564 8732
rect 39620 8730 39644 8732
rect 39700 8730 39724 8732
rect 39780 8730 39786 8732
rect 39540 8678 39542 8730
rect 39722 8678 39724 8730
rect 39478 8676 39484 8678
rect 39540 8676 39564 8678
rect 39620 8676 39644 8678
rect 39700 8676 39724 8678
rect 39780 8676 39786 8678
rect 39478 8656 39786 8676
rect 39478 7644 39786 7664
rect 39478 7642 39484 7644
rect 39540 7642 39564 7644
rect 39620 7642 39644 7644
rect 39700 7642 39724 7644
rect 39780 7642 39786 7644
rect 39540 7590 39542 7642
rect 39722 7590 39724 7642
rect 39478 7588 39484 7590
rect 39540 7588 39564 7590
rect 39620 7588 39644 7590
rect 39700 7588 39724 7590
rect 39780 7588 39786 7590
rect 39478 7568 39786 7588
rect 39478 6556 39786 6576
rect 39478 6554 39484 6556
rect 39540 6554 39564 6556
rect 39620 6554 39644 6556
rect 39700 6554 39724 6556
rect 39780 6554 39786 6556
rect 39540 6502 39542 6554
rect 39722 6502 39724 6554
rect 39478 6500 39484 6502
rect 39540 6500 39564 6502
rect 39620 6500 39644 6502
rect 39700 6500 39724 6502
rect 39780 6500 39786 6502
rect 39478 6480 39786 6500
rect 39478 5468 39786 5488
rect 39478 5466 39484 5468
rect 39540 5466 39564 5468
rect 39620 5466 39644 5468
rect 39700 5466 39724 5468
rect 39780 5466 39786 5468
rect 39540 5414 39542 5466
rect 39722 5414 39724 5466
rect 39478 5412 39484 5414
rect 39540 5412 39564 5414
rect 39620 5412 39644 5414
rect 39700 5412 39724 5414
rect 39780 5412 39786 5414
rect 39478 5392 39786 5412
rect 39478 4380 39786 4400
rect 39478 4378 39484 4380
rect 39540 4378 39564 4380
rect 39620 4378 39644 4380
rect 39700 4378 39724 4380
rect 39780 4378 39786 4380
rect 39540 4326 39542 4378
rect 39722 4326 39724 4378
rect 39478 4324 39484 4326
rect 39540 4324 39564 4326
rect 39620 4324 39644 4326
rect 39700 4324 39724 4326
rect 39780 4324 39786 4326
rect 39478 4304 39786 4324
rect 39478 3292 39786 3312
rect 39478 3290 39484 3292
rect 39540 3290 39564 3292
rect 39620 3290 39644 3292
rect 39700 3290 39724 3292
rect 39780 3290 39786 3292
rect 39540 3238 39542 3290
rect 39722 3238 39724 3290
rect 39478 3236 39484 3238
rect 39540 3236 39564 3238
rect 39620 3236 39644 3238
rect 39700 3236 39724 3238
rect 39780 3236 39786 3238
rect 39478 3216 39786 3236
rect 39868 2650 39896 14334
rect 41512 14340 41564 14346
rect 41512 14282 41564 14288
rect 41604 14272 41656 14278
rect 41604 14214 41656 14220
rect 40224 11212 40276 11218
rect 40224 11154 40276 11160
rect 40236 11082 40264 11154
rect 40224 11076 40276 11082
rect 40224 11018 40276 11024
rect 40236 6914 40264 11018
rect 40144 6886 40264 6914
rect 40144 3534 40172 6886
rect 40132 3528 40184 3534
rect 40132 3470 40184 3476
rect 41616 2650 41644 14214
rect 42352 2650 42380 15302
rect 42996 11286 43024 17138
rect 43536 16652 43588 16658
rect 43536 16594 43588 16600
rect 42984 11280 43036 11286
rect 42984 11222 43036 11228
rect 43548 2650 43576 16594
rect 44008 16590 44036 19450
rect 44928 19378 44956 21200
rect 45376 19508 45428 19514
rect 45376 19450 45428 19456
rect 44916 19372 44968 19378
rect 44916 19314 44968 19320
rect 45008 16992 45060 16998
rect 45008 16934 45060 16940
rect 45020 16794 45048 16934
rect 45008 16788 45060 16794
rect 45008 16730 45060 16736
rect 45008 16652 45060 16658
rect 45008 16594 45060 16600
rect 43996 16584 44048 16590
rect 43996 16526 44048 16532
rect 43628 16448 43680 16454
rect 43628 16390 43680 16396
rect 43640 16114 43668 16390
rect 43628 16108 43680 16114
rect 43628 16050 43680 16056
rect 45020 2650 45048 16594
rect 45388 16590 45416 19450
rect 46584 19378 46612 21270
rect 47766 21270 48084 21298
rect 47766 21200 47822 21270
rect 48056 19378 48084 21270
rect 49146 21270 49464 21298
rect 49146 21200 49202 21270
rect 48964 19508 49016 19514
rect 48964 19450 49016 19456
rect 46572 19372 46624 19378
rect 46572 19314 46624 19320
rect 48044 19372 48096 19378
rect 48044 19314 48096 19320
rect 46388 19168 46440 19174
rect 46388 19110 46440 19116
rect 47860 19168 47912 19174
rect 47860 19110 47912 19116
rect 46020 17672 46072 17678
rect 46020 17614 46072 17620
rect 46032 17338 46060 17614
rect 46400 17338 46428 19110
rect 47584 17672 47636 17678
rect 47584 17614 47636 17620
rect 46756 17536 46808 17542
rect 46756 17478 46808 17484
rect 46020 17332 46072 17338
rect 46020 17274 46072 17280
rect 46388 17332 46440 17338
rect 46388 17274 46440 17280
rect 46768 17270 46796 17478
rect 47596 17338 47624 17614
rect 47872 17338 47900 19110
rect 48228 17740 48280 17746
rect 48228 17682 48280 17688
rect 47584 17332 47636 17338
rect 47584 17274 47636 17280
rect 47860 17332 47912 17338
rect 47860 17274 47912 17280
rect 46756 17264 46808 17270
rect 46756 17206 46808 17212
rect 48240 17134 48268 17682
rect 48976 17678 49004 19450
rect 49436 19378 49464 21270
rect 50618 21270 50936 21298
rect 50618 21200 50674 21270
rect 50908 19378 50936 21270
rect 51998 21270 52224 21298
rect 51998 21200 52054 21270
rect 51172 19508 51224 19514
rect 51172 19450 51224 19456
rect 49424 19372 49476 19378
rect 49424 19314 49476 19320
rect 50896 19372 50948 19378
rect 50896 19314 50948 19320
rect 49110 19068 49418 19088
rect 49110 19066 49116 19068
rect 49172 19066 49196 19068
rect 49252 19066 49276 19068
rect 49332 19066 49356 19068
rect 49412 19066 49418 19068
rect 49172 19014 49174 19066
rect 49354 19014 49356 19066
rect 49110 19012 49116 19014
rect 49172 19012 49196 19014
rect 49252 19012 49276 19014
rect 49332 19012 49356 19014
rect 49412 19012 49418 19014
rect 49110 18992 49418 19012
rect 51080 18896 51132 18902
rect 51080 18838 51132 18844
rect 50804 18624 50856 18630
rect 50804 18566 50856 18572
rect 50988 18624 51040 18630
rect 50988 18566 51040 18572
rect 50816 18290 50844 18566
rect 50804 18284 50856 18290
rect 50804 18226 50856 18232
rect 49110 17980 49418 18000
rect 49110 17978 49116 17980
rect 49172 17978 49196 17980
rect 49252 17978 49276 17980
rect 49332 17978 49356 17980
rect 49412 17978 49418 17980
rect 49172 17926 49174 17978
rect 49354 17926 49356 17978
rect 49110 17924 49116 17926
rect 49172 17924 49196 17926
rect 49252 17924 49276 17926
rect 49332 17924 49356 17926
rect 49412 17924 49418 17926
rect 49110 17904 49418 17924
rect 48964 17672 49016 17678
rect 48964 17614 49016 17620
rect 49516 17536 49568 17542
rect 49516 17478 49568 17484
rect 46296 17128 46348 17134
rect 46296 17070 46348 17076
rect 48044 17128 48096 17134
rect 48044 17070 48096 17076
rect 48228 17128 48280 17134
rect 48228 17070 48280 17076
rect 45376 16584 45428 16590
rect 45376 16526 45428 16532
rect 46308 2650 46336 17070
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 25044 2644 25096 2650
rect 25044 2586 25096 2592
rect 27436 2644 27488 2650
rect 27436 2586 27488 2592
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 30748 2644 30800 2650
rect 30748 2586 30800 2592
rect 32128 2644 32180 2650
rect 32128 2586 32180 2592
rect 33600 2644 33652 2650
rect 33600 2586 33652 2592
rect 34980 2644 35032 2650
rect 34980 2586 35032 2592
rect 36360 2644 36412 2650
rect 36360 2586 36412 2592
rect 37740 2644 37792 2650
rect 37740 2586 37792 2592
rect 39856 2644 39908 2650
rect 39856 2586 39908 2592
rect 41604 2644 41656 2650
rect 41604 2586 41656 2592
rect 42340 2644 42392 2650
rect 42340 2586 42392 2592
rect 43536 2644 43588 2650
rect 43536 2586 43588 2592
rect 45008 2644 45060 2650
rect 45008 2586 45060 2592
rect 46296 2644 46348 2650
rect 46296 2586 46348 2592
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 48056 2514 48084 17070
rect 48240 16998 48268 17070
rect 48228 16992 48280 16998
rect 48228 16934 48280 16940
rect 49110 16892 49418 16912
rect 49110 16890 49116 16892
rect 49172 16890 49196 16892
rect 49252 16890 49276 16892
rect 49332 16890 49356 16892
rect 49412 16890 49418 16892
rect 49172 16838 49174 16890
rect 49354 16838 49356 16890
rect 49110 16836 49116 16838
rect 49172 16836 49196 16838
rect 49252 16836 49276 16838
rect 49332 16836 49356 16838
rect 49412 16836 49418 16838
rect 49110 16816 49418 16836
rect 49110 15804 49418 15824
rect 49110 15802 49116 15804
rect 49172 15802 49196 15804
rect 49252 15802 49276 15804
rect 49332 15802 49356 15804
rect 49412 15802 49418 15804
rect 49172 15750 49174 15802
rect 49354 15750 49356 15802
rect 49110 15748 49116 15750
rect 49172 15748 49196 15750
rect 49252 15748 49276 15750
rect 49332 15748 49356 15750
rect 49412 15748 49418 15750
rect 49110 15728 49418 15748
rect 49110 14716 49418 14736
rect 49110 14714 49116 14716
rect 49172 14714 49196 14716
rect 49252 14714 49276 14716
rect 49332 14714 49356 14716
rect 49412 14714 49418 14716
rect 49172 14662 49174 14714
rect 49354 14662 49356 14714
rect 49110 14660 49116 14662
rect 49172 14660 49196 14662
rect 49252 14660 49276 14662
rect 49332 14660 49356 14662
rect 49412 14660 49418 14662
rect 49110 14640 49418 14660
rect 49110 13628 49418 13648
rect 49110 13626 49116 13628
rect 49172 13626 49196 13628
rect 49252 13626 49276 13628
rect 49332 13626 49356 13628
rect 49412 13626 49418 13628
rect 49172 13574 49174 13626
rect 49354 13574 49356 13626
rect 49110 13572 49116 13574
rect 49172 13572 49196 13574
rect 49252 13572 49276 13574
rect 49332 13572 49356 13574
rect 49412 13572 49418 13574
rect 49110 13552 49418 13572
rect 49110 12540 49418 12560
rect 49110 12538 49116 12540
rect 49172 12538 49196 12540
rect 49252 12538 49276 12540
rect 49332 12538 49356 12540
rect 49412 12538 49418 12540
rect 49172 12486 49174 12538
rect 49354 12486 49356 12538
rect 49110 12484 49116 12486
rect 49172 12484 49196 12486
rect 49252 12484 49276 12486
rect 49332 12484 49356 12486
rect 49412 12484 49418 12486
rect 49110 12464 49418 12484
rect 49110 11452 49418 11472
rect 49110 11450 49116 11452
rect 49172 11450 49196 11452
rect 49252 11450 49276 11452
rect 49332 11450 49356 11452
rect 49412 11450 49418 11452
rect 49172 11398 49174 11450
rect 49354 11398 49356 11450
rect 49110 11396 49116 11398
rect 49172 11396 49196 11398
rect 49252 11396 49276 11398
rect 49332 11396 49356 11398
rect 49412 11396 49418 11398
rect 49110 11376 49418 11396
rect 49110 10364 49418 10384
rect 49110 10362 49116 10364
rect 49172 10362 49196 10364
rect 49252 10362 49276 10364
rect 49332 10362 49356 10364
rect 49412 10362 49418 10364
rect 49172 10310 49174 10362
rect 49354 10310 49356 10362
rect 49110 10308 49116 10310
rect 49172 10308 49196 10310
rect 49252 10308 49276 10310
rect 49332 10308 49356 10310
rect 49412 10308 49418 10310
rect 49110 10288 49418 10308
rect 49110 9276 49418 9296
rect 49110 9274 49116 9276
rect 49172 9274 49196 9276
rect 49252 9274 49276 9276
rect 49332 9274 49356 9276
rect 49412 9274 49418 9276
rect 49172 9222 49174 9274
rect 49354 9222 49356 9274
rect 49110 9220 49116 9222
rect 49172 9220 49196 9222
rect 49252 9220 49276 9222
rect 49332 9220 49356 9222
rect 49412 9220 49418 9222
rect 49110 9200 49418 9220
rect 49110 8188 49418 8208
rect 49110 8186 49116 8188
rect 49172 8186 49196 8188
rect 49252 8186 49276 8188
rect 49332 8186 49356 8188
rect 49412 8186 49418 8188
rect 49172 8134 49174 8186
rect 49354 8134 49356 8186
rect 49110 8132 49116 8134
rect 49172 8132 49196 8134
rect 49252 8132 49276 8134
rect 49332 8132 49356 8134
rect 49412 8132 49418 8134
rect 49110 8112 49418 8132
rect 49110 7100 49418 7120
rect 49110 7098 49116 7100
rect 49172 7098 49196 7100
rect 49252 7098 49276 7100
rect 49332 7098 49356 7100
rect 49412 7098 49418 7100
rect 49172 7046 49174 7098
rect 49354 7046 49356 7098
rect 49110 7044 49116 7046
rect 49172 7044 49196 7046
rect 49252 7044 49276 7046
rect 49332 7044 49356 7046
rect 49412 7044 49418 7046
rect 49110 7024 49418 7044
rect 49110 6012 49418 6032
rect 49110 6010 49116 6012
rect 49172 6010 49196 6012
rect 49252 6010 49276 6012
rect 49332 6010 49356 6012
rect 49412 6010 49418 6012
rect 49172 5958 49174 6010
rect 49354 5958 49356 6010
rect 49110 5956 49116 5958
rect 49172 5956 49196 5958
rect 49252 5956 49276 5958
rect 49332 5956 49356 5958
rect 49412 5956 49418 5958
rect 49110 5936 49418 5956
rect 49110 4924 49418 4944
rect 49110 4922 49116 4924
rect 49172 4922 49196 4924
rect 49252 4922 49276 4924
rect 49332 4922 49356 4924
rect 49412 4922 49418 4924
rect 49172 4870 49174 4922
rect 49354 4870 49356 4922
rect 49110 4868 49116 4870
rect 49172 4868 49196 4870
rect 49252 4868 49276 4870
rect 49332 4868 49356 4870
rect 49412 4868 49418 4870
rect 49110 4848 49418 4868
rect 49110 3836 49418 3856
rect 49110 3834 49116 3836
rect 49172 3834 49196 3836
rect 49252 3834 49276 3836
rect 49332 3834 49356 3836
rect 49412 3834 49418 3836
rect 49172 3782 49174 3834
rect 49354 3782 49356 3834
rect 49110 3780 49116 3782
rect 49172 3780 49196 3782
rect 49252 3780 49276 3782
rect 49332 3780 49356 3782
rect 49412 3780 49418 3782
rect 49110 3760 49418 3780
rect 48412 3392 48464 3398
rect 48412 3334 48464 3340
rect 48424 3194 48452 3334
rect 48412 3188 48464 3194
rect 48412 3130 48464 3136
rect 49528 3058 49556 17478
rect 50252 15020 50304 15026
rect 50252 14962 50304 14968
rect 50264 14414 50292 14962
rect 50252 14408 50304 14414
rect 50252 14350 50304 14356
rect 50344 14408 50396 14414
rect 50344 14350 50396 14356
rect 50356 13870 50384 14350
rect 50344 13864 50396 13870
rect 50344 13806 50396 13812
rect 50344 12300 50396 12306
rect 50344 12242 50396 12248
rect 50356 11762 50384 12242
rect 50344 11756 50396 11762
rect 50344 11698 50396 11704
rect 50344 9580 50396 9586
rect 50344 9522 50396 9528
rect 50356 8974 50384 9522
rect 50344 8968 50396 8974
rect 50344 8910 50396 8916
rect 50436 8968 50488 8974
rect 50436 8910 50488 8916
rect 50448 8566 50476 8910
rect 50436 8560 50488 8566
rect 50436 8502 50488 8508
rect 50344 6792 50396 6798
rect 50344 6734 50396 6740
rect 50356 6118 50384 6734
rect 50344 6112 50396 6118
rect 50344 6054 50396 6060
rect 49516 3052 49568 3058
rect 49516 2994 49568 3000
rect 48964 2984 49016 2990
rect 48964 2926 49016 2932
rect 48044 2508 48096 2514
rect 48044 2450 48096 2456
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 24860 2440 24912 2446
rect 24860 2382 24912 2388
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 29184 2440 29236 2446
rect 29184 2382 29236 2388
rect 30656 2440 30708 2446
rect 30656 2382 30708 2388
rect 32036 2440 32088 2446
rect 32036 2382 32088 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 34888 2440 34940 2446
rect 34888 2382 34940 2388
rect 36360 2440 36412 2446
rect 36360 2382 36412 2388
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 39212 2440 39264 2446
rect 39212 2382 39264 2388
rect 40592 2440 40644 2446
rect 40592 2382 40644 2388
rect 42064 2440 42116 2446
rect 42064 2382 42116 2388
rect 43444 2440 43496 2446
rect 43444 2382 43496 2388
rect 44916 2440 44968 2446
rect 44916 2382 44968 2388
rect 46296 2440 46348 2446
rect 46296 2382 46348 2388
rect 47768 2440 47820 2446
rect 47768 2382 47820 2388
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 10704 1170 10732 2246
rect 10612 1142 10732 1170
rect 10612 800 10640 1142
rect 12084 800 12112 2246
rect 13464 800 13492 2246
rect 14936 800 14964 2382
rect 16316 800 16344 2382
rect 17788 800 17816 2382
rect 19168 800 19196 2382
rect 20214 2204 20522 2224
rect 20214 2202 20220 2204
rect 20276 2202 20300 2204
rect 20356 2202 20380 2204
rect 20436 2202 20460 2204
rect 20516 2202 20522 2204
rect 20276 2150 20278 2202
rect 20458 2150 20460 2202
rect 20214 2148 20220 2150
rect 20276 2148 20300 2150
rect 20356 2148 20380 2150
rect 20436 2148 20460 2150
rect 20516 2148 20522 2150
rect 20214 2128 20522 2148
rect 20640 800 20668 2382
rect 22020 800 22048 2382
rect 23492 800 23520 2382
rect 24872 800 24900 2382
rect 26344 800 26372 2382
rect 27724 800 27752 2382
rect 29196 800 29224 2382
rect 30668 800 30696 2382
rect 32048 800 32076 2382
rect 33520 800 33548 2382
rect 34900 800 34928 2382
rect 36372 800 36400 2382
rect 37752 800 37780 2382
rect 39224 800 39252 2382
rect 39478 2204 39786 2224
rect 39478 2202 39484 2204
rect 39540 2202 39564 2204
rect 39620 2202 39644 2204
rect 39700 2202 39724 2204
rect 39780 2202 39786 2204
rect 39540 2150 39542 2202
rect 39722 2150 39724 2202
rect 39478 2148 39484 2150
rect 39540 2148 39564 2150
rect 39620 2148 39644 2150
rect 39700 2148 39724 2150
rect 39780 2148 39786 2150
rect 39478 2128 39786 2148
rect 40604 800 40632 2382
rect 42076 800 42104 2382
rect 43456 800 43484 2382
rect 44928 800 44956 2382
rect 46308 800 46336 2382
rect 47780 800 47808 2382
rect 48976 1578 49004 2926
rect 49110 2748 49418 2768
rect 49110 2746 49116 2748
rect 49172 2746 49196 2748
rect 49252 2746 49276 2748
rect 49332 2746 49356 2748
rect 49412 2746 49418 2748
rect 49172 2694 49174 2746
rect 49354 2694 49356 2746
rect 49110 2692 49116 2694
rect 49172 2692 49196 2694
rect 49252 2692 49276 2694
rect 49332 2692 49356 2694
rect 49412 2692 49418 2694
rect 49110 2672 49418 2692
rect 51000 2514 51028 18566
rect 51092 17542 51120 18838
rect 51184 18766 51212 19450
rect 52196 19378 52224 21270
rect 53470 21270 53788 21298
rect 53470 21200 53526 21270
rect 53012 19848 53064 19854
rect 53012 19790 53064 19796
rect 52184 19372 52236 19378
rect 52184 19314 52236 19320
rect 52276 19168 52328 19174
rect 52276 19110 52328 19116
rect 51172 18760 51224 18766
rect 51172 18702 51224 18708
rect 52288 18630 52316 19110
rect 52368 18760 52420 18766
rect 52368 18702 52420 18708
rect 52000 18624 52052 18630
rect 52000 18566 52052 18572
rect 52276 18624 52328 18630
rect 52276 18566 52328 18572
rect 52012 18290 52040 18566
rect 52000 18284 52052 18290
rect 52000 18226 52052 18232
rect 51080 17536 51132 17542
rect 51080 17478 51132 17484
rect 52380 2514 52408 18702
rect 53024 18426 53052 19790
rect 53380 19780 53432 19786
rect 53380 19722 53432 19728
rect 53392 19378 53420 19722
rect 53380 19372 53432 19378
rect 53380 19314 53432 19320
rect 53564 18624 53616 18630
rect 53564 18566 53616 18572
rect 53576 18426 53604 18566
rect 53012 18420 53064 18426
rect 53012 18362 53064 18368
rect 53564 18420 53616 18426
rect 53564 18362 53616 18368
rect 53760 18290 53788 21270
rect 54772 21270 54906 21298
rect 53932 19712 53984 19718
rect 53932 19654 53984 19660
rect 53840 18624 53892 18630
rect 53840 18566 53892 18572
rect 53748 18284 53800 18290
rect 53748 18226 53800 18232
rect 52460 13932 52512 13938
rect 52460 13874 52512 13880
rect 52472 13326 52500 13874
rect 52460 13320 52512 13326
rect 52460 13262 52512 13268
rect 52552 13320 52604 13326
rect 52552 13262 52604 13268
rect 52564 12714 52592 13262
rect 52552 12708 52604 12714
rect 52552 12650 52604 12656
rect 53852 3058 53880 18566
rect 53944 18154 53972 19654
rect 54024 19372 54076 19378
rect 54024 19314 54076 19320
rect 54036 18970 54064 19314
rect 54024 18964 54076 18970
rect 54024 18906 54076 18912
rect 54772 18290 54800 21270
rect 54850 21200 54906 21270
rect 55770 20088 55826 20097
rect 55770 20023 55826 20032
rect 55784 19378 55812 20023
rect 55588 19372 55640 19378
rect 55588 19314 55640 19320
rect 55772 19372 55824 19378
rect 55772 19314 55824 19320
rect 55600 18970 55628 19314
rect 55588 18964 55640 18970
rect 55588 18906 55640 18912
rect 55864 18828 55916 18834
rect 55864 18770 55916 18776
rect 55496 18692 55548 18698
rect 55496 18634 55548 18640
rect 54760 18284 54812 18290
rect 54760 18226 54812 18232
rect 53932 18148 53984 18154
rect 53932 18090 53984 18096
rect 53840 3052 53892 3058
rect 53840 2994 53892 3000
rect 53472 2984 53524 2990
rect 53472 2926 53524 2932
rect 50988 2508 51040 2514
rect 50988 2450 51040 2456
rect 52368 2508 52420 2514
rect 52368 2450 52420 2456
rect 50620 2440 50672 2446
rect 50620 2382 50672 2388
rect 52000 2440 52052 2446
rect 52000 2382 52052 2388
rect 48976 1550 49188 1578
rect 49160 800 49188 1550
rect 50632 800 50660 2382
rect 52012 800 52040 2382
rect 53484 800 53512 2926
rect 55508 2514 55536 18634
rect 55680 18624 55732 18630
rect 55680 18566 55732 18572
rect 55692 18426 55720 18566
rect 55680 18420 55732 18426
rect 55680 18362 55732 18368
rect 55876 17882 55904 18770
rect 55968 17882 55996 21655
rect 56322 21200 56378 22000
rect 57702 21298 57758 22000
rect 57348 21270 57758 21298
rect 56230 21176 56286 21185
rect 56230 21111 56286 21120
rect 56046 20632 56102 20641
rect 56046 20567 56102 20576
rect 56060 18426 56088 20567
rect 56244 19514 56272 21111
rect 56232 19508 56284 19514
rect 56232 19450 56284 19456
rect 56048 18420 56100 18426
rect 56048 18362 56100 18368
rect 55864 17876 55916 17882
rect 55864 17818 55916 17824
rect 55956 17876 56008 17882
rect 55956 17818 56008 17824
rect 55772 17604 55824 17610
rect 55772 17546 55824 17552
rect 55784 17066 55812 17546
rect 56336 17202 56364 21200
rect 57152 19848 57204 19854
rect 57152 19790 57204 19796
rect 56968 19780 57020 19786
rect 56968 19722 57020 19728
rect 56506 19680 56562 19689
rect 56506 19615 56562 19624
rect 56520 19514 56548 19615
rect 56508 19508 56560 19514
rect 56508 19450 56560 19456
rect 56692 18692 56744 18698
rect 56692 18634 56744 18640
rect 56508 18624 56560 18630
rect 56508 18566 56560 18572
rect 56520 18358 56548 18566
rect 56508 18352 56560 18358
rect 56508 18294 56560 18300
rect 56600 18284 56652 18290
rect 56600 18226 56652 18232
rect 56324 17196 56376 17202
rect 56324 17138 56376 17144
rect 55772 17060 55824 17066
rect 55772 17002 55824 17008
rect 55784 5914 55812 17002
rect 56612 16454 56640 18226
rect 56600 16448 56652 16454
rect 56600 16390 56652 16396
rect 56600 15496 56652 15502
rect 56600 15438 56652 15444
rect 56612 14958 56640 15438
rect 56600 14952 56652 14958
rect 56600 14894 56652 14900
rect 55772 5908 55824 5914
rect 55772 5850 55824 5856
rect 56508 5228 56560 5234
rect 56508 5170 56560 5176
rect 56520 4729 56548 5170
rect 56506 4720 56562 4729
rect 56506 4655 56562 4664
rect 56508 4548 56560 4554
rect 56508 4490 56560 4496
rect 56520 4321 56548 4490
rect 56600 4480 56652 4486
rect 56600 4422 56652 4428
rect 56506 4312 56562 4321
rect 56506 4247 56562 4256
rect 56048 4208 56100 4214
rect 56048 4150 56100 4156
rect 55680 3936 55732 3942
rect 55680 3878 55732 3884
rect 55692 3194 55720 3878
rect 55772 3460 55824 3466
rect 55772 3402 55824 3408
rect 55680 3188 55732 3194
rect 55680 3130 55732 3136
rect 55588 3052 55640 3058
rect 55588 2994 55640 3000
rect 55496 2508 55548 2514
rect 55496 2450 55548 2456
rect 54852 2440 54904 2446
rect 54852 2382 54904 2388
rect 54864 800 54892 2382
rect 55128 2372 55180 2378
rect 55128 2314 55180 2320
rect 5000 734 5212 762
rect 6366 0 6422 800
rect 7746 0 7802 800
rect 9218 0 9274 800
rect 10598 0 10654 800
rect 12070 0 12126 800
rect 13450 0 13506 800
rect 14922 0 14978 800
rect 16302 0 16358 800
rect 17774 0 17830 800
rect 19154 0 19210 800
rect 20626 0 20682 800
rect 22006 0 22062 800
rect 23478 0 23534 800
rect 24858 0 24914 800
rect 26330 0 26386 800
rect 27710 0 27766 800
rect 29182 0 29238 800
rect 30654 0 30710 800
rect 32034 0 32090 800
rect 33506 0 33562 800
rect 34886 0 34942 800
rect 36358 0 36414 800
rect 37738 0 37794 800
rect 39210 0 39266 800
rect 40590 0 40646 800
rect 42062 0 42118 800
rect 43442 0 43498 800
rect 44914 0 44970 800
rect 46294 0 46350 800
rect 47766 0 47822 800
rect 49146 0 49202 800
rect 50618 0 50674 800
rect 51998 0 52054 800
rect 53470 0 53526 800
rect 54850 0 54906 800
rect 55140 82 55168 2314
rect 55600 2281 55628 2994
rect 55784 2689 55812 3402
rect 56060 3233 56088 4150
rect 56508 3460 56560 3466
rect 56508 3402 56560 3408
rect 56046 3224 56102 3233
rect 56046 3159 56102 3168
rect 56324 2984 56376 2990
rect 56324 2926 56376 2932
rect 55770 2680 55826 2689
rect 55770 2615 55826 2624
rect 55586 2272 55642 2281
rect 55586 2207 55642 2216
rect 56336 800 56364 2926
rect 56520 1193 56548 3402
rect 56612 3126 56640 4422
rect 56600 3120 56652 3126
rect 56600 3062 56652 3068
rect 56704 3058 56732 18634
rect 56876 18624 56928 18630
rect 56876 18566 56928 18572
rect 56784 18216 56836 18222
rect 56784 18158 56836 18164
rect 56796 17814 56824 18158
rect 56784 17808 56836 17814
rect 56784 17750 56836 17756
rect 56796 11218 56824 17750
rect 56888 17066 56916 18566
rect 56980 17882 57008 19722
rect 57060 19712 57112 19718
rect 57060 19654 57112 19660
rect 57072 19378 57100 19654
rect 57164 19378 57192 19790
rect 57060 19372 57112 19378
rect 57060 19314 57112 19320
rect 57152 19372 57204 19378
rect 57152 19314 57204 19320
rect 57244 19168 57296 19174
rect 57242 19136 57244 19145
rect 57296 19136 57298 19145
rect 57242 19071 57298 19080
rect 57244 18284 57296 18290
rect 57244 18226 57296 18232
rect 56968 17876 57020 17882
rect 56968 17818 57020 17824
rect 57256 17746 57284 18226
rect 57244 17740 57296 17746
rect 57244 17682 57296 17688
rect 57152 17672 57204 17678
rect 57152 17614 57204 17620
rect 56968 17604 57020 17610
rect 56968 17546 57020 17552
rect 56876 17060 56928 17066
rect 56876 17002 56928 17008
rect 56784 11212 56836 11218
rect 56784 11154 56836 11160
rect 56876 5636 56928 5642
rect 56876 5578 56928 5584
rect 56888 5273 56916 5578
rect 56874 5264 56930 5273
rect 56874 5199 56930 5208
rect 56784 5024 56836 5030
rect 56784 4966 56836 4972
rect 56796 3398 56824 4966
rect 56980 3534 57008 17546
rect 57164 16794 57192 17614
rect 57242 17096 57298 17105
rect 57242 17031 57244 17040
rect 57296 17031 57298 17040
rect 57244 17002 57296 17008
rect 57152 16788 57204 16794
rect 57152 16730 57204 16736
rect 57060 16720 57112 16726
rect 57060 16662 57112 16668
rect 57072 16590 57100 16662
rect 57060 16584 57112 16590
rect 57060 16526 57112 16532
rect 57348 16114 57376 21270
rect 57702 21200 57758 21270
rect 59174 21200 59230 22000
rect 57888 19508 57940 19514
rect 57888 19450 57940 19456
rect 57900 18601 57928 19450
rect 58072 18624 58124 18630
rect 57886 18592 57942 18601
rect 58072 18566 58124 18572
rect 57886 18527 57942 18536
rect 57704 18352 57756 18358
rect 57704 18294 57756 18300
rect 57428 18080 57480 18086
rect 57428 18022 57480 18028
rect 57440 16590 57468 18022
rect 57520 17536 57572 17542
rect 57520 17478 57572 17484
rect 57428 16584 57480 16590
rect 57428 16526 57480 16532
rect 57532 16250 57560 17478
rect 57612 17196 57664 17202
rect 57612 17138 57664 17144
rect 57624 16522 57652 17138
rect 57612 16516 57664 16522
rect 57612 16458 57664 16464
rect 57520 16244 57572 16250
rect 57520 16186 57572 16192
rect 57336 16108 57388 16114
rect 57336 16050 57388 16056
rect 57428 16108 57480 16114
rect 57428 16050 57480 16056
rect 57440 15094 57468 16050
rect 57428 15088 57480 15094
rect 57428 15030 57480 15036
rect 57060 10668 57112 10674
rect 57060 10610 57112 10616
rect 57152 10668 57204 10674
rect 57152 10610 57204 10616
rect 57072 10062 57100 10610
rect 57060 10056 57112 10062
rect 57060 9998 57112 10004
rect 57164 9994 57192 10610
rect 57244 10464 57296 10470
rect 57242 10432 57244 10441
rect 57296 10432 57298 10441
rect 57242 10367 57298 10376
rect 57152 9988 57204 9994
rect 57152 9930 57204 9936
rect 57520 7744 57572 7750
rect 57520 7686 57572 7692
rect 57428 7404 57480 7410
rect 57428 7346 57480 7352
rect 57440 7206 57468 7346
rect 57428 7200 57480 7206
rect 57428 7142 57480 7148
rect 57440 6254 57468 7142
rect 57532 6662 57560 7686
rect 57716 6914 57744 18294
rect 57888 18080 57940 18086
rect 58084 18057 58112 18566
rect 57888 18022 57940 18028
rect 58070 18048 58126 18057
rect 57900 17649 57928 18022
rect 58070 17983 58126 17992
rect 57886 17640 57942 17649
rect 57886 17575 57942 17584
rect 58072 16992 58124 16998
rect 58072 16934 58124 16940
rect 57888 16584 57940 16590
rect 58084 16561 58112 16934
rect 59188 16726 59216 21200
rect 59176 16720 59228 16726
rect 59176 16662 59228 16668
rect 57888 16526 57940 16532
rect 58070 16552 58126 16561
rect 57900 15910 57928 16526
rect 58070 16487 58126 16496
rect 58072 16448 58124 16454
rect 58072 16390 58124 16396
rect 58084 16017 58112 16390
rect 58070 16008 58126 16017
rect 58070 15943 58126 15952
rect 57888 15904 57940 15910
rect 57888 15846 57940 15852
rect 58072 15904 58124 15910
rect 58072 15846 58124 15852
rect 58084 15609 58112 15846
rect 58070 15600 58126 15609
rect 58070 15535 58126 15544
rect 57888 15360 57940 15366
rect 57888 15302 57940 15308
rect 57900 15065 57928 15302
rect 57886 15056 57942 15065
rect 57886 14991 57942 15000
rect 58072 14816 58124 14822
rect 58072 14758 58124 14764
rect 58084 14521 58112 14758
rect 58070 14512 58126 14521
rect 58070 14447 58126 14456
rect 58072 14272 58124 14278
rect 58072 14214 58124 14220
rect 57888 14068 57940 14074
rect 57888 14010 57940 14016
rect 57900 13433 57928 14010
rect 58084 13977 58112 14214
rect 58070 13968 58126 13977
rect 58070 13903 58126 13912
rect 57886 13424 57942 13433
rect 57886 13359 57942 13368
rect 58072 13184 58124 13190
rect 58072 13126 58124 13132
rect 58084 13025 58112 13126
rect 58070 13016 58126 13025
rect 58070 12951 58126 12960
rect 58072 12640 58124 12646
rect 58072 12582 58124 12588
rect 58084 12481 58112 12582
rect 58070 12472 58126 12481
rect 58070 12407 58126 12416
rect 58072 12096 58124 12102
rect 58072 12038 58124 12044
rect 58084 11937 58112 12038
rect 58070 11928 58126 11937
rect 58070 11863 58126 11872
rect 58072 11552 58124 11558
rect 58072 11494 58124 11500
rect 58084 11393 58112 11494
rect 58070 11384 58126 11393
rect 58070 11319 58126 11328
rect 57888 11280 57940 11286
rect 57888 11222 57940 11228
rect 57900 10985 57928 11222
rect 57886 10976 57942 10985
rect 57886 10911 57942 10920
rect 58072 10464 58124 10470
rect 58072 10406 58124 10412
rect 57888 9920 57940 9926
rect 58084 9897 58112 10406
rect 57888 9862 57940 9868
rect 58070 9888 58126 9897
rect 57900 9353 57928 9862
rect 58070 9823 58126 9832
rect 58072 9376 58124 9382
rect 57886 9344 57942 9353
rect 58072 9318 58124 9324
rect 57886 9279 57942 9288
rect 58084 8945 58112 9318
rect 58070 8936 58126 8945
rect 58070 8871 58126 8880
rect 58072 8832 58124 8838
rect 58072 8774 58124 8780
rect 58084 8401 58112 8774
rect 58070 8392 58126 8401
rect 57888 8356 57940 8362
rect 58070 8327 58126 8336
rect 57888 8298 57940 8304
rect 57900 7857 57928 8298
rect 57886 7848 57942 7857
rect 57886 7783 57942 7792
rect 58072 7744 58124 7750
rect 58072 7686 58124 7692
rect 57980 7540 58032 7546
rect 57980 7482 58032 7488
rect 57624 6886 57744 6914
rect 57520 6656 57572 6662
rect 57520 6598 57572 6604
rect 57428 6248 57480 6254
rect 57428 6190 57480 6196
rect 57624 4690 57652 6886
rect 57992 5846 58020 7482
rect 58084 7313 58112 7686
rect 58070 7304 58126 7313
rect 58070 7239 58126 7248
rect 58072 7200 58124 7206
rect 58072 7142 58124 7148
rect 58084 6769 58112 7142
rect 58070 6760 58126 6769
rect 58070 6695 58126 6704
rect 58072 6656 58124 6662
rect 58072 6598 58124 6604
rect 58084 6361 58112 6598
rect 58070 6352 58126 6361
rect 58070 6287 58126 6296
rect 58072 6112 58124 6118
rect 58072 6054 58124 6060
rect 57980 5840 58032 5846
rect 58084 5817 58112 6054
rect 57980 5782 58032 5788
rect 58070 5808 58126 5817
rect 58070 5743 58126 5752
rect 57796 5636 57848 5642
rect 57796 5578 57848 5584
rect 57612 4684 57664 4690
rect 57612 4626 57664 4632
rect 57152 4208 57204 4214
rect 57152 4150 57204 4156
rect 57060 3936 57112 3942
rect 57060 3878 57112 3884
rect 57072 3602 57100 3878
rect 57060 3596 57112 3602
rect 57060 3538 57112 3544
rect 56968 3528 57020 3534
rect 56968 3470 57020 3476
rect 56784 3392 56836 3398
rect 56784 3334 56836 3340
rect 56692 3052 56744 3058
rect 56692 2994 56744 3000
rect 56968 2372 57020 2378
rect 56968 2314 57020 2320
rect 56506 1184 56562 1193
rect 56506 1119 56562 1128
rect 55218 232 55274 241
rect 55218 167 55274 176
rect 55232 82 55260 167
rect 55140 54 55260 82
rect 56322 0 56378 800
rect 56980 649 57008 2314
rect 57164 1737 57192 4150
rect 57808 3777 57836 5578
rect 59176 4616 59228 4622
rect 59176 4558 59228 4564
rect 57794 3768 57850 3777
rect 57794 3703 57850 3712
rect 57704 3596 57756 3602
rect 57704 3538 57756 3544
rect 57150 1728 57206 1737
rect 57150 1663 57206 1672
rect 57716 800 57744 3538
rect 59188 800 59216 4558
rect 56966 640 57022 649
rect 56966 575 57022 584
rect 57702 0 57758 800
rect 59174 0 59230 800
<< via2 >>
rect 10588 19066 10644 19068
rect 10668 19066 10724 19068
rect 10748 19066 10804 19068
rect 10828 19066 10884 19068
rect 10588 19014 10634 19066
rect 10634 19014 10644 19066
rect 10668 19014 10698 19066
rect 10698 19014 10710 19066
rect 10710 19014 10724 19066
rect 10748 19014 10762 19066
rect 10762 19014 10774 19066
rect 10774 19014 10804 19066
rect 10828 19014 10838 19066
rect 10838 19014 10884 19066
rect 10588 19012 10644 19014
rect 10668 19012 10724 19014
rect 10748 19012 10804 19014
rect 10828 19012 10884 19014
rect 10588 17978 10644 17980
rect 10668 17978 10724 17980
rect 10748 17978 10804 17980
rect 10828 17978 10884 17980
rect 10588 17926 10634 17978
rect 10634 17926 10644 17978
rect 10668 17926 10698 17978
rect 10698 17926 10710 17978
rect 10710 17926 10724 17978
rect 10748 17926 10762 17978
rect 10762 17926 10774 17978
rect 10774 17926 10804 17978
rect 10828 17926 10838 17978
rect 10838 17926 10884 17978
rect 10588 17924 10644 17926
rect 10668 17924 10724 17926
rect 10748 17924 10804 17926
rect 10828 17924 10884 17926
rect 10588 16890 10644 16892
rect 10668 16890 10724 16892
rect 10748 16890 10804 16892
rect 10828 16890 10884 16892
rect 10588 16838 10634 16890
rect 10634 16838 10644 16890
rect 10668 16838 10698 16890
rect 10698 16838 10710 16890
rect 10710 16838 10724 16890
rect 10748 16838 10762 16890
rect 10762 16838 10774 16890
rect 10774 16838 10804 16890
rect 10828 16838 10838 16890
rect 10838 16838 10884 16890
rect 10588 16836 10644 16838
rect 10668 16836 10724 16838
rect 10748 16836 10804 16838
rect 10828 16836 10884 16838
rect 10588 15802 10644 15804
rect 10668 15802 10724 15804
rect 10748 15802 10804 15804
rect 10828 15802 10884 15804
rect 10588 15750 10634 15802
rect 10634 15750 10644 15802
rect 10668 15750 10698 15802
rect 10698 15750 10710 15802
rect 10710 15750 10724 15802
rect 10748 15750 10762 15802
rect 10762 15750 10774 15802
rect 10774 15750 10804 15802
rect 10828 15750 10838 15802
rect 10838 15750 10884 15802
rect 10588 15748 10644 15750
rect 10668 15748 10724 15750
rect 10748 15748 10804 15750
rect 10828 15748 10884 15750
rect 10588 14714 10644 14716
rect 10668 14714 10724 14716
rect 10748 14714 10804 14716
rect 10828 14714 10884 14716
rect 10588 14662 10634 14714
rect 10634 14662 10644 14714
rect 10668 14662 10698 14714
rect 10698 14662 10710 14714
rect 10710 14662 10724 14714
rect 10748 14662 10762 14714
rect 10762 14662 10774 14714
rect 10774 14662 10804 14714
rect 10828 14662 10838 14714
rect 10838 14662 10884 14714
rect 10588 14660 10644 14662
rect 10668 14660 10724 14662
rect 10748 14660 10804 14662
rect 10828 14660 10884 14662
rect 10588 13626 10644 13628
rect 10668 13626 10724 13628
rect 10748 13626 10804 13628
rect 10828 13626 10884 13628
rect 10588 13574 10634 13626
rect 10634 13574 10644 13626
rect 10668 13574 10698 13626
rect 10698 13574 10710 13626
rect 10710 13574 10724 13626
rect 10748 13574 10762 13626
rect 10762 13574 10774 13626
rect 10774 13574 10804 13626
rect 10828 13574 10838 13626
rect 10838 13574 10884 13626
rect 10588 13572 10644 13574
rect 10668 13572 10724 13574
rect 10748 13572 10804 13574
rect 10828 13572 10884 13574
rect 10588 12538 10644 12540
rect 10668 12538 10724 12540
rect 10748 12538 10804 12540
rect 10828 12538 10884 12540
rect 10588 12486 10634 12538
rect 10634 12486 10644 12538
rect 10668 12486 10698 12538
rect 10698 12486 10710 12538
rect 10710 12486 10724 12538
rect 10748 12486 10762 12538
rect 10762 12486 10774 12538
rect 10774 12486 10804 12538
rect 10828 12486 10838 12538
rect 10838 12486 10884 12538
rect 10588 12484 10644 12486
rect 10668 12484 10724 12486
rect 10748 12484 10804 12486
rect 10828 12484 10884 12486
rect 10588 11450 10644 11452
rect 10668 11450 10724 11452
rect 10748 11450 10804 11452
rect 10828 11450 10884 11452
rect 10588 11398 10634 11450
rect 10634 11398 10644 11450
rect 10668 11398 10698 11450
rect 10698 11398 10710 11450
rect 10710 11398 10724 11450
rect 10748 11398 10762 11450
rect 10762 11398 10774 11450
rect 10774 11398 10804 11450
rect 10828 11398 10838 11450
rect 10838 11398 10884 11450
rect 10588 11396 10644 11398
rect 10668 11396 10724 11398
rect 10748 11396 10804 11398
rect 10828 11396 10884 11398
rect 10588 10362 10644 10364
rect 10668 10362 10724 10364
rect 10748 10362 10804 10364
rect 10828 10362 10884 10364
rect 10588 10310 10634 10362
rect 10634 10310 10644 10362
rect 10668 10310 10698 10362
rect 10698 10310 10710 10362
rect 10710 10310 10724 10362
rect 10748 10310 10762 10362
rect 10762 10310 10774 10362
rect 10774 10310 10804 10362
rect 10828 10310 10838 10362
rect 10838 10310 10884 10362
rect 10588 10308 10644 10310
rect 10668 10308 10724 10310
rect 10748 10308 10804 10310
rect 10828 10308 10884 10310
rect 10588 9274 10644 9276
rect 10668 9274 10724 9276
rect 10748 9274 10804 9276
rect 10828 9274 10884 9276
rect 10588 9222 10634 9274
rect 10634 9222 10644 9274
rect 10668 9222 10698 9274
rect 10698 9222 10710 9274
rect 10710 9222 10724 9274
rect 10748 9222 10762 9274
rect 10762 9222 10774 9274
rect 10774 9222 10804 9274
rect 10828 9222 10838 9274
rect 10838 9222 10884 9274
rect 10588 9220 10644 9222
rect 10668 9220 10724 9222
rect 10748 9220 10804 9222
rect 10828 9220 10884 9222
rect 10588 8186 10644 8188
rect 10668 8186 10724 8188
rect 10748 8186 10804 8188
rect 10828 8186 10884 8188
rect 10588 8134 10634 8186
rect 10634 8134 10644 8186
rect 10668 8134 10698 8186
rect 10698 8134 10710 8186
rect 10710 8134 10724 8186
rect 10748 8134 10762 8186
rect 10762 8134 10774 8186
rect 10774 8134 10804 8186
rect 10828 8134 10838 8186
rect 10838 8134 10884 8186
rect 10588 8132 10644 8134
rect 10668 8132 10724 8134
rect 10748 8132 10804 8134
rect 10828 8132 10884 8134
rect 10588 7098 10644 7100
rect 10668 7098 10724 7100
rect 10748 7098 10804 7100
rect 10828 7098 10884 7100
rect 10588 7046 10634 7098
rect 10634 7046 10644 7098
rect 10668 7046 10698 7098
rect 10698 7046 10710 7098
rect 10710 7046 10724 7098
rect 10748 7046 10762 7098
rect 10762 7046 10774 7098
rect 10774 7046 10804 7098
rect 10828 7046 10838 7098
rect 10838 7046 10884 7098
rect 10588 7044 10644 7046
rect 10668 7044 10724 7046
rect 10748 7044 10804 7046
rect 10828 7044 10884 7046
rect 10588 6010 10644 6012
rect 10668 6010 10724 6012
rect 10748 6010 10804 6012
rect 10828 6010 10884 6012
rect 10588 5958 10634 6010
rect 10634 5958 10644 6010
rect 10668 5958 10698 6010
rect 10698 5958 10710 6010
rect 10710 5958 10724 6010
rect 10748 5958 10762 6010
rect 10762 5958 10774 6010
rect 10774 5958 10804 6010
rect 10828 5958 10838 6010
rect 10838 5958 10884 6010
rect 10588 5956 10644 5958
rect 10668 5956 10724 5958
rect 10748 5956 10804 5958
rect 10828 5956 10884 5958
rect 10588 4922 10644 4924
rect 10668 4922 10724 4924
rect 10748 4922 10804 4924
rect 10828 4922 10884 4924
rect 10588 4870 10634 4922
rect 10634 4870 10644 4922
rect 10668 4870 10698 4922
rect 10698 4870 10710 4922
rect 10710 4870 10724 4922
rect 10748 4870 10762 4922
rect 10762 4870 10774 4922
rect 10774 4870 10804 4922
rect 10828 4870 10838 4922
rect 10838 4870 10884 4922
rect 10588 4868 10644 4870
rect 10668 4868 10724 4870
rect 10748 4868 10804 4870
rect 10828 4868 10884 4870
rect 10588 3834 10644 3836
rect 10668 3834 10724 3836
rect 10748 3834 10804 3836
rect 10828 3834 10884 3836
rect 10588 3782 10634 3834
rect 10634 3782 10644 3834
rect 10668 3782 10698 3834
rect 10698 3782 10710 3834
rect 10710 3782 10724 3834
rect 10748 3782 10762 3834
rect 10762 3782 10774 3834
rect 10774 3782 10804 3834
rect 10828 3782 10838 3834
rect 10838 3782 10884 3834
rect 10588 3780 10644 3782
rect 10668 3780 10724 3782
rect 10748 3780 10804 3782
rect 10828 3780 10884 3782
rect 10588 2746 10644 2748
rect 10668 2746 10724 2748
rect 10748 2746 10804 2748
rect 10828 2746 10884 2748
rect 10588 2694 10634 2746
rect 10634 2694 10644 2746
rect 10668 2694 10698 2746
rect 10698 2694 10710 2746
rect 10710 2694 10724 2746
rect 10748 2694 10762 2746
rect 10762 2694 10774 2746
rect 10774 2694 10804 2746
rect 10828 2694 10838 2746
rect 10838 2694 10884 2746
rect 10588 2692 10644 2694
rect 10668 2692 10724 2694
rect 10748 2692 10804 2694
rect 10828 2692 10884 2694
rect 20220 19610 20276 19612
rect 20300 19610 20356 19612
rect 20380 19610 20436 19612
rect 20460 19610 20516 19612
rect 20220 19558 20266 19610
rect 20266 19558 20276 19610
rect 20300 19558 20330 19610
rect 20330 19558 20342 19610
rect 20342 19558 20356 19610
rect 20380 19558 20394 19610
rect 20394 19558 20406 19610
rect 20406 19558 20436 19610
rect 20460 19558 20470 19610
rect 20470 19558 20516 19610
rect 20220 19556 20276 19558
rect 20300 19556 20356 19558
rect 20380 19556 20436 19558
rect 20460 19556 20516 19558
rect 20220 18522 20276 18524
rect 20300 18522 20356 18524
rect 20380 18522 20436 18524
rect 20460 18522 20516 18524
rect 20220 18470 20266 18522
rect 20266 18470 20276 18522
rect 20300 18470 20330 18522
rect 20330 18470 20342 18522
rect 20342 18470 20356 18522
rect 20380 18470 20394 18522
rect 20394 18470 20406 18522
rect 20406 18470 20436 18522
rect 20460 18470 20470 18522
rect 20470 18470 20516 18522
rect 20220 18468 20276 18470
rect 20300 18468 20356 18470
rect 20380 18468 20436 18470
rect 20460 18468 20516 18470
rect 20220 17434 20276 17436
rect 20300 17434 20356 17436
rect 20380 17434 20436 17436
rect 20460 17434 20516 17436
rect 20220 17382 20266 17434
rect 20266 17382 20276 17434
rect 20300 17382 20330 17434
rect 20330 17382 20342 17434
rect 20342 17382 20356 17434
rect 20380 17382 20394 17434
rect 20394 17382 20406 17434
rect 20406 17382 20436 17434
rect 20460 17382 20470 17434
rect 20470 17382 20516 17434
rect 20220 17380 20276 17382
rect 20300 17380 20356 17382
rect 20380 17380 20436 17382
rect 20460 17380 20516 17382
rect 20220 16346 20276 16348
rect 20300 16346 20356 16348
rect 20380 16346 20436 16348
rect 20460 16346 20516 16348
rect 20220 16294 20266 16346
rect 20266 16294 20276 16346
rect 20300 16294 20330 16346
rect 20330 16294 20342 16346
rect 20342 16294 20356 16346
rect 20380 16294 20394 16346
rect 20394 16294 20406 16346
rect 20406 16294 20436 16346
rect 20460 16294 20470 16346
rect 20470 16294 20516 16346
rect 20220 16292 20276 16294
rect 20300 16292 20356 16294
rect 20380 16292 20436 16294
rect 20460 16292 20516 16294
rect 20220 15258 20276 15260
rect 20300 15258 20356 15260
rect 20380 15258 20436 15260
rect 20460 15258 20516 15260
rect 20220 15206 20266 15258
rect 20266 15206 20276 15258
rect 20300 15206 20330 15258
rect 20330 15206 20342 15258
rect 20342 15206 20356 15258
rect 20380 15206 20394 15258
rect 20394 15206 20406 15258
rect 20406 15206 20436 15258
rect 20460 15206 20470 15258
rect 20470 15206 20516 15258
rect 20220 15204 20276 15206
rect 20300 15204 20356 15206
rect 20380 15204 20436 15206
rect 20460 15204 20516 15206
rect 20220 14170 20276 14172
rect 20300 14170 20356 14172
rect 20380 14170 20436 14172
rect 20460 14170 20516 14172
rect 20220 14118 20266 14170
rect 20266 14118 20276 14170
rect 20300 14118 20330 14170
rect 20330 14118 20342 14170
rect 20342 14118 20356 14170
rect 20380 14118 20394 14170
rect 20394 14118 20406 14170
rect 20406 14118 20436 14170
rect 20460 14118 20470 14170
rect 20470 14118 20516 14170
rect 20220 14116 20276 14118
rect 20300 14116 20356 14118
rect 20380 14116 20436 14118
rect 20460 14116 20516 14118
rect 20220 13082 20276 13084
rect 20300 13082 20356 13084
rect 20380 13082 20436 13084
rect 20460 13082 20516 13084
rect 20220 13030 20266 13082
rect 20266 13030 20276 13082
rect 20300 13030 20330 13082
rect 20330 13030 20342 13082
rect 20342 13030 20356 13082
rect 20380 13030 20394 13082
rect 20394 13030 20406 13082
rect 20406 13030 20436 13082
rect 20460 13030 20470 13082
rect 20470 13030 20516 13082
rect 20220 13028 20276 13030
rect 20300 13028 20356 13030
rect 20380 13028 20436 13030
rect 20460 13028 20516 13030
rect 20220 11994 20276 11996
rect 20300 11994 20356 11996
rect 20380 11994 20436 11996
rect 20460 11994 20516 11996
rect 20220 11942 20266 11994
rect 20266 11942 20276 11994
rect 20300 11942 20330 11994
rect 20330 11942 20342 11994
rect 20342 11942 20356 11994
rect 20380 11942 20394 11994
rect 20394 11942 20406 11994
rect 20406 11942 20436 11994
rect 20460 11942 20470 11994
rect 20470 11942 20516 11994
rect 20220 11940 20276 11942
rect 20300 11940 20356 11942
rect 20380 11940 20436 11942
rect 20460 11940 20516 11942
rect 20220 10906 20276 10908
rect 20300 10906 20356 10908
rect 20380 10906 20436 10908
rect 20460 10906 20516 10908
rect 20220 10854 20266 10906
rect 20266 10854 20276 10906
rect 20300 10854 20330 10906
rect 20330 10854 20342 10906
rect 20342 10854 20356 10906
rect 20380 10854 20394 10906
rect 20394 10854 20406 10906
rect 20406 10854 20436 10906
rect 20460 10854 20470 10906
rect 20470 10854 20516 10906
rect 20220 10852 20276 10854
rect 20300 10852 20356 10854
rect 20380 10852 20436 10854
rect 20460 10852 20516 10854
rect 20220 9818 20276 9820
rect 20300 9818 20356 9820
rect 20380 9818 20436 9820
rect 20460 9818 20516 9820
rect 20220 9766 20266 9818
rect 20266 9766 20276 9818
rect 20300 9766 20330 9818
rect 20330 9766 20342 9818
rect 20342 9766 20356 9818
rect 20380 9766 20394 9818
rect 20394 9766 20406 9818
rect 20406 9766 20436 9818
rect 20460 9766 20470 9818
rect 20470 9766 20516 9818
rect 20220 9764 20276 9766
rect 20300 9764 20356 9766
rect 20380 9764 20436 9766
rect 20460 9764 20516 9766
rect 20220 8730 20276 8732
rect 20300 8730 20356 8732
rect 20380 8730 20436 8732
rect 20460 8730 20516 8732
rect 20220 8678 20266 8730
rect 20266 8678 20276 8730
rect 20300 8678 20330 8730
rect 20330 8678 20342 8730
rect 20342 8678 20356 8730
rect 20380 8678 20394 8730
rect 20394 8678 20406 8730
rect 20406 8678 20436 8730
rect 20460 8678 20470 8730
rect 20470 8678 20516 8730
rect 20220 8676 20276 8678
rect 20300 8676 20356 8678
rect 20380 8676 20436 8678
rect 20460 8676 20516 8678
rect 20220 7642 20276 7644
rect 20300 7642 20356 7644
rect 20380 7642 20436 7644
rect 20460 7642 20516 7644
rect 20220 7590 20266 7642
rect 20266 7590 20276 7642
rect 20300 7590 20330 7642
rect 20330 7590 20342 7642
rect 20342 7590 20356 7642
rect 20380 7590 20394 7642
rect 20394 7590 20406 7642
rect 20406 7590 20436 7642
rect 20460 7590 20470 7642
rect 20470 7590 20516 7642
rect 20220 7588 20276 7590
rect 20300 7588 20356 7590
rect 20380 7588 20436 7590
rect 20460 7588 20516 7590
rect 20220 6554 20276 6556
rect 20300 6554 20356 6556
rect 20380 6554 20436 6556
rect 20460 6554 20516 6556
rect 20220 6502 20266 6554
rect 20266 6502 20276 6554
rect 20300 6502 20330 6554
rect 20330 6502 20342 6554
rect 20342 6502 20356 6554
rect 20380 6502 20394 6554
rect 20394 6502 20406 6554
rect 20406 6502 20436 6554
rect 20460 6502 20470 6554
rect 20470 6502 20516 6554
rect 20220 6500 20276 6502
rect 20300 6500 20356 6502
rect 20380 6500 20436 6502
rect 20460 6500 20516 6502
rect 20220 5466 20276 5468
rect 20300 5466 20356 5468
rect 20380 5466 20436 5468
rect 20460 5466 20516 5468
rect 20220 5414 20266 5466
rect 20266 5414 20276 5466
rect 20300 5414 20330 5466
rect 20330 5414 20342 5466
rect 20342 5414 20356 5466
rect 20380 5414 20394 5466
rect 20394 5414 20406 5466
rect 20406 5414 20436 5466
rect 20460 5414 20470 5466
rect 20470 5414 20516 5466
rect 20220 5412 20276 5414
rect 20300 5412 20356 5414
rect 20380 5412 20436 5414
rect 20460 5412 20516 5414
rect 20220 4378 20276 4380
rect 20300 4378 20356 4380
rect 20380 4378 20436 4380
rect 20460 4378 20516 4380
rect 20220 4326 20266 4378
rect 20266 4326 20276 4378
rect 20300 4326 20330 4378
rect 20330 4326 20342 4378
rect 20342 4326 20356 4378
rect 20380 4326 20394 4378
rect 20394 4326 20406 4378
rect 20406 4326 20436 4378
rect 20460 4326 20470 4378
rect 20470 4326 20516 4378
rect 20220 4324 20276 4326
rect 20300 4324 20356 4326
rect 20380 4324 20436 4326
rect 20460 4324 20516 4326
rect 20220 3290 20276 3292
rect 20300 3290 20356 3292
rect 20380 3290 20436 3292
rect 20460 3290 20516 3292
rect 20220 3238 20266 3290
rect 20266 3238 20276 3290
rect 20300 3238 20330 3290
rect 20330 3238 20342 3290
rect 20342 3238 20356 3290
rect 20380 3238 20394 3290
rect 20394 3238 20406 3290
rect 20406 3238 20436 3290
rect 20460 3238 20470 3290
rect 20470 3238 20516 3290
rect 20220 3236 20276 3238
rect 20300 3236 20356 3238
rect 20380 3236 20436 3238
rect 20460 3236 20516 3238
rect 29852 19066 29908 19068
rect 29932 19066 29988 19068
rect 30012 19066 30068 19068
rect 30092 19066 30148 19068
rect 29852 19014 29898 19066
rect 29898 19014 29908 19066
rect 29932 19014 29962 19066
rect 29962 19014 29974 19066
rect 29974 19014 29988 19066
rect 30012 19014 30026 19066
rect 30026 19014 30038 19066
rect 30038 19014 30068 19066
rect 30092 19014 30102 19066
rect 30102 19014 30148 19066
rect 29852 19012 29908 19014
rect 29932 19012 29988 19014
rect 30012 19012 30068 19014
rect 30092 19012 30148 19014
rect 29852 17978 29908 17980
rect 29932 17978 29988 17980
rect 30012 17978 30068 17980
rect 30092 17978 30148 17980
rect 29852 17926 29898 17978
rect 29898 17926 29908 17978
rect 29932 17926 29962 17978
rect 29962 17926 29974 17978
rect 29974 17926 29988 17978
rect 30012 17926 30026 17978
rect 30026 17926 30038 17978
rect 30038 17926 30068 17978
rect 30092 17926 30102 17978
rect 30102 17926 30148 17978
rect 29852 17924 29908 17926
rect 29932 17924 29988 17926
rect 30012 17924 30068 17926
rect 30092 17924 30148 17926
rect 29852 16890 29908 16892
rect 29932 16890 29988 16892
rect 30012 16890 30068 16892
rect 30092 16890 30148 16892
rect 29852 16838 29898 16890
rect 29898 16838 29908 16890
rect 29932 16838 29962 16890
rect 29962 16838 29974 16890
rect 29974 16838 29988 16890
rect 30012 16838 30026 16890
rect 30026 16838 30038 16890
rect 30038 16838 30068 16890
rect 30092 16838 30102 16890
rect 30102 16838 30148 16890
rect 29852 16836 29908 16838
rect 29932 16836 29988 16838
rect 30012 16836 30068 16838
rect 30092 16836 30148 16838
rect 29852 15802 29908 15804
rect 29932 15802 29988 15804
rect 30012 15802 30068 15804
rect 30092 15802 30148 15804
rect 29852 15750 29898 15802
rect 29898 15750 29908 15802
rect 29932 15750 29962 15802
rect 29962 15750 29974 15802
rect 29974 15750 29988 15802
rect 30012 15750 30026 15802
rect 30026 15750 30038 15802
rect 30038 15750 30068 15802
rect 30092 15750 30102 15802
rect 30102 15750 30148 15802
rect 29852 15748 29908 15750
rect 29932 15748 29988 15750
rect 30012 15748 30068 15750
rect 30092 15748 30148 15750
rect 29852 14714 29908 14716
rect 29932 14714 29988 14716
rect 30012 14714 30068 14716
rect 30092 14714 30148 14716
rect 29852 14662 29898 14714
rect 29898 14662 29908 14714
rect 29932 14662 29962 14714
rect 29962 14662 29974 14714
rect 29974 14662 29988 14714
rect 30012 14662 30026 14714
rect 30026 14662 30038 14714
rect 30038 14662 30068 14714
rect 30092 14662 30102 14714
rect 30102 14662 30148 14714
rect 29852 14660 29908 14662
rect 29932 14660 29988 14662
rect 30012 14660 30068 14662
rect 30092 14660 30148 14662
rect 29852 13626 29908 13628
rect 29932 13626 29988 13628
rect 30012 13626 30068 13628
rect 30092 13626 30148 13628
rect 29852 13574 29898 13626
rect 29898 13574 29908 13626
rect 29932 13574 29962 13626
rect 29962 13574 29974 13626
rect 29974 13574 29988 13626
rect 30012 13574 30026 13626
rect 30026 13574 30038 13626
rect 30038 13574 30068 13626
rect 30092 13574 30102 13626
rect 30102 13574 30148 13626
rect 29852 13572 29908 13574
rect 29932 13572 29988 13574
rect 30012 13572 30068 13574
rect 30092 13572 30148 13574
rect 29852 12538 29908 12540
rect 29932 12538 29988 12540
rect 30012 12538 30068 12540
rect 30092 12538 30148 12540
rect 29852 12486 29898 12538
rect 29898 12486 29908 12538
rect 29932 12486 29962 12538
rect 29962 12486 29974 12538
rect 29974 12486 29988 12538
rect 30012 12486 30026 12538
rect 30026 12486 30038 12538
rect 30038 12486 30068 12538
rect 30092 12486 30102 12538
rect 30102 12486 30148 12538
rect 29852 12484 29908 12486
rect 29932 12484 29988 12486
rect 30012 12484 30068 12486
rect 30092 12484 30148 12486
rect 29852 11450 29908 11452
rect 29932 11450 29988 11452
rect 30012 11450 30068 11452
rect 30092 11450 30148 11452
rect 29852 11398 29898 11450
rect 29898 11398 29908 11450
rect 29932 11398 29962 11450
rect 29962 11398 29974 11450
rect 29974 11398 29988 11450
rect 30012 11398 30026 11450
rect 30026 11398 30038 11450
rect 30038 11398 30068 11450
rect 30092 11398 30102 11450
rect 30102 11398 30148 11450
rect 29852 11396 29908 11398
rect 29932 11396 29988 11398
rect 30012 11396 30068 11398
rect 30092 11396 30148 11398
rect 29852 10362 29908 10364
rect 29932 10362 29988 10364
rect 30012 10362 30068 10364
rect 30092 10362 30148 10364
rect 29852 10310 29898 10362
rect 29898 10310 29908 10362
rect 29932 10310 29962 10362
rect 29962 10310 29974 10362
rect 29974 10310 29988 10362
rect 30012 10310 30026 10362
rect 30026 10310 30038 10362
rect 30038 10310 30068 10362
rect 30092 10310 30102 10362
rect 30102 10310 30148 10362
rect 29852 10308 29908 10310
rect 29932 10308 29988 10310
rect 30012 10308 30068 10310
rect 30092 10308 30148 10310
rect 29852 9274 29908 9276
rect 29932 9274 29988 9276
rect 30012 9274 30068 9276
rect 30092 9274 30148 9276
rect 29852 9222 29898 9274
rect 29898 9222 29908 9274
rect 29932 9222 29962 9274
rect 29962 9222 29974 9274
rect 29974 9222 29988 9274
rect 30012 9222 30026 9274
rect 30026 9222 30038 9274
rect 30038 9222 30068 9274
rect 30092 9222 30102 9274
rect 30102 9222 30148 9274
rect 29852 9220 29908 9222
rect 29932 9220 29988 9222
rect 30012 9220 30068 9222
rect 30092 9220 30148 9222
rect 29852 8186 29908 8188
rect 29932 8186 29988 8188
rect 30012 8186 30068 8188
rect 30092 8186 30148 8188
rect 29852 8134 29898 8186
rect 29898 8134 29908 8186
rect 29932 8134 29962 8186
rect 29962 8134 29974 8186
rect 29974 8134 29988 8186
rect 30012 8134 30026 8186
rect 30026 8134 30038 8186
rect 30038 8134 30068 8186
rect 30092 8134 30102 8186
rect 30102 8134 30148 8186
rect 29852 8132 29908 8134
rect 29932 8132 29988 8134
rect 30012 8132 30068 8134
rect 30092 8132 30148 8134
rect 29852 7098 29908 7100
rect 29932 7098 29988 7100
rect 30012 7098 30068 7100
rect 30092 7098 30148 7100
rect 29852 7046 29898 7098
rect 29898 7046 29908 7098
rect 29932 7046 29962 7098
rect 29962 7046 29974 7098
rect 29974 7046 29988 7098
rect 30012 7046 30026 7098
rect 30026 7046 30038 7098
rect 30038 7046 30068 7098
rect 30092 7046 30102 7098
rect 30102 7046 30148 7098
rect 29852 7044 29908 7046
rect 29932 7044 29988 7046
rect 30012 7044 30068 7046
rect 30092 7044 30148 7046
rect 29852 6010 29908 6012
rect 29932 6010 29988 6012
rect 30012 6010 30068 6012
rect 30092 6010 30148 6012
rect 29852 5958 29898 6010
rect 29898 5958 29908 6010
rect 29932 5958 29962 6010
rect 29962 5958 29974 6010
rect 29974 5958 29988 6010
rect 30012 5958 30026 6010
rect 30026 5958 30038 6010
rect 30038 5958 30068 6010
rect 30092 5958 30102 6010
rect 30102 5958 30148 6010
rect 29852 5956 29908 5958
rect 29932 5956 29988 5958
rect 30012 5956 30068 5958
rect 30092 5956 30148 5958
rect 29852 4922 29908 4924
rect 29932 4922 29988 4924
rect 30012 4922 30068 4924
rect 30092 4922 30148 4924
rect 29852 4870 29898 4922
rect 29898 4870 29908 4922
rect 29932 4870 29962 4922
rect 29962 4870 29974 4922
rect 29974 4870 29988 4922
rect 30012 4870 30026 4922
rect 30026 4870 30038 4922
rect 30038 4870 30068 4922
rect 30092 4870 30102 4922
rect 30102 4870 30148 4922
rect 29852 4868 29908 4870
rect 29932 4868 29988 4870
rect 30012 4868 30068 4870
rect 30092 4868 30148 4870
rect 29852 3834 29908 3836
rect 29932 3834 29988 3836
rect 30012 3834 30068 3836
rect 30092 3834 30148 3836
rect 29852 3782 29898 3834
rect 29898 3782 29908 3834
rect 29932 3782 29962 3834
rect 29962 3782 29974 3834
rect 29974 3782 29988 3834
rect 30012 3782 30026 3834
rect 30026 3782 30038 3834
rect 30038 3782 30068 3834
rect 30092 3782 30102 3834
rect 30102 3782 30148 3834
rect 29852 3780 29908 3782
rect 29932 3780 29988 3782
rect 30012 3780 30068 3782
rect 30092 3780 30148 3782
rect 29852 2746 29908 2748
rect 29932 2746 29988 2748
rect 30012 2746 30068 2748
rect 30092 2746 30148 2748
rect 29852 2694 29898 2746
rect 29898 2694 29908 2746
rect 29932 2694 29962 2746
rect 29962 2694 29974 2746
rect 29974 2694 29988 2746
rect 30012 2694 30026 2746
rect 30026 2694 30038 2746
rect 30038 2694 30068 2746
rect 30092 2694 30102 2746
rect 30102 2694 30148 2746
rect 29852 2692 29908 2694
rect 29932 2692 29988 2694
rect 30012 2692 30068 2694
rect 30092 2692 30148 2694
rect 39484 19610 39540 19612
rect 39564 19610 39620 19612
rect 39644 19610 39700 19612
rect 39724 19610 39780 19612
rect 39484 19558 39530 19610
rect 39530 19558 39540 19610
rect 39564 19558 39594 19610
rect 39594 19558 39606 19610
rect 39606 19558 39620 19610
rect 39644 19558 39658 19610
rect 39658 19558 39670 19610
rect 39670 19558 39700 19610
rect 39724 19558 39734 19610
rect 39734 19558 39780 19610
rect 39484 19556 39540 19558
rect 39564 19556 39620 19558
rect 39644 19556 39700 19558
rect 39724 19556 39780 19558
rect 39484 18522 39540 18524
rect 39564 18522 39620 18524
rect 39644 18522 39700 18524
rect 39724 18522 39780 18524
rect 39484 18470 39530 18522
rect 39530 18470 39540 18522
rect 39564 18470 39594 18522
rect 39594 18470 39606 18522
rect 39606 18470 39620 18522
rect 39644 18470 39658 18522
rect 39658 18470 39670 18522
rect 39670 18470 39700 18522
rect 39724 18470 39734 18522
rect 39734 18470 39780 18522
rect 39484 18468 39540 18470
rect 39564 18468 39620 18470
rect 39644 18468 39700 18470
rect 39724 18468 39780 18470
rect 39484 17434 39540 17436
rect 39564 17434 39620 17436
rect 39644 17434 39700 17436
rect 39724 17434 39780 17436
rect 39484 17382 39530 17434
rect 39530 17382 39540 17434
rect 39564 17382 39594 17434
rect 39594 17382 39606 17434
rect 39606 17382 39620 17434
rect 39644 17382 39658 17434
rect 39658 17382 39670 17434
rect 39670 17382 39700 17434
rect 39724 17382 39734 17434
rect 39734 17382 39780 17434
rect 39484 17380 39540 17382
rect 39564 17380 39620 17382
rect 39644 17380 39700 17382
rect 39724 17380 39780 17382
rect 39484 16346 39540 16348
rect 39564 16346 39620 16348
rect 39644 16346 39700 16348
rect 39724 16346 39780 16348
rect 39484 16294 39530 16346
rect 39530 16294 39540 16346
rect 39564 16294 39594 16346
rect 39594 16294 39606 16346
rect 39606 16294 39620 16346
rect 39644 16294 39658 16346
rect 39658 16294 39670 16346
rect 39670 16294 39700 16346
rect 39724 16294 39734 16346
rect 39734 16294 39780 16346
rect 39484 16292 39540 16294
rect 39564 16292 39620 16294
rect 39644 16292 39700 16294
rect 39724 16292 39780 16294
rect 39484 15258 39540 15260
rect 39564 15258 39620 15260
rect 39644 15258 39700 15260
rect 39724 15258 39780 15260
rect 39484 15206 39530 15258
rect 39530 15206 39540 15258
rect 39564 15206 39594 15258
rect 39594 15206 39606 15258
rect 39606 15206 39620 15258
rect 39644 15206 39658 15258
rect 39658 15206 39670 15258
rect 39670 15206 39700 15258
rect 39724 15206 39734 15258
rect 39734 15206 39780 15258
rect 39484 15204 39540 15206
rect 39564 15204 39620 15206
rect 39644 15204 39700 15206
rect 39724 15204 39780 15206
rect 55954 21664 56010 21720
rect 39484 14170 39540 14172
rect 39564 14170 39620 14172
rect 39644 14170 39700 14172
rect 39724 14170 39780 14172
rect 39484 14118 39530 14170
rect 39530 14118 39540 14170
rect 39564 14118 39594 14170
rect 39594 14118 39606 14170
rect 39606 14118 39620 14170
rect 39644 14118 39658 14170
rect 39658 14118 39670 14170
rect 39670 14118 39700 14170
rect 39724 14118 39734 14170
rect 39734 14118 39780 14170
rect 39484 14116 39540 14118
rect 39564 14116 39620 14118
rect 39644 14116 39700 14118
rect 39724 14116 39780 14118
rect 39484 13082 39540 13084
rect 39564 13082 39620 13084
rect 39644 13082 39700 13084
rect 39724 13082 39780 13084
rect 39484 13030 39530 13082
rect 39530 13030 39540 13082
rect 39564 13030 39594 13082
rect 39594 13030 39606 13082
rect 39606 13030 39620 13082
rect 39644 13030 39658 13082
rect 39658 13030 39670 13082
rect 39670 13030 39700 13082
rect 39724 13030 39734 13082
rect 39734 13030 39780 13082
rect 39484 13028 39540 13030
rect 39564 13028 39620 13030
rect 39644 13028 39700 13030
rect 39724 13028 39780 13030
rect 39484 11994 39540 11996
rect 39564 11994 39620 11996
rect 39644 11994 39700 11996
rect 39724 11994 39780 11996
rect 39484 11942 39530 11994
rect 39530 11942 39540 11994
rect 39564 11942 39594 11994
rect 39594 11942 39606 11994
rect 39606 11942 39620 11994
rect 39644 11942 39658 11994
rect 39658 11942 39670 11994
rect 39670 11942 39700 11994
rect 39724 11942 39734 11994
rect 39734 11942 39780 11994
rect 39484 11940 39540 11942
rect 39564 11940 39620 11942
rect 39644 11940 39700 11942
rect 39724 11940 39780 11942
rect 39484 10906 39540 10908
rect 39564 10906 39620 10908
rect 39644 10906 39700 10908
rect 39724 10906 39780 10908
rect 39484 10854 39530 10906
rect 39530 10854 39540 10906
rect 39564 10854 39594 10906
rect 39594 10854 39606 10906
rect 39606 10854 39620 10906
rect 39644 10854 39658 10906
rect 39658 10854 39670 10906
rect 39670 10854 39700 10906
rect 39724 10854 39734 10906
rect 39734 10854 39780 10906
rect 39484 10852 39540 10854
rect 39564 10852 39620 10854
rect 39644 10852 39700 10854
rect 39724 10852 39780 10854
rect 39484 9818 39540 9820
rect 39564 9818 39620 9820
rect 39644 9818 39700 9820
rect 39724 9818 39780 9820
rect 39484 9766 39530 9818
rect 39530 9766 39540 9818
rect 39564 9766 39594 9818
rect 39594 9766 39606 9818
rect 39606 9766 39620 9818
rect 39644 9766 39658 9818
rect 39658 9766 39670 9818
rect 39670 9766 39700 9818
rect 39724 9766 39734 9818
rect 39734 9766 39780 9818
rect 39484 9764 39540 9766
rect 39564 9764 39620 9766
rect 39644 9764 39700 9766
rect 39724 9764 39780 9766
rect 39484 8730 39540 8732
rect 39564 8730 39620 8732
rect 39644 8730 39700 8732
rect 39724 8730 39780 8732
rect 39484 8678 39530 8730
rect 39530 8678 39540 8730
rect 39564 8678 39594 8730
rect 39594 8678 39606 8730
rect 39606 8678 39620 8730
rect 39644 8678 39658 8730
rect 39658 8678 39670 8730
rect 39670 8678 39700 8730
rect 39724 8678 39734 8730
rect 39734 8678 39780 8730
rect 39484 8676 39540 8678
rect 39564 8676 39620 8678
rect 39644 8676 39700 8678
rect 39724 8676 39780 8678
rect 39484 7642 39540 7644
rect 39564 7642 39620 7644
rect 39644 7642 39700 7644
rect 39724 7642 39780 7644
rect 39484 7590 39530 7642
rect 39530 7590 39540 7642
rect 39564 7590 39594 7642
rect 39594 7590 39606 7642
rect 39606 7590 39620 7642
rect 39644 7590 39658 7642
rect 39658 7590 39670 7642
rect 39670 7590 39700 7642
rect 39724 7590 39734 7642
rect 39734 7590 39780 7642
rect 39484 7588 39540 7590
rect 39564 7588 39620 7590
rect 39644 7588 39700 7590
rect 39724 7588 39780 7590
rect 39484 6554 39540 6556
rect 39564 6554 39620 6556
rect 39644 6554 39700 6556
rect 39724 6554 39780 6556
rect 39484 6502 39530 6554
rect 39530 6502 39540 6554
rect 39564 6502 39594 6554
rect 39594 6502 39606 6554
rect 39606 6502 39620 6554
rect 39644 6502 39658 6554
rect 39658 6502 39670 6554
rect 39670 6502 39700 6554
rect 39724 6502 39734 6554
rect 39734 6502 39780 6554
rect 39484 6500 39540 6502
rect 39564 6500 39620 6502
rect 39644 6500 39700 6502
rect 39724 6500 39780 6502
rect 39484 5466 39540 5468
rect 39564 5466 39620 5468
rect 39644 5466 39700 5468
rect 39724 5466 39780 5468
rect 39484 5414 39530 5466
rect 39530 5414 39540 5466
rect 39564 5414 39594 5466
rect 39594 5414 39606 5466
rect 39606 5414 39620 5466
rect 39644 5414 39658 5466
rect 39658 5414 39670 5466
rect 39670 5414 39700 5466
rect 39724 5414 39734 5466
rect 39734 5414 39780 5466
rect 39484 5412 39540 5414
rect 39564 5412 39620 5414
rect 39644 5412 39700 5414
rect 39724 5412 39780 5414
rect 39484 4378 39540 4380
rect 39564 4378 39620 4380
rect 39644 4378 39700 4380
rect 39724 4378 39780 4380
rect 39484 4326 39530 4378
rect 39530 4326 39540 4378
rect 39564 4326 39594 4378
rect 39594 4326 39606 4378
rect 39606 4326 39620 4378
rect 39644 4326 39658 4378
rect 39658 4326 39670 4378
rect 39670 4326 39700 4378
rect 39724 4326 39734 4378
rect 39734 4326 39780 4378
rect 39484 4324 39540 4326
rect 39564 4324 39620 4326
rect 39644 4324 39700 4326
rect 39724 4324 39780 4326
rect 39484 3290 39540 3292
rect 39564 3290 39620 3292
rect 39644 3290 39700 3292
rect 39724 3290 39780 3292
rect 39484 3238 39530 3290
rect 39530 3238 39540 3290
rect 39564 3238 39594 3290
rect 39594 3238 39606 3290
rect 39606 3238 39620 3290
rect 39644 3238 39658 3290
rect 39658 3238 39670 3290
rect 39670 3238 39700 3290
rect 39724 3238 39734 3290
rect 39734 3238 39780 3290
rect 39484 3236 39540 3238
rect 39564 3236 39620 3238
rect 39644 3236 39700 3238
rect 39724 3236 39780 3238
rect 49116 19066 49172 19068
rect 49196 19066 49252 19068
rect 49276 19066 49332 19068
rect 49356 19066 49412 19068
rect 49116 19014 49162 19066
rect 49162 19014 49172 19066
rect 49196 19014 49226 19066
rect 49226 19014 49238 19066
rect 49238 19014 49252 19066
rect 49276 19014 49290 19066
rect 49290 19014 49302 19066
rect 49302 19014 49332 19066
rect 49356 19014 49366 19066
rect 49366 19014 49412 19066
rect 49116 19012 49172 19014
rect 49196 19012 49252 19014
rect 49276 19012 49332 19014
rect 49356 19012 49412 19014
rect 49116 17978 49172 17980
rect 49196 17978 49252 17980
rect 49276 17978 49332 17980
rect 49356 17978 49412 17980
rect 49116 17926 49162 17978
rect 49162 17926 49172 17978
rect 49196 17926 49226 17978
rect 49226 17926 49238 17978
rect 49238 17926 49252 17978
rect 49276 17926 49290 17978
rect 49290 17926 49302 17978
rect 49302 17926 49332 17978
rect 49356 17926 49366 17978
rect 49366 17926 49412 17978
rect 49116 17924 49172 17926
rect 49196 17924 49252 17926
rect 49276 17924 49332 17926
rect 49356 17924 49412 17926
rect 49116 16890 49172 16892
rect 49196 16890 49252 16892
rect 49276 16890 49332 16892
rect 49356 16890 49412 16892
rect 49116 16838 49162 16890
rect 49162 16838 49172 16890
rect 49196 16838 49226 16890
rect 49226 16838 49238 16890
rect 49238 16838 49252 16890
rect 49276 16838 49290 16890
rect 49290 16838 49302 16890
rect 49302 16838 49332 16890
rect 49356 16838 49366 16890
rect 49366 16838 49412 16890
rect 49116 16836 49172 16838
rect 49196 16836 49252 16838
rect 49276 16836 49332 16838
rect 49356 16836 49412 16838
rect 49116 15802 49172 15804
rect 49196 15802 49252 15804
rect 49276 15802 49332 15804
rect 49356 15802 49412 15804
rect 49116 15750 49162 15802
rect 49162 15750 49172 15802
rect 49196 15750 49226 15802
rect 49226 15750 49238 15802
rect 49238 15750 49252 15802
rect 49276 15750 49290 15802
rect 49290 15750 49302 15802
rect 49302 15750 49332 15802
rect 49356 15750 49366 15802
rect 49366 15750 49412 15802
rect 49116 15748 49172 15750
rect 49196 15748 49252 15750
rect 49276 15748 49332 15750
rect 49356 15748 49412 15750
rect 49116 14714 49172 14716
rect 49196 14714 49252 14716
rect 49276 14714 49332 14716
rect 49356 14714 49412 14716
rect 49116 14662 49162 14714
rect 49162 14662 49172 14714
rect 49196 14662 49226 14714
rect 49226 14662 49238 14714
rect 49238 14662 49252 14714
rect 49276 14662 49290 14714
rect 49290 14662 49302 14714
rect 49302 14662 49332 14714
rect 49356 14662 49366 14714
rect 49366 14662 49412 14714
rect 49116 14660 49172 14662
rect 49196 14660 49252 14662
rect 49276 14660 49332 14662
rect 49356 14660 49412 14662
rect 49116 13626 49172 13628
rect 49196 13626 49252 13628
rect 49276 13626 49332 13628
rect 49356 13626 49412 13628
rect 49116 13574 49162 13626
rect 49162 13574 49172 13626
rect 49196 13574 49226 13626
rect 49226 13574 49238 13626
rect 49238 13574 49252 13626
rect 49276 13574 49290 13626
rect 49290 13574 49302 13626
rect 49302 13574 49332 13626
rect 49356 13574 49366 13626
rect 49366 13574 49412 13626
rect 49116 13572 49172 13574
rect 49196 13572 49252 13574
rect 49276 13572 49332 13574
rect 49356 13572 49412 13574
rect 49116 12538 49172 12540
rect 49196 12538 49252 12540
rect 49276 12538 49332 12540
rect 49356 12538 49412 12540
rect 49116 12486 49162 12538
rect 49162 12486 49172 12538
rect 49196 12486 49226 12538
rect 49226 12486 49238 12538
rect 49238 12486 49252 12538
rect 49276 12486 49290 12538
rect 49290 12486 49302 12538
rect 49302 12486 49332 12538
rect 49356 12486 49366 12538
rect 49366 12486 49412 12538
rect 49116 12484 49172 12486
rect 49196 12484 49252 12486
rect 49276 12484 49332 12486
rect 49356 12484 49412 12486
rect 49116 11450 49172 11452
rect 49196 11450 49252 11452
rect 49276 11450 49332 11452
rect 49356 11450 49412 11452
rect 49116 11398 49162 11450
rect 49162 11398 49172 11450
rect 49196 11398 49226 11450
rect 49226 11398 49238 11450
rect 49238 11398 49252 11450
rect 49276 11398 49290 11450
rect 49290 11398 49302 11450
rect 49302 11398 49332 11450
rect 49356 11398 49366 11450
rect 49366 11398 49412 11450
rect 49116 11396 49172 11398
rect 49196 11396 49252 11398
rect 49276 11396 49332 11398
rect 49356 11396 49412 11398
rect 49116 10362 49172 10364
rect 49196 10362 49252 10364
rect 49276 10362 49332 10364
rect 49356 10362 49412 10364
rect 49116 10310 49162 10362
rect 49162 10310 49172 10362
rect 49196 10310 49226 10362
rect 49226 10310 49238 10362
rect 49238 10310 49252 10362
rect 49276 10310 49290 10362
rect 49290 10310 49302 10362
rect 49302 10310 49332 10362
rect 49356 10310 49366 10362
rect 49366 10310 49412 10362
rect 49116 10308 49172 10310
rect 49196 10308 49252 10310
rect 49276 10308 49332 10310
rect 49356 10308 49412 10310
rect 49116 9274 49172 9276
rect 49196 9274 49252 9276
rect 49276 9274 49332 9276
rect 49356 9274 49412 9276
rect 49116 9222 49162 9274
rect 49162 9222 49172 9274
rect 49196 9222 49226 9274
rect 49226 9222 49238 9274
rect 49238 9222 49252 9274
rect 49276 9222 49290 9274
rect 49290 9222 49302 9274
rect 49302 9222 49332 9274
rect 49356 9222 49366 9274
rect 49366 9222 49412 9274
rect 49116 9220 49172 9222
rect 49196 9220 49252 9222
rect 49276 9220 49332 9222
rect 49356 9220 49412 9222
rect 49116 8186 49172 8188
rect 49196 8186 49252 8188
rect 49276 8186 49332 8188
rect 49356 8186 49412 8188
rect 49116 8134 49162 8186
rect 49162 8134 49172 8186
rect 49196 8134 49226 8186
rect 49226 8134 49238 8186
rect 49238 8134 49252 8186
rect 49276 8134 49290 8186
rect 49290 8134 49302 8186
rect 49302 8134 49332 8186
rect 49356 8134 49366 8186
rect 49366 8134 49412 8186
rect 49116 8132 49172 8134
rect 49196 8132 49252 8134
rect 49276 8132 49332 8134
rect 49356 8132 49412 8134
rect 49116 7098 49172 7100
rect 49196 7098 49252 7100
rect 49276 7098 49332 7100
rect 49356 7098 49412 7100
rect 49116 7046 49162 7098
rect 49162 7046 49172 7098
rect 49196 7046 49226 7098
rect 49226 7046 49238 7098
rect 49238 7046 49252 7098
rect 49276 7046 49290 7098
rect 49290 7046 49302 7098
rect 49302 7046 49332 7098
rect 49356 7046 49366 7098
rect 49366 7046 49412 7098
rect 49116 7044 49172 7046
rect 49196 7044 49252 7046
rect 49276 7044 49332 7046
rect 49356 7044 49412 7046
rect 49116 6010 49172 6012
rect 49196 6010 49252 6012
rect 49276 6010 49332 6012
rect 49356 6010 49412 6012
rect 49116 5958 49162 6010
rect 49162 5958 49172 6010
rect 49196 5958 49226 6010
rect 49226 5958 49238 6010
rect 49238 5958 49252 6010
rect 49276 5958 49290 6010
rect 49290 5958 49302 6010
rect 49302 5958 49332 6010
rect 49356 5958 49366 6010
rect 49366 5958 49412 6010
rect 49116 5956 49172 5958
rect 49196 5956 49252 5958
rect 49276 5956 49332 5958
rect 49356 5956 49412 5958
rect 49116 4922 49172 4924
rect 49196 4922 49252 4924
rect 49276 4922 49332 4924
rect 49356 4922 49412 4924
rect 49116 4870 49162 4922
rect 49162 4870 49172 4922
rect 49196 4870 49226 4922
rect 49226 4870 49238 4922
rect 49238 4870 49252 4922
rect 49276 4870 49290 4922
rect 49290 4870 49302 4922
rect 49302 4870 49332 4922
rect 49356 4870 49366 4922
rect 49366 4870 49412 4922
rect 49116 4868 49172 4870
rect 49196 4868 49252 4870
rect 49276 4868 49332 4870
rect 49356 4868 49412 4870
rect 49116 3834 49172 3836
rect 49196 3834 49252 3836
rect 49276 3834 49332 3836
rect 49356 3834 49412 3836
rect 49116 3782 49162 3834
rect 49162 3782 49172 3834
rect 49196 3782 49226 3834
rect 49226 3782 49238 3834
rect 49238 3782 49252 3834
rect 49276 3782 49290 3834
rect 49290 3782 49302 3834
rect 49302 3782 49332 3834
rect 49356 3782 49366 3834
rect 49366 3782 49412 3834
rect 49116 3780 49172 3782
rect 49196 3780 49252 3782
rect 49276 3780 49332 3782
rect 49356 3780 49412 3782
rect 20220 2202 20276 2204
rect 20300 2202 20356 2204
rect 20380 2202 20436 2204
rect 20460 2202 20516 2204
rect 20220 2150 20266 2202
rect 20266 2150 20276 2202
rect 20300 2150 20330 2202
rect 20330 2150 20342 2202
rect 20342 2150 20356 2202
rect 20380 2150 20394 2202
rect 20394 2150 20406 2202
rect 20406 2150 20436 2202
rect 20460 2150 20470 2202
rect 20470 2150 20516 2202
rect 20220 2148 20276 2150
rect 20300 2148 20356 2150
rect 20380 2148 20436 2150
rect 20460 2148 20516 2150
rect 39484 2202 39540 2204
rect 39564 2202 39620 2204
rect 39644 2202 39700 2204
rect 39724 2202 39780 2204
rect 39484 2150 39530 2202
rect 39530 2150 39540 2202
rect 39564 2150 39594 2202
rect 39594 2150 39606 2202
rect 39606 2150 39620 2202
rect 39644 2150 39658 2202
rect 39658 2150 39670 2202
rect 39670 2150 39700 2202
rect 39724 2150 39734 2202
rect 39734 2150 39780 2202
rect 39484 2148 39540 2150
rect 39564 2148 39620 2150
rect 39644 2148 39700 2150
rect 39724 2148 39780 2150
rect 49116 2746 49172 2748
rect 49196 2746 49252 2748
rect 49276 2746 49332 2748
rect 49356 2746 49412 2748
rect 49116 2694 49162 2746
rect 49162 2694 49172 2746
rect 49196 2694 49226 2746
rect 49226 2694 49238 2746
rect 49238 2694 49252 2746
rect 49276 2694 49290 2746
rect 49290 2694 49302 2746
rect 49302 2694 49332 2746
rect 49356 2694 49366 2746
rect 49366 2694 49412 2746
rect 49116 2692 49172 2694
rect 49196 2692 49252 2694
rect 49276 2692 49332 2694
rect 49356 2692 49412 2694
rect 55770 20032 55826 20088
rect 56230 21120 56286 21176
rect 56046 20576 56102 20632
rect 56506 19624 56562 19680
rect 56506 4664 56562 4720
rect 56506 4256 56562 4312
rect 56046 3168 56102 3224
rect 55770 2624 55826 2680
rect 55586 2216 55642 2272
rect 57242 19116 57244 19136
rect 57244 19116 57296 19136
rect 57296 19116 57298 19136
rect 57242 19080 57298 19116
rect 56874 5208 56930 5264
rect 57242 17060 57298 17096
rect 57242 17040 57244 17060
rect 57244 17040 57296 17060
rect 57296 17040 57298 17060
rect 57886 18536 57942 18592
rect 57242 10412 57244 10432
rect 57244 10412 57296 10432
rect 57296 10412 57298 10432
rect 57242 10376 57298 10412
rect 58070 17992 58126 18048
rect 57886 17584 57942 17640
rect 58070 16496 58126 16552
rect 58070 15952 58126 16008
rect 58070 15544 58126 15600
rect 57886 15000 57942 15056
rect 58070 14456 58126 14512
rect 58070 13912 58126 13968
rect 57886 13368 57942 13424
rect 58070 12960 58126 13016
rect 58070 12416 58126 12472
rect 58070 11872 58126 11928
rect 58070 11328 58126 11384
rect 57886 10920 57942 10976
rect 58070 9832 58126 9888
rect 57886 9288 57942 9344
rect 58070 8880 58126 8936
rect 58070 8336 58126 8392
rect 57886 7792 57942 7848
rect 58070 7248 58126 7304
rect 58070 6704 58126 6760
rect 58070 6296 58126 6352
rect 58070 5752 58126 5808
rect 56506 1128 56562 1184
rect 55218 176 55274 232
rect 57794 3712 57850 3768
rect 57150 1672 57206 1728
rect 56966 584 57022 640
<< metal3 >>
rect 55949 21722 56015 21725
rect 59200 21722 60000 21752
rect 55949 21720 60000 21722
rect 55949 21664 55954 21720
rect 56010 21664 60000 21720
rect 55949 21662 60000 21664
rect 55949 21659 56015 21662
rect 59200 21632 60000 21662
rect 56225 21178 56291 21181
rect 59200 21178 60000 21208
rect 56225 21176 60000 21178
rect 56225 21120 56230 21176
rect 56286 21120 60000 21176
rect 56225 21118 60000 21120
rect 56225 21115 56291 21118
rect 59200 21088 60000 21118
rect 56041 20634 56107 20637
rect 59200 20634 60000 20664
rect 56041 20632 60000 20634
rect 56041 20576 56046 20632
rect 56102 20576 60000 20632
rect 56041 20574 60000 20576
rect 56041 20571 56107 20574
rect 59200 20544 60000 20574
rect 55765 20090 55831 20093
rect 59200 20090 60000 20120
rect 55765 20088 60000 20090
rect 55765 20032 55770 20088
rect 55826 20032 60000 20088
rect 55765 20030 60000 20032
rect 55765 20027 55831 20030
rect 59200 20000 60000 20030
rect 56501 19682 56567 19685
rect 59200 19682 60000 19712
rect 56501 19680 60000 19682
rect 56501 19624 56506 19680
rect 56562 19624 60000 19680
rect 56501 19622 60000 19624
rect 56501 19619 56567 19622
rect 20208 19616 20528 19617
rect 20208 19552 20216 19616
rect 20280 19552 20296 19616
rect 20360 19552 20376 19616
rect 20440 19552 20456 19616
rect 20520 19552 20528 19616
rect 20208 19551 20528 19552
rect 39472 19616 39792 19617
rect 39472 19552 39480 19616
rect 39544 19552 39560 19616
rect 39624 19552 39640 19616
rect 39704 19552 39720 19616
rect 39784 19552 39792 19616
rect 59200 19592 60000 19622
rect 39472 19551 39792 19552
rect 57237 19138 57303 19141
rect 59200 19138 60000 19168
rect 57237 19136 60000 19138
rect 57237 19080 57242 19136
rect 57298 19080 60000 19136
rect 57237 19078 60000 19080
rect 57237 19075 57303 19078
rect 10576 19072 10896 19073
rect 10576 19008 10584 19072
rect 10648 19008 10664 19072
rect 10728 19008 10744 19072
rect 10808 19008 10824 19072
rect 10888 19008 10896 19072
rect 10576 19007 10896 19008
rect 29840 19072 30160 19073
rect 29840 19008 29848 19072
rect 29912 19008 29928 19072
rect 29992 19008 30008 19072
rect 30072 19008 30088 19072
rect 30152 19008 30160 19072
rect 29840 19007 30160 19008
rect 49104 19072 49424 19073
rect 49104 19008 49112 19072
rect 49176 19008 49192 19072
rect 49256 19008 49272 19072
rect 49336 19008 49352 19072
rect 49416 19008 49424 19072
rect 59200 19048 60000 19078
rect 49104 19007 49424 19008
rect 57881 18594 57947 18597
rect 59200 18594 60000 18624
rect 57881 18592 60000 18594
rect 57881 18536 57886 18592
rect 57942 18536 60000 18592
rect 57881 18534 60000 18536
rect 57881 18531 57947 18534
rect 20208 18528 20528 18529
rect 20208 18464 20216 18528
rect 20280 18464 20296 18528
rect 20360 18464 20376 18528
rect 20440 18464 20456 18528
rect 20520 18464 20528 18528
rect 20208 18463 20528 18464
rect 39472 18528 39792 18529
rect 39472 18464 39480 18528
rect 39544 18464 39560 18528
rect 39624 18464 39640 18528
rect 39704 18464 39720 18528
rect 39784 18464 39792 18528
rect 59200 18504 60000 18534
rect 39472 18463 39792 18464
rect 58065 18050 58131 18053
rect 59200 18050 60000 18080
rect 58065 18048 60000 18050
rect 58065 17992 58070 18048
rect 58126 17992 60000 18048
rect 58065 17990 60000 17992
rect 58065 17987 58131 17990
rect 10576 17984 10896 17985
rect 10576 17920 10584 17984
rect 10648 17920 10664 17984
rect 10728 17920 10744 17984
rect 10808 17920 10824 17984
rect 10888 17920 10896 17984
rect 10576 17919 10896 17920
rect 29840 17984 30160 17985
rect 29840 17920 29848 17984
rect 29912 17920 29928 17984
rect 29992 17920 30008 17984
rect 30072 17920 30088 17984
rect 30152 17920 30160 17984
rect 29840 17919 30160 17920
rect 49104 17984 49424 17985
rect 49104 17920 49112 17984
rect 49176 17920 49192 17984
rect 49256 17920 49272 17984
rect 49336 17920 49352 17984
rect 49416 17920 49424 17984
rect 59200 17960 60000 17990
rect 49104 17919 49424 17920
rect 57881 17642 57947 17645
rect 59200 17642 60000 17672
rect 57881 17640 60000 17642
rect 57881 17584 57886 17640
rect 57942 17584 60000 17640
rect 57881 17582 60000 17584
rect 57881 17579 57947 17582
rect 59200 17552 60000 17582
rect 20208 17440 20528 17441
rect 20208 17376 20216 17440
rect 20280 17376 20296 17440
rect 20360 17376 20376 17440
rect 20440 17376 20456 17440
rect 20520 17376 20528 17440
rect 20208 17375 20528 17376
rect 39472 17440 39792 17441
rect 39472 17376 39480 17440
rect 39544 17376 39560 17440
rect 39624 17376 39640 17440
rect 39704 17376 39720 17440
rect 39784 17376 39792 17440
rect 39472 17375 39792 17376
rect 57237 17098 57303 17101
rect 59200 17098 60000 17128
rect 57237 17096 60000 17098
rect 57237 17040 57242 17096
rect 57298 17040 60000 17096
rect 57237 17038 60000 17040
rect 57237 17035 57303 17038
rect 59200 17008 60000 17038
rect 10576 16896 10896 16897
rect 10576 16832 10584 16896
rect 10648 16832 10664 16896
rect 10728 16832 10744 16896
rect 10808 16832 10824 16896
rect 10888 16832 10896 16896
rect 10576 16831 10896 16832
rect 29840 16896 30160 16897
rect 29840 16832 29848 16896
rect 29912 16832 29928 16896
rect 29992 16832 30008 16896
rect 30072 16832 30088 16896
rect 30152 16832 30160 16896
rect 29840 16831 30160 16832
rect 49104 16896 49424 16897
rect 49104 16832 49112 16896
rect 49176 16832 49192 16896
rect 49256 16832 49272 16896
rect 49336 16832 49352 16896
rect 49416 16832 49424 16896
rect 49104 16831 49424 16832
rect 58065 16554 58131 16557
rect 59200 16554 60000 16584
rect 58065 16552 60000 16554
rect 58065 16496 58070 16552
rect 58126 16496 60000 16552
rect 58065 16494 60000 16496
rect 58065 16491 58131 16494
rect 59200 16464 60000 16494
rect 20208 16352 20528 16353
rect 20208 16288 20216 16352
rect 20280 16288 20296 16352
rect 20360 16288 20376 16352
rect 20440 16288 20456 16352
rect 20520 16288 20528 16352
rect 20208 16287 20528 16288
rect 39472 16352 39792 16353
rect 39472 16288 39480 16352
rect 39544 16288 39560 16352
rect 39624 16288 39640 16352
rect 39704 16288 39720 16352
rect 39784 16288 39792 16352
rect 39472 16287 39792 16288
rect 58065 16010 58131 16013
rect 59200 16010 60000 16040
rect 58065 16008 60000 16010
rect 58065 15952 58070 16008
rect 58126 15952 60000 16008
rect 58065 15950 60000 15952
rect 58065 15947 58131 15950
rect 59200 15920 60000 15950
rect 10576 15808 10896 15809
rect 10576 15744 10584 15808
rect 10648 15744 10664 15808
rect 10728 15744 10744 15808
rect 10808 15744 10824 15808
rect 10888 15744 10896 15808
rect 10576 15743 10896 15744
rect 29840 15808 30160 15809
rect 29840 15744 29848 15808
rect 29912 15744 29928 15808
rect 29992 15744 30008 15808
rect 30072 15744 30088 15808
rect 30152 15744 30160 15808
rect 29840 15743 30160 15744
rect 49104 15808 49424 15809
rect 49104 15744 49112 15808
rect 49176 15744 49192 15808
rect 49256 15744 49272 15808
rect 49336 15744 49352 15808
rect 49416 15744 49424 15808
rect 49104 15743 49424 15744
rect 58065 15602 58131 15605
rect 59200 15602 60000 15632
rect 58065 15600 60000 15602
rect 58065 15544 58070 15600
rect 58126 15544 60000 15600
rect 58065 15542 60000 15544
rect 58065 15539 58131 15542
rect 59200 15512 60000 15542
rect 20208 15264 20528 15265
rect 20208 15200 20216 15264
rect 20280 15200 20296 15264
rect 20360 15200 20376 15264
rect 20440 15200 20456 15264
rect 20520 15200 20528 15264
rect 20208 15199 20528 15200
rect 39472 15264 39792 15265
rect 39472 15200 39480 15264
rect 39544 15200 39560 15264
rect 39624 15200 39640 15264
rect 39704 15200 39720 15264
rect 39784 15200 39792 15264
rect 39472 15199 39792 15200
rect 57881 15058 57947 15061
rect 59200 15058 60000 15088
rect 57881 15056 60000 15058
rect 57881 15000 57886 15056
rect 57942 15000 60000 15056
rect 57881 14998 60000 15000
rect 57881 14995 57947 14998
rect 59200 14968 60000 14998
rect 10576 14720 10896 14721
rect 10576 14656 10584 14720
rect 10648 14656 10664 14720
rect 10728 14656 10744 14720
rect 10808 14656 10824 14720
rect 10888 14656 10896 14720
rect 10576 14655 10896 14656
rect 29840 14720 30160 14721
rect 29840 14656 29848 14720
rect 29912 14656 29928 14720
rect 29992 14656 30008 14720
rect 30072 14656 30088 14720
rect 30152 14656 30160 14720
rect 29840 14655 30160 14656
rect 49104 14720 49424 14721
rect 49104 14656 49112 14720
rect 49176 14656 49192 14720
rect 49256 14656 49272 14720
rect 49336 14656 49352 14720
rect 49416 14656 49424 14720
rect 49104 14655 49424 14656
rect 58065 14514 58131 14517
rect 59200 14514 60000 14544
rect 58065 14512 60000 14514
rect 58065 14456 58070 14512
rect 58126 14456 60000 14512
rect 58065 14454 60000 14456
rect 58065 14451 58131 14454
rect 59200 14424 60000 14454
rect 20208 14176 20528 14177
rect 20208 14112 20216 14176
rect 20280 14112 20296 14176
rect 20360 14112 20376 14176
rect 20440 14112 20456 14176
rect 20520 14112 20528 14176
rect 20208 14111 20528 14112
rect 39472 14176 39792 14177
rect 39472 14112 39480 14176
rect 39544 14112 39560 14176
rect 39624 14112 39640 14176
rect 39704 14112 39720 14176
rect 39784 14112 39792 14176
rect 39472 14111 39792 14112
rect 58065 13970 58131 13973
rect 59200 13970 60000 14000
rect 58065 13968 60000 13970
rect 58065 13912 58070 13968
rect 58126 13912 60000 13968
rect 58065 13910 60000 13912
rect 58065 13907 58131 13910
rect 59200 13880 60000 13910
rect 10576 13632 10896 13633
rect 10576 13568 10584 13632
rect 10648 13568 10664 13632
rect 10728 13568 10744 13632
rect 10808 13568 10824 13632
rect 10888 13568 10896 13632
rect 10576 13567 10896 13568
rect 29840 13632 30160 13633
rect 29840 13568 29848 13632
rect 29912 13568 29928 13632
rect 29992 13568 30008 13632
rect 30072 13568 30088 13632
rect 30152 13568 30160 13632
rect 29840 13567 30160 13568
rect 49104 13632 49424 13633
rect 49104 13568 49112 13632
rect 49176 13568 49192 13632
rect 49256 13568 49272 13632
rect 49336 13568 49352 13632
rect 49416 13568 49424 13632
rect 49104 13567 49424 13568
rect 57881 13426 57947 13429
rect 59200 13426 60000 13456
rect 57881 13424 60000 13426
rect 57881 13368 57886 13424
rect 57942 13368 60000 13424
rect 57881 13366 60000 13368
rect 57881 13363 57947 13366
rect 59200 13336 60000 13366
rect 20208 13088 20528 13089
rect 20208 13024 20216 13088
rect 20280 13024 20296 13088
rect 20360 13024 20376 13088
rect 20440 13024 20456 13088
rect 20520 13024 20528 13088
rect 20208 13023 20528 13024
rect 39472 13088 39792 13089
rect 39472 13024 39480 13088
rect 39544 13024 39560 13088
rect 39624 13024 39640 13088
rect 39704 13024 39720 13088
rect 39784 13024 39792 13088
rect 39472 13023 39792 13024
rect 58065 13018 58131 13021
rect 59200 13018 60000 13048
rect 58065 13016 60000 13018
rect 58065 12960 58070 13016
rect 58126 12960 60000 13016
rect 58065 12958 60000 12960
rect 58065 12955 58131 12958
rect 59200 12928 60000 12958
rect 10576 12544 10896 12545
rect 10576 12480 10584 12544
rect 10648 12480 10664 12544
rect 10728 12480 10744 12544
rect 10808 12480 10824 12544
rect 10888 12480 10896 12544
rect 10576 12479 10896 12480
rect 29840 12544 30160 12545
rect 29840 12480 29848 12544
rect 29912 12480 29928 12544
rect 29992 12480 30008 12544
rect 30072 12480 30088 12544
rect 30152 12480 30160 12544
rect 29840 12479 30160 12480
rect 49104 12544 49424 12545
rect 49104 12480 49112 12544
rect 49176 12480 49192 12544
rect 49256 12480 49272 12544
rect 49336 12480 49352 12544
rect 49416 12480 49424 12544
rect 49104 12479 49424 12480
rect 58065 12474 58131 12477
rect 59200 12474 60000 12504
rect 58065 12472 60000 12474
rect 58065 12416 58070 12472
rect 58126 12416 60000 12472
rect 58065 12414 60000 12416
rect 58065 12411 58131 12414
rect 59200 12384 60000 12414
rect 20208 12000 20528 12001
rect 20208 11936 20216 12000
rect 20280 11936 20296 12000
rect 20360 11936 20376 12000
rect 20440 11936 20456 12000
rect 20520 11936 20528 12000
rect 20208 11935 20528 11936
rect 39472 12000 39792 12001
rect 39472 11936 39480 12000
rect 39544 11936 39560 12000
rect 39624 11936 39640 12000
rect 39704 11936 39720 12000
rect 39784 11936 39792 12000
rect 39472 11935 39792 11936
rect 58065 11930 58131 11933
rect 59200 11930 60000 11960
rect 58065 11928 60000 11930
rect 58065 11872 58070 11928
rect 58126 11872 60000 11928
rect 58065 11870 60000 11872
rect 58065 11867 58131 11870
rect 59200 11840 60000 11870
rect 10576 11456 10896 11457
rect 10576 11392 10584 11456
rect 10648 11392 10664 11456
rect 10728 11392 10744 11456
rect 10808 11392 10824 11456
rect 10888 11392 10896 11456
rect 10576 11391 10896 11392
rect 29840 11456 30160 11457
rect 29840 11392 29848 11456
rect 29912 11392 29928 11456
rect 29992 11392 30008 11456
rect 30072 11392 30088 11456
rect 30152 11392 30160 11456
rect 29840 11391 30160 11392
rect 49104 11456 49424 11457
rect 49104 11392 49112 11456
rect 49176 11392 49192 11456
rect 49256 11392 49272 11456
rect 49336 11392 49352 11456
rect 49416 11392 49424 11456
rect 49104 11391 49424 11392
rect 58065 11386 58131 11389
rect 59200 11386 60000 11416
rect 58065 11384 60000 11386
rect 58065 11328 58070 11384
rect 58126 11328 60000 11384
rect 58065 11326 60000 11328
rect 58065 11323 58131 11326
rect 59200 11296 60000 11326
rect 57881 10978 57947 10981
rect 59200 10978 60000 11008
rect 57881 10976 60000 10978
rect 57881 10920 57886 10976
rect 57942 10920 60000 10976
rect 57881 10918 60000 10920
rect 57881 10915 57947 10918
rect 20208 10912 20528 10913
rect 20208 10848 20216 10912
rect 20280 10848 20296 10912
rect 20360 10848 20376 10912
rect 20440 10848 20456 10912
rect 20520 10848 20528 10912
rect 20208 10847 20528 10848
rect 39472 10912 39792 10913
rect 39472 10848 39480 10912
rect 39544 10848 39560 10912
rect 39624 10848 39640 10912
rect 39704 10848 39720 10912
rect 39784 10848 39792 10912
rect 59200 10888 60000 10918
rect 39472 10847 39792 10848
rect 57237 10434 57303 10437
rect 59200 10434 60000 10464
rect 57237 10432 60000 10434
rect 57237 10376 57242 10432
rect 57298 10376 60000 10432
rect 57237 10374 60000 10376
rect 57237 10371 57303 10374
rect 10576 10368 10896 10369
rect 10576 10304 10584 10368
rect 10648 10304 10664 10368
rect 10728 10304 10744 10368
rect 10808 10304 10824 10368
rect 10888 10304 10896 10368
rect 10576 10303 10896 10304
rect 29840 10368 30160 10369
rect 29840 10304 29848 10368
rect 29912 10304 29928 10368
rect 29992 10304 30008 10368
rect 30072 10304 30088 10368
rect 30152 10304 30160 10368
rect 29840 10303 30160 10304
rect 49104 10368 49424 10369
rect 49104 10304 49112 10368
rect 49176 10304 49192 10368
rect 49256 10304 49272 10368
rect 49336 10304 49352 10368
rect 49416 10304 49424 10368
rect 59200 10344 60000 10374
rect 49104 10303 49424 10304
rect 58065 9890 58131 9893
rect 59200 9890 60000 9920
rect 58065 9888 60000 9890
rect 58065 9832 58070 9888
rect 58126 9832 60000 9888
rect 58065 9830 60000 9832
rect 58065 9827 58131 9830
rect 20208 9824 20528 9825
rect 20208 9760 20216 9824
rect 20280 9760 20296 9824
rect 20360 9760 20376 9824
rect 20440 9760 20456 9824
rect 20520 9760 20528 9824
rect 20208 9759 20528 9760
rect 39472 9824 39792 9825
rect 39472 9760 39480 9824
rect 39544 9760 39560 9824
rect 39624 9760 39640 9824
rect 39704 9760 39720 9824
rect 39784 9760 39792 9824
rect 59200 9800 60000 9830
rect 39472 9759 39792 9760
rect 57881 9346 57947 9349
rect 59200 9346 60000 9376
rect 57881 9344 60000 9346
rect 57881 9288 57886 9344
rect 57942 9288 60000 9344
rect 57881 9286 60000 9288
rect 57881 9283 57947 9286
rect 10576 9280 10896 9281
rect 10576 9216 10584 9280
rect 10648 9216 10664 9280
rect 10728 9216 10744 9280
rect 10808 9216 10824 9280
rect 10888 9216 10896 9280
rect 10576 9215 10896 9216
rect 29840 9280 30160 9281
rect 29840 9216 29848 9280
rect 29912 9216 29928 9280
rect 29992 9216 30008 9280
rect 30072 9216 30088 9280
rect 30152 9216 30160 9280
rect 29840 9215 30160 9216
rect 49104 9280 49424 9281
rect 49104 9216 49112 9280
rect 49176 9216 49192 9280
rect 49256 9216 49272 9280
rect 49336 9216 49352 9280
rect 49416 9216 49424 9280
rect 59200 9256 60000 9286
rect 49104 9215 49424 9216
rect 58065 8938 58131 8941
rect 59200 8938 60000 8968
rect 58065 8936 60000 8938
rect 58065 8880 58070 8936
rect 58126 8880 60000 8936
rect 58065 8878 60000 8880
rect 58065 8875 58131 8878
rect 59200 8848 60000 8878
rect 20208 8736 20528 8737
rect 20208 8672 20216 8736
rect 20280 8672 20296 8736
rect 20360 8672 20376 8736
rect 20440 8672 20456 8736
rect 20520 8672 20528 8736
rect 20208 8671 20528 8672
rect 39472 8736 39792 8737
rect 39472 8672 39480 8736
rect 39544 8672 39560 8736
rect 39624 8672 39640 8736
rect 39704 8672 39720 8736
rect 39784 8672 39792 8736
rect 39472 8671 39792 8672
rect 58065 8394 58131 8397
rect 59200 8394 60000 8424
rect 58065 8392 60000 8394
rect 58065 8336 58070 8392
rect 58126 8336 60000 8392
rect 58065 8334 60000 8336
rect 58065 8331 58131 8334
rect 59200 8304 60000 8334
rect 10576 8192 10896 8193
rect 10576 8128 10584 8192
rect 10648 8128 10664 8192
rect 10728 8128 10744 8192
rect 10808 8128 10824 8192
rect 10888 8128 10896 8192
rect 10576 8127 10896 8128
rect 29840 8192 30160 8193
rect 29840 8128 29848 8192
rect 29912 8128 29928 8192
rect 29992 8128 30008 8192
rect 30072 8128 30088 8192
rect 30152 8128 30160 8192
rect 29840 8127 30160 8128
rect 49104 8192 49424 8193
rect 49104 8128 49112 8192
rect 49176 8128 49192 8192
rect 49256 8128 49272 8192
rect 49336 8128 49352 8192
rect 49416 8128 49424 8192
rect 49104 8127 49424 8128
rect 57881 7850 57947 7853
rect 59200 7850 60000 7880
rect 57881 7848 60000 7850
rect 57881 7792 57886 7848
rect 57942 7792 60000 7848
rect 57881 7790 60000 7792
rect 57881 7787 57947 7790
rect 59200 7760 60000 7790
rect 20208 7648 20528 7649
rect 20208 7584 20216 7648
rect 20280 7584 20296 7648
rect 20360 7584 20376 7648
rect 20440 7584 20456 7648
rect 20520 7584 20528 7648
rect 20208 7583 20528 7584
rect 39472 7648 39792 7649
rect 39472 7584 39480 7648
rect 39544 7584 39560 7648
rect 39624 7584 39640 7648
rect 39704 7584 39720 7648
rect 39784 7584 39792 7648
rect 39472 7583 39792 7584
rect 58065 7306 58131 7309
rect 59200 7306 60000 7336
rect 58065 7304 60000 7306
rect 58065 7248 58070 7304
rect 58126 7248 60000 7304
rect 58065 7246 60000 7248
rect 58065 7243 58131 7246
rect 59200 7216 60000 7246
rect 10576 7104 10896 7105
rect 10576 7040 10584 7104
rect 10648 7040 10664 7104
rect 10728 7040 10744 7104
rect 10808 7040 10824 7104
rect 10888 7040 10896 7104
rect 10576 7039 10896 7040
rect 29840 7104 30160 7105
rect 29840 7040 29848 7104
rect 29912 7040 29928 7104
rect 29992 7040 30008 7104
rect 30072 7040 30088 7104
rect 30152 7040 30160 7104
rect 29840 7039 30160 7040
rect 49104 7104 49424 7105
rect 49104 7040 49112 7104
rect 49176 7040 49192 7104
rect 49256 7040 49272 7104
rect 49336 7040 49352 7104
rect 49416 7040 49424 7104
rect 49104 7039 49424 7040
rect 58065 6762 58131 6765
rect 59200 6762 60000 6792
rect 58065 6760 60000 6762
rect 58065 6704 58070 6760
rect 58126 6704 60000 6760
rect 58065 6702 60000 6704
rect 58065 6699 58131 6702
rect 59200 6672 60000 6702
rect 20208 6560 20528 6561
rect 20208 6496 20216 6560
rect 20280 6496 20296 6560
rect 20360 6496 20376 6560
rect 20440 6496 20456 6560
rect 20520 6496 20528 6560
rect 20208 6495 20528 6496
rect 39472 6560 39792 6561
rect 39472 6496 39480 6560
rect 39544 6496 39560 6560
rect 39624 6496 39640 6560
rect 39704 6496 39720 6560
rect 39784 6496 39792 6560
rect 39472 6495 39792 6496
rect 58065 6354 58131 6357
rect 59200 6354 60000 6384
rect 58065 6352 60000 6354
rect 58065 6296 58070 6352
rect 58126 6296 60000 6352
rect 58065 6294 60000 6296
rect 58065 6291 58131 6294
rect 59200 6264 60000 6294
rect 10576 6016 10896 6017
rect 10576 5952 10584 6016
rect 10648 5952 10664 6016
rect 10728 5952 10744 6016
rect 10808 5952 10824 6016
rect 10888 5952 10896 6016
rect 10576 5951 10896 5952
rect 29840 6016 30160 6017
rect 29840 5952 29848 6016
rect 29912 5952 29928 6016
rect 29992 5952 30008 6016
rect 30072 5952 30088 6016
rect 30152 5952 30160 6016
rect 29840 5951 30160 5952
rect 49104 6016 49424 6017
rect 49104 5952 49112 6016
rect 49176 5952 49192 6016
rect 49256 5952 49272 6016
rect 49336 5952 49352 6016
rect 49416 5952 49424 6016
rect 49104 5951 49424 5952
rect 58065 5810 58131 5813
rect 59200 5810 60000 5840
rect 58065 5808 60000 5810
rect 58065 5752 58070 5808
rect 58126 5752 60000 5808
rect 58065 5750 60000 5752
rect 58065 5747 58131 5750
rect 59200 5720 60000 5750
rect 20208 5472 20528 5473
rect 20208 5408 20216 5472
rect 20280 5408 20296 5472
rect 20360 5408 20376 5472
rect 20440 5408 20456 5472
rect 20520 5408 20528 5472
rect 20208 5407 20528 5408
rect 39472 5472 39792 5473
rect 39472 5408 39480 5472
rect 39544 5408 39560 5472
rect 39624 5408 39640 5472
rect 39704 5408 39720 5472
rect 39784 5408 39792 5472
rect 39472 5407 39792 5408
rect 56869 5266 56935 5269
rect 59200 5266 60000 5296
rect 56869 5264 60000 5266
rect 56869 5208 56874 5264
rect 56930 5208 60000 5264
rect 56869 5206 60000 5208
rect 56869 5203 56935 5206
rect 59200 5176 60000 5206
rect 10576 4928 10896 4929
rect 10576 4864 10584 4928
rect 10648 4864 10664 4928
rect 10728 4864 10744 4928
rect 10808 4864 10824 4928
rect 10888 4864 10896 4928
rect 10576 4863 10896 4864
rect 29840 4928 30160 4929
rect 29840 4864 29848 4928
rect 29912 4864 29928 4928
rect 29992 4864 30008 4928
rect 30072 4864 30088 4928
rect 30152 4864 30160 4928
rect 29840 4863 30160 4864
rect 49104 4928 49424 4929
rect 49104 4864 49112 4928
rect 49176 4864 49192 4928
rect 49256 4864 49272 4928
rect 49336 4864 49352 4928
rect 49416 4864 49424 4928
rect 49104 4863 49424 4864
rect 56501 4722 56567 4725
rect 59200 4722 60000 4752
rect 56501 4720 60000 4722
rect 56501 4664 56506 4720
rect 56562 4664 60000 4720
rect 56501 4662 60000 4664
rect 56501 4659 56567 4662
rect 59200 4632 60000 4662
rect 20208 4384 20528 4385
rect 20208 4320 20216 4384
rect 20280 4320 20296 4384
rect 20360 4320 20376 4384
rect 20440 4320 20456 4384
rect 20520 4320 20528 4384
rect 20208 4319 20528 4320
rect 39472 4384 39792 4385
rect 39472 4320 39480 4384
rect 39544 4320 39560 4384
rect 39624 4320 39640 4384
rect 39704 4320 39720 4384
rect 39784 4320 39792 4384
rect 39472 4319 39792 4320
rect 56501 4314 56567 4317
rect 59200 4314 60000 4344
rect 56501 4312 60000 4314
rect 56501 4256 56506 4312
rect 56562 4256 60000 4312
rect 56501 4254 60000 4256
rect 56501 4251 56567 4254
rect 59200 4224 60000 4254
rect 10576 3840 10896 3841
rect 10576 3776 10584 3840
rect 10648 3776 10664 3840
rect 10728 3776 10744 3840
rect 10808 3776 10824 3840
rect 10888 3776 10896 3840
rect 10576 3775 10896 3776
rect 29840 3840 30160 3841
rect 29840 3776 29848 3840
rect 29912 3776 29928 3840
rect 29992 3776 30008 3840
rect 30072 3776 30088 3840
rect 30152 3776 30160 3840
rect 29840 3775 30160 3776
rect 49104 3840 49424 3841
rect 49104 3776 49112 3840
rect 49176 3776 49192 3840
rect 49256 3776 49272 3840
rect 49336 3776 49352 3840
rect 49416 3776 49424 3840
rect 49104 3775 49424 3776
rect 57789 3770 57855 3773
rect 59200 3770 60000 3800
rect 57789 3768 60000 3770
rect 57789 3712 57794 3768
rect 57850 3712 60000 3768
rect 57789 3710 60000 3712
rect 57789 3707 57855 3710
rect 59200 3680 60000 3710
rect 20208 3296 20528 3297
rect 20208 3232 20216 3296
rect 20280 3232 20296 3296
rect 20360 3232 20376 3296
rect 20440 3232 20456 3296
rect 20520 3232 20528 3296
rect 20208 3231 20528 3232
rect 39472 3296 39792 3297
rect 39472 3232 39480 3296
rect 39544 3232 39560 3296
rect 39624 3232 39640 3296
rect 39704 3232 39720 3296
rect 39784 3232 39792 3296
rect 39472 3231 39792 3232
rect 56041 3226 56107 3229
rect 59200 3226 60000 3256
rect 56041 3224 60000 3226
rect 56041 3168 56046 3224
rect 56102 3168 60000 3224
rect 56041 3166 60000 3168
rect 56041 3163 56107 3166
rect 59200 3136 60000 3166
rect 10576 2752 10896 2753
rect 10576 2688 10584 2752
rect 10648 2688 10664 2752
rect 10728 2688 10744 2752
rect 10808 2688 10824 2752
rect 10888 2688 10896 2752
rect 10576 2687 10896 2688
rect 29840 2752 30160 2753
rect 29840 2688 29848 2752
rect 29912 2688 29928 2752
rect 29992 2688 30008 2752
rect 30072 2688 30088 2752
rect 30152 2688 30160 2752
rect 29840 2687 30160 2688
rect 49104 2752 49424 2753
rect 49104 2688 49112 2752
rect 49176 2688 49192 2752
rect 49256 2688 49272 2752
rect 49336 2688 49352 2752
rect 49416 2688 49424 2752
rect 49104 2687 49424 2688
rect 55765 2682 55831 2685
rect 59200 2682 60000 2712
rect 55765 2680 60000 2682
rect 55765 2624 55770 2680
rect 55826 2624 60000 2680
rect 55765 2622 60000 2624
rect 55765 2619 55831 2622
rect 59200 2592 60000 2622
rect 55581 2274 55647 2277
rect 59200 2274 60000 2304
rect 55581 2272 60000 2274
rect 55581 2216 55586 2272
rect 55642 2216 60000 2272
rect 55581 2214 60000 2216
rect 55581 2211 55647 2214
rect 20208 2208 20528 2209
rect 20208 2144 20216 2208
rect 20280 2144 20296 2208
rect 20360 2144 20376 2208
rect 20440 2144 20456 2208
rect 20520 2144 20528 2208
rect 20208 2143 20528 2144
rect 39472 2208 39792 2209
rect 39472 2144 39480 2208
rect 39544 2144 39560 2208
rect 39624 2144 39640 2208
rect 39704 2144 39720 2208
rect 39784 2144 39792 2208
rect 59200 2184 60000 2214
rect 39472 2143 39792 2144
rect 57145 1730 57211 1733
rect 59200 1730 60000 1760
rect 57145 1728 60000 1730
rect 57145 1672 57150 1728
rect 57206 1672 60000 1728
rect 57145 1670 60000 1672
rect 57145 1667 57211 1670
rect 59200 1640 60000 1670
rect 56501 1186 56567 1189
rect 59200 1186 60000 1216
rect 56501 1184 60000 1186
rect 56501 1128 56506 1184
rect 56562 1128 60000 1184
rect 56501 1126 60000 1128
rect 56501 1123 56567 1126
rect 59200 1096 60000 1126
rect 56961 642 57027 645
rect 59200 642 60000 672
rect 56961 640 60000 642
rect 56961 584 56966 640
rect 57022 584 60000 640
rect 56961 582 60000 584
rect 56961 579 57027 582
rect 59200 552 60000 582
rect 55213 234 55279 237
rect 59200 234 60000 264
rect 55213 232 60000 234
rect 55213 176 55218 232
rect 55274 176 60000 232
rect 55213 174 60000 176
rect 55213 171 55279 174
rect 59200 144 60000 174
<< via3 >>
rect 20216 19612 20280 19616
rect 20216 19556 20220 19612
rect 20220 19556 20276 19612
rect 20276 19556 20280 19612
rect 20216 19552 20280 19556
rect 20296 19612 20360 19616
rect 20296 19556 20300 19612
rect 20300 19556 20356 19612
rect 20356 19556 20360 19612
rect 20296 19552 20360 19556
rect 20376 19612 20440 19616
rect 20376 19556 20380 19612
rect 20380 19556 20436 19612
rect 20436 19556 20440 19612
rect 20376 19552 20440 19556
rect 20456 19612 20520 19616
rect 20456 19556 20460 19612
rect 20460 19556 20516 19612
rect 20516 19556 20520 19612
rect 20456 19552 20520 19556
rect 39480 19612 39544 19616
rect 39480 19556 39484 19612
rect 39484 19556 39540 19612
rect 39540 19556 39544 19612
rect 39480 19552 39544 19556
rect 39560 19612 39624 19616
rect 39560 19556 39564 19612
rect 39564 19556 39620 19612
rect 39620 19556 39624 19612
rect 39560 19552 39624 19556
rect 39640 19612 39704 19616
rect 39640 19556 39644 19612
rect 39644 19556 39700 19612
rect 39700 19556 39704 19612
rect 39640 19552 39704 19556
rect 39720 19612 39784 19616
rect 39720 19556 39724 19612
rect 39724 19556 39780 19612
rect 39780 19556 39784 19612
rect 39720 19552 39784 19556
rect 10584 19068 10648 19072
rect 10584 19012 10588 19068
rect 10588 19012 10644 19068
rect 10644 19012 10648 19068
rect 10584 19008 10648 19012
rect 10664 19068 10728 19072
rect 10664 19012 10668 19068
rect 10668 19012 10724 19068
rect 10724 19012 10728 19068
rect 10664 19008 10728 19012
rect 10744 19068 10808 19072
rect 10744 19012 10748 19068
rect 10748 19012 10804 19068
rect 10804 19012 10808 19068
rect 10744 19008 10808 19012
rect 10824 19068 10888 19072
rect 10824 19012 10828 19068
rect 10828 19012 10884 19068
rect 10884 19012 10888 19068
rect 10824 19008 10888 19012
rect 29848 19068 29912 19072
rect 29848 19012 29852 19068
rect 29852 19012 29908 19068
rect 29908 19012 29912 19068
rect 29848 19008 29912 19012
rect 29928 19068 29992 19072
rect 29928 19012 29932 19068
rect 29932 19012 29988 19068
rect 29988 19012 29992 19068
rect 29928 19008 29992 19012
rect 30008 19068 30072 19072
rect 30008 19012 30012 19068
rect 30012 19012 30068 19068
rect 30068 19012 30072 19068
rect 30008 19008 30072 19012
rect 30088 19068 30152 19072
rect 30088 19012 30092 19068
rect 30092 19012 30148 19068
rect 30148 19012 30152 19068
rect 30088 19008 30152 19012
rect 49112 19068 49176 19072
rect 49112 19012 49116 19068
rect 49116 19012 49172 19068
rect 49172 19012 49176 19068
rect 49112 19008 49176 19012
rect 49192 19068 49256 19072
rect 49192 19012 49196 19068
rect 49196 19012 49252 19068
rect 49252 19012 49256 19068
rect 49192 19008 49256 19012
rect 49272 19068 49336 19072
rect 49272 19012 49276 19068
rect 49276 19012 49332 19068
rect 49332 19012 49336 19068
rect 49272 19008 49336 19012
rect 49352 19068 49416 19072
rect 49352 19012 49356 19068
rect 49356 19012 49412 19068
rect 49412 19012 49416 19068
rect 49352 19008 49416 19012
rect 20216 18524 20280 18528
rect 20216 18468 20220 18524
rect 20220 18468 20276 18524
rect 20276 18468 20280 18524
rect 20216 18464 20280 18468
rect 20296 18524 20360 18528
rect 20296 18468 20300 18524
rect 20300 18468 20356 18524
rect 20356 18468 20360 18524
rect 20296 18464 20360 18468
rect 20376 18524 20440 18528
rect 20376 18468 20380 18524
rect 20380 18468 20436 18524
rect 20436 18468 20440 18524
rect 20376 18464 20440 18468
rect 20456 18524 20520 18528
rect 20456 18468 20460 18524
rect 20460 18468 20516 18524
rect 20516 18468 20520 18524
rect 20456 18464 20520 18468
rect 39480 18524 39544 18528
rect 39480 18468 39484 18524
rect 39484 18468 39540 18524
rect 39540 18468 39544 18524
rect 39480 18464 39544 18468
rect 39560 18524 39624 18528
rect 39560 18468 39564 18524
rect 39564 18468 39620 18524
rect 39620 18468 39624 18524
rect 39560 18464 39624 18468
rect 39640 18524 39704 18528
rect 39640 18468 39644 18524
rect 39644 18468 39700 18524
rect 39700 18468 39704 18524
rect 39640 18464 39704 18468
rect 39720 18524 39784 18528
rect 39720 18468 39724 18524
rect 39724 18468 39780 18524
rect 39780 18468 39784 18524
rect 39720 18464 39784 18468
rect 10584 17980 10648 17984
rect 10584 17924 10588 17980
rect 10588 17924 10644 17980
rect 10644 17924 10648 17980
rect 10584 17920 10648 17924
rect 10664 17980 10728 17984
rect 10664 17924 10668 17980
rect 10668 17924 10724 17980
rect 10724 17924 10728 17980
rect 10664 17920 10728 17924
rect 10744 17980 10808 17984
rect 10744 17924 10748 17980
rect 10748 17924 10804 17980
rect 10804 17924 10808 17980
rect 10744 17920 10808 17924
rect 10824 17980 10888 17984
rect 10824 17924 10828 17980
rect 10828 17924 10884 17980
rect 10884 17924 10888 17980
rect 10824 17920 10888 17924
rect 29848 17980 29912 17984
rect 29848 17924 29852 17980
rect 29852 17924 29908 17980
rect 29908 17924 29912 17980
rect 29848 17920 29912 17924
rect 29928 17980 29992 17984
rect 29928 17924 29932 17980
rect 29932 17924 29988 17980
rect 29988 17924 29992 17980
rect 29928 17920 29992 17924
rect 30008 17980 30072 17984
rect 30008 17924 30012 17980
rect 30012 17924 30068 17980
rect 30068 17924 30072 17980
rect 30008 17920 30072 17924
rect 30088 17980 30152 17984
rect 30088 17924 30092 17980
rect 30092 17924 30148 17980
rect 30148 17924 30152 17980
rect 30088 17920 30152 17924
rect 49112 17980 49176 17984
rect 49112 17924 49116 17980
rect 49116 17924 49172 17980
rect 49172 17924 49176 17980
rect 49112 17920 49176 17924
rect 49192 17980 49256 17984
rect 49192 17924 49196 17980
rect 49196 17924 49252 17980
rect 49252 17924 49256 17980
rect 49192 17920 49256 17924
rect 49272 17980 49336 17984
rect 49272 17924 49276 17980
rect 49276 17924 49332 17980
rect 49332 17924 49336 17980
rect 49272 17920 49336 17924
rect 49352 17980 49416 17984
rect 49352 17924 49356 17980
rect 49356 17924 49412 17980
rect 49412 17924 49416 17980
rect 49352 17920 49416 17924
rect 20216 17436 20280 17440
rect 20216 17380 20220 17436
rect 20220 17380 20276 17436
rect 20276 17380 20280 17436
rect 20216 17376 20280 17380
rect 20296 17436 20360 17440
rect 20296 17380 20300 17436
rect 20300 17380 20356 17436
rect 20356 17380 20360 17436
rect 20296 17376 20360 17380
rect 20376 17436 20440 17440
rect 20376 17380 20380 17436
rect 20380 17380 20436 17436
rect 20436 17380 20440 17436
rect 20376 17376 20440 17380
rect 20456 17436 20520 17440
rect 20456 17380 20460 17436
rect 20460 17380 20516 17436
rect 20516 17380 20520 17436
rect 20456 17376 20520 17380
rect 39480 17436 39544 17440
rect 39480 17380 39484 17436
rect 39484 17380 39540 17436
rect 39540 17380 39544 17436
rect 39480 17376 39544 17380
rect 39560 17436 39624 17440
rect 39560 17380 39564 17436
rect 39564 17380 39620 17436
rect 39620 17380 39624 17436
rect 39560 17376 39624 17380
rect 39640 17436 39704 17440
rect 39640 17380 39644 17436
rect 39644 17380 39700 17436
rect 39700 17380 39704 17436
rect 39640 17376 39704 17380
rect 39720 17436 39784 17440
rect 39720 17380 39724 17436
rect 39724 17380 39780 17436
rect 39780 17380 39784 17436
rect 39720 17376 39784 17380
rect 10584 16892 10648 16896
rect 10584 16836 10588 16892
rect 10588 16836 10644 16892
rect 10644 16836 10648 16892
rect 10584 16832 10648 16836
rect 10664 16892 10728 16896
rect 10664 16836 10668 16892
rect 10668 16836 10724 16892
rect 10724 16836 10728 16892
rect 10664 16832 10728 16836
rect 10744 16892 10808 16896
rect 10744 16836 10748 16892
rect 10748 16836 10804 16892
rect 10804 16836 10808 16892
rect 10744 16832 10808 16836
rect 10824 16892 10888 16896
rect 10824 16836 10828 16892
rect 10828 16836 10884 16892
rect 10884 16836 10888 16892
rect 10824 16832 10888 16836
rect 29848 16892 29912 16896
rect 29848 16836 29852 16892
rect 29852 16836 29908 16892
rect 29908 16836 29912 16892
rect 29848 16832 29912 16836
rect 29928 16892 29992 16896
rect 29928 16836 29932 16892
rect 29932 16836 29988 16892
rect 29988 16836 29992 16892
rect 29928 16832 29992 16836
rect 30008 16892 30072 16896
rect 30008 16836 30012 16892
rect 30012 16836 30068 16892
rect 30068 16836 30072 16892
rect 30008 16832 30072 16836
rect 30088 16892 30152 16896
rect 30088 16836 30092 16892
rect 30092 16836 30148 16892
rect 30148 16836 30152 16892
rect 30088 16832 30152 16836
rect 49112 16892 49176 16896
rect 49112 16836 49116 16892
rect 49116 16836 49172 16892
rect 49172 16836 49176 16892
rect 49112 16832 49176 16836
rect 49192 16892 49256 16896
rect 49192 16836 49196 16892
rect 49196 16836 49252 16892
rect 49252 16836 49256 16892
rect 49192 16832 49256 16836
rect 49272 16892 49336 16896
rect 49272 16836 49276 16892
rect 49276 16836 49332 16892
rect 49332 16836 49336 16892
rect 49272 16832 49336 16836
rect 49352 16892 49416 16896
rect 49352 16836 49356 16892
rect 49356 16836 49412 16892
rect 49412 16836 49416 16892
rect 49352 16832 49416 16836
rect 20216 16348 20280 16352
rect 20216 16292 20220 16348
rect 20220 16292 20276 16348
rect 20276 16292 20280 16348
rect 20216 16288 20280 16292
rect 20296 16348 20360 16352
rect 20296 16292 20300 16348
rect 20300 16292 20356 16348
rect 20356 16292 20360 16348
rect 20296 16288 20360 16292
rect 20376 16348 20440 16352
rect 20376 16292 20380 16348
rect 20380 16292 20436 16348
rect 20436 16292 20440 16348
rect 20376 16288 20440 16292
rect 20456 16348 20520 16352
rect 20456 16292 20460 16348
rect 20460 16292 20516 16348
rect 20516 16292 20520 16348
rect 20456 16288 20520 16292
rect 39480 16348 39544 16352
rect 39480 16292 39484 16348
rect 39484 16292 39540 16348
rect 39540 16292 39544 16348
rect 39480 16288 39544 16292
rect 39560 16348 39624 16352
rect 39560 16292 39564 16348
rect 39564 16292 39620 16348
rect 39620 16292 39624 16348
rect 39560 16288 39624 16292
rect 39640 16348 39704 16352
rect 39640 16292 39644 16348
rect 39644 16292 39700 16348
rect 39700 16292 39704 16348
rect 39640 16288 39704 16292
rect 39720 16348 39784 16352
rect 39720 16292 39724 16348
rect 39724 16292 39780 16348
rect 39780 16292 39784 16348
rect 39720 16288 39784 16292
rect 10584 15804 10648 15808
rect 10584 15748 10588 15804
rect 10588 15748 10644 15804
rect 10644 15748 10648 15804
rect 10584 15744 10648 15748
rect 10664 15804 10728 15808
rect 10664 15748 10668 15804
rect 10668 15748 10724 15804
rect 10724 15748 10728 15804
rect 10664 15744 10728 15748
rect 10744 15804 10808 15808
rect 10744 15748 10748 15804
rect 10748 15748 10804 15804
rect 10804 15748 10808 15804
rect 10744 15744 10808 15748
rect 10824 15804 10888 15808
rect 10824 15748 10828 15804
rect 10828 15748 10884 15804
rect 10884 15748 10888 15804
rect 10824 15744 10888 15748
rect 29848 15804 29912 15808
rect 29848 15748 29852 15804
rect 29852 15748 29908 15804
rect 29908 15748 29912 15804
rect 29848 15744 29912 15748
rect 29928 15804 29992 15808
rect 29928 15748 29932 15804
rect 29932 15748 29988 15804
rect 29988 15748 29992 15804
rect 29928 15744 29992 15748
rect 30008 15804 30072 15808
rect 30008 15748 30012 15804
rect 30012 15748 30068 15804
rect 30068 15748 30072 15804
rect 30008 15744 30072 15748
rect 30088 15804 30152 15808
rect 30088 15748 30092 15804
rect 30092 15748 30148 15804
rect 30148 15748 30152 15804
rect 30088 15744 30152 15748
rect 49112 15804 49176 15808
rect 49112 15748 49116 15804
rect 49116 15748 49172 15804
rect 49172 15748 49176 15804
rect 49112 15744 49176 15748
rect 49192 15804 49256 15808
rect 49192 15748 49196 15804
rect 49196 15748 49252 15804
rect 49252 15748 49256 15804
rect 49192 15744 49256 15748
rect 49272 15804 49336 15808
rect 49272 15748 49276 15804
rect 49276 15748 49332 15804
rect 49332 15748 49336 15804
rect 49272 15744 49336 15748
rect 49352 15804 49416 15808
rect 49352 15748 49356 15804
rect 49356 15748 49412 15804
rect 49412 15748 49416 15804
rect 49352 15744 49416 15748
rect 20216 15260 20280 15264
rect 20216 15204 20220 15260
rect 20220 15204 20276 15260
rect 20276 15204 20280 15260
rect 20216 15200 20280 15204
rect 20296 15260 20360 15264
rect 20296 15204 20300 15260
rect 20300 15204 20356 15260
rect 20356 15204 20360 15260
rect 20296 15200 20360 15204
rect 20376 15260 20440 15264
rect 20376 15204 20380 15260
rect 20380 15204 20436 15260
rect 20436 15204 20440 15260
rect 20376 15200 20440 15204
rect 20456 15260 20520 15264
rect 20456 15204 20460 15260
rect 20460 15204 20516 15260
rect 20516 15204 20520 15260
rect 20456 15200 20520 15204
rect 39480 15260 39544 15264
rect 39480 15204 39484 15260
rect 39484 15204 39540 15260
rect 39540 15204 39544 15260
rect 39480 15200 39544 15204
rect 39560 15260 39624 15264
rect 39560 15204 39564 15260
rect 39564 15204 39620 15260
rect 39620 15204 39624 15260
rect 39560 15200 39624 15204
rect 39640 15260 39704 15264
rect 39640 15204 39644 15260
rect 39644 15204 39700 15260
rect 39700 15204 39704 15260
rect 39640 15200 39704 15204
rect 39720 15260 39784 15264
rect 39720 15204 39724 15260
rect 39724 15204 39780 15260
rect 39780 15204 39784 15260
rect 39720 15200 39784 15204
rect 10584 14716 10648 14720
rect 10584 14660 10588 14716
rect 10588 14660 10644 14716
rect 10644 14660 10648 14716
rect 10584 14656 10648 14660
rect 10664 14716 10728 14720
rect 10664 14660 10668 14716
rect 10668 14660 10724 14716
rect 10724 14660 10728 14716
rect 10664 14656 10728 14660
rect 10744 14716 10808 14720
rect 10744 14660 10748 14716
rect 10748 14660 10804 14716
rect 10804 14660 10808 14716
rect 10744 14656 10808 14660
rect 10824 14716 10888 14720
rect 10824 14660 10828 14716
rect 10828 14660 10884 14716
rect 10884 14660 10888 14716
rect 10824 14656 10888 14660
rect 29848 14716 29912 14720
rect 29848 14660 29852 14716
rect 29852 14660 29908 14716
rect 29908 14660 29912 14716
rect 29848 14656 29912 14660
rect 29928 14716 29992 14720
rect 29928 14660 29932 14716
rect 29932 14660 29988 14716
rect 29988 14660 29992 14716
rect 29928 14656 29992 14660
rect 30008 14716 30072 14720
rect 30008 14660 30012 14716
rect 30012 14660 30068 14716
rect 30068 14660 30072 14716
rect 30008 14656 30072 14660
rect 30088 14716 30152 14720
rect 30088 14660 30092 14716
rect 30092 14660 30148 14716
rect 30148 14660 30152 14716
rect 30088 14656 30152 14660
rect 49112 14716 49176 14720
rect 49112 14660 49116 14716
rect 49116 14660 49172 14716
rect 49172 14660 49176 14716
rect 49112 14656 49176 14660
rect 49192 14716 49256 14720
rect 49192 14660 49196 14716
rect 49196 14660 49252 14716
rect 49252 14660 49256 14716
rect 49192 14656 49256 14660
rect 49272 14716 49336 14720
rect 49272 14660 49276 14716
rect 49276 14660 49332 14716
rect 49332 14660 49336 14716
rect 49272 14656 49336 14660
rect 49352 14716 49416 14720
rect 49352 14660 49356 14716
rect 49356 14660 49412 14716
rect 49412 14660 49416 14716
rect 49352 14656 49416 14660
rect 20216 14172 20280 14176
rect 20216 14116 20220 14172
rect 20220 14116 20276 14172
rect 20276 14116 20280 14172
rect 20216 14112 20280 14116
rect 20296 14172 20360 14176
rect 20296 14116 20300 14172
rect 20300 14116 20356 14172
rect 20356 14116 20360 14172
rect 20296 14112 20360 14116
rect 20376 14172 20440 14176
rect 20376 14116 20380 14172
rect 20380 14116 20436 14172
rect 20436 14116 20440 14172
rect 20376 14112 20440 14116
rect 20456 14172 20520 14176
rect 20456 14116 20460 14172
rect 20460 14116 20516 14172
rect 20516 14116 20520 14172
rect 20456 14112 20520 14116
rect 39480 14172 39544 14176
rect 39480 14116 39484 14172
rect 39484 14116 39540 14172
rect 39540 14116 39544 14172
rect 39480 14112 39544 14116
rect 39560 14172 39624 14176
rect 39560 14116 39564 14172
rect 39564 14116 39620 14172
rect 39620 14116 39624 14172
rect 39560 14112 39624 14116
rect 39640 14172 39704 14176
rect 39640 14116 39644 14172
rect 39644 14116 39700 14172
rect 39700 14116 39704 14172
rect 39640 14112 39704 14116
rect 39720 14172 39784 14176
rect 39720 14116 39724 14172
rect 39724 14116 39780 14172
rect 39780 14116 39784 14172
rect 39720 14112 39784 14116
rect 10584 13628 10648 13632
rect 10584 13572 10588 13628
rect 10588 13572 10644 13628
rect 10644 13572 10648 13628
rect 10584 13568 10648 13572
rect 10664 13628 10728 13632
rect 10664 13572 10668 13628
rect 10668 13572 10724 13628
rect 10724 13572 10728 13628
rect 10664 13568 10728 13572
rect 10744 13628 10808 13632
rect 10744 13572 10748 13628
rect 10748 13572 10804 13628
rect 10804 13572 10808 13628
rect 10744 13568 10808 13572
rect 10824 13628 10888 13632
rect 10824 13572 10828 13628
rect 10828 13572 10884 13628
rect 10884 13572 10888 13628
rect 10824 13568 10888 13572
rect 29848 13628 29912 13632
rect 29848 13572 29852 13628
rect 29852 13572 29908 13628
rect 29908 13572 29912 13628
rect 29848 13568 29912 13572
rect 29928 13628 29992 13632
rect 29928 13572 29932 13628
rect 29932 13572 29988 13628
rect 29988 13572 29992 13628
rect 29928 13568 29992 13572
rect 30008 13628 30072 13632
rect 30008 13572 30012 13628
rect 30012 13572 30068 13628
rect 30068 13572 30072 13628
rect 30008 13568 30072 13572
rect 30088 13628 30152 13632
rect 30088 13572 30092 13628
rect 30092 13572 30148 13628
rect 30148 13572 30152 13628
rect 30088 13568 30152 13572
rect 49112 13628 49176 13632
rect 49112 13572 49116 13628
rect 49116 13572 49172 13628
rect 49172 13572 49176 13628
rect 49112 13568 49176 13572
rect 49192 13628 49256 13632
rect 49192 13572 49196 13628
rect 49196 13572 49252 13628
rect 49252 13572 49256 13628
rect 49192 13568 49256 13572
rect 49272 13628 49336 13632
rect 49272 13572 49276 13628
rect 49276 13572 49332 13628
rect 49332 13572 49336 13628
rect 49272 13568 49336 13572
rect 49352 13628 49416 13632
rect 49352 13572 49356 13628
rect 49356 13572 49412 13628
rect 49412 13572 49416 13628
rect 49352 13568 49416 13572
rect 20216 13084 20280 13088
rect 20216 13028 20220 13084
rect 20220 13028 20276 13084
rect 20276 13028 20280 13084
rect 20216 13024 20280 13028
rect 20296 13084 20360 13088
rect 20296 13028 20300 13084
rect 20300 13028 20356 13084
rect 20356 13028 20360 13084
rect 20296 13024 20360 13028
rect 20376 13084 20440 13088
rect 20376 13028 20380 13084
rect 20380 13028 20436 13084
rect 20436 13028 20440 13084
rect 20376 13024 20440 13028
rect 20456 13084 20520 13088
rect 20456 13028 20460 13084
rect 20460 13028 20516 13084
rect 20516 13028 20520 13084
rect 20456 13024 20520 13028
rect 39480 13084 39544 13088
rect 39480 13028 39484 13084
rect 39484 13028 39540 13084
rect 39540 13028 39544 13084
rect 39480 13024 39544 13028
rect 39560 13084 39624 13088
rect 39560 13028 39564 13084
rect 39564 13028 39620 13084
rect 39620 13028 39624 13084
rect 39560 13024 39624 13028
rect 39640 13084 39704 13088
rect 39640 13028 39644 13084
rect 39644 13028 39700 13084
rect 39700 13028 39704 13084
rect 39640 13024 39704 13028
rect 39720 13084 39784 13088
rect 39720 13028 39724 13084
rect 39724 13028 39780 13084
rect 39780 13028 39784 13084
rect 39720 13024 39784 13028
rect 10584 12540 10648 12544
rect 10584 12484 10588 12540
rect 10588 12484 10644 12540
rect 10644 12484 10648 12540
rect 10584 12480 10648 12484
rect 10664 12540 10728 12544
rect 10664 12484 10668 12540
rect 10668 12484 10724 12540
rect 10724 12484 10728 12540
rect 10664 12480 10728 12484
rect 10744 12540 10808 12544
rect 10744 12484 10748 12540
rect 10748 12484 10804 12540
rect 10804 12484 10808 12540
rect 10744 12480 10808 12484
rect 10824 12540 10888 12544
rect 10824 12484 10828 12540
rect 10828 12484 10884 12540
rect 10884 12484 10888 12540
rect 10824 12480 10888 12484
rect 29848 12540 29912 12544
rect 29848 12484 29852 12540
rect 29852 12484 29908 12540
rect 29908 12484 29912 12540
rect 29848 12480 29912 12484
rect 29928 12540 29992 12544
rect 29928 12484 29932 12540
rect 29932 12484 29988 12540
rect 29988 12484 29992 12540
rect 29928 12480 29992 12484
rect 30008 12540 30072 12544
rect 30008 12484 30012 12540
rect 30012 12484 30068 12540
rect 30068 12484 30072 12540
rect 30008 12480 30072 12484
rect 30088 12540 30152 12544
rect 30088 12484 30092 12540
rect 30092 12484 30148 12540
rect 30148 12484 30152 12540
rect 30088 12480 30152 12484
rect 49112 12540 49176 12544
rect 49112 12484 49116 12540
rect 49116 12484 49172 12540
rect 49172 12484 49176 12540
rect 49112 12480 49176 12484
rect 49192 12540 49256 12544
rect 49192 12484 49196 12540
rect 49196 12484 49252 12540
rect 49252 12484 49256 12540
rect 49192 12480 49256 12484
rect 49272 12540 49336 12544
rect 49272 12484 49276 12540
rect 49276 12484 49332 12540
rect 49332 12484 49336 12540
rect 49272 12480 49336 12484
rect 49352 12540 49416 12544
rect 49352 12484 49356 12540
rect 49356 12484 49412 12540
rect 49412 12484 49416 12540
rect 49352 12480 49416 12484
rect 20216 11996 20280 12000
rect 20216 11940 20220 11996
rect 20220 11940 20276 11996
rect 20276 11940 20280 11996
rect 20216 11936 20280 11940
rect 20296 11996 20360 12000
rect 20296 11940 20300 11996
rect 20300 11940 20356 11996
rect 20356 11940 20360 11996
rect 20296 11936 20360 11940
rect 20376 11996 20440 12000
rect 20376 11940 20380 11996
rect 20380 11940 20436 11996
rect 20436 11940 20440 11996
rect 20376 11936 20440 11940
rect 20456 11996 20520 12000
rect 20456 11940 20460 11996
rect 20460 11940 20516 11996
rect 20516 11940 20520 11996
rect 20456 11936 20520 11940
rect 39480 11996 39544 12000
rect 39480 11940 39484 11996
rect 39484 11940 39540 11996
rect 39540 11940 39544 11996
rect 39480 11936 39544 11940
rect 39560 11996 39624 12000
rect 39560 11940 39564 11996
rect 39564 11940 39620 11996
rect 39620 11940 39624 11996
rect 39560 11936 39624 11940
rect 39640 11996 39704 12000
rect 39640 11940 39644 11996
rect 39644 11940 39700 11996
rect 39700 11940 39704 11996
rect 39640 11936 39704 11940
rect 39720 11996 39784 12000
rect 39720 11940 39724 11996
rect 39724 11940 39780 11996
rect 39780 11940 39784 11996
rect 39720 11936 39784 11940
rect 10584 11452 10648 11456
rect 10584 11396 10588 11452
rect 10588 11396 10644 11452
rect 10644 11396 10648 11452
rect 10584 11392 10648 11396
rect 10664 11452 10728 11456
rect 10664 11396 10668 11452
rect 10668 11396 10724 11452
rect 10724 11396 10728 11452
rect 10664 11392 10728 11396
rect 10744 11452 10808 11456
rect 10744 11396 10748 11452
rect 10748 11396 10804 11452
rect 10804 11396 10808 11452
rect 10744 11392 10808 11396
rect 10824 11452 10888 11456
rect 10824 11396 10828 11452
rect 10828 11396 10884 11452
rect 10884 11396 10888 11452
rect 10824 11392 10888 11396
rect 29848 11452 29912 11456
rect 29848 11396 29852 11452
rect 29852 11396 29908 11452
rect 29908 11396 29912 11452
rect 29848 11392 29912 11396
rect 29928 11452 29992 11456
rect 29928 11396 29932 11452
rect 29932 11396 29988 11452
rect 29988 11396 29992 11452
rect 29928 11392 29992 11396
rect 30008 11452 30072 11456
rect 30008 11396 30012 11452
rect 30012 11396 30068 11452
rect 30068 11396 30072 11452
rect 30008 11392 30072 11396
rect 30088 11452 30152 11456
rect 30088 11396 30092 11452
rect 30092 11396 30148 11452
rect 30148 11396 30152 11452
rect 30088 11392 30152 11396
rect 49112 11452 49176 11456
rect 49112 11396 49116 11452
rect 49116 11396 49172 11452
rect 49172 11396 49176 11452
rect 49112 11392 49176 11396
rect 49192 11452 49256 11456
rect 49192 11396 49196 11452
rect 49196 11396 49252 11452
rect 49252 11396 49256 11452
rect 49192 11392 49256 11396
rect 49272 11452 49336 11456
rect 49272 11396 49276 11452
rect 49276 11396 49332 11452
rect 49332 11396 49336 11452
rect 49272 11392 49336 11396
rect 49352 11452 49416 11456
rect 49352 11396 49356 11452
rect 49356 11396 49412 11452
rect 49412 11396 49416 11452
rect 49352 11392 49416 11396
rect 20216 10908 20280 10912
rect 20216 10852 20220 10908
rect 20220 10852 20276 10908
rect 20276 10852 20280 10908
rect 20216 10848 20280 10852
rect 20296 10908 20360 10912
rect 20296 10852 20300 10908
rect 20300 10852 20356 10908
rect 20356 10852 20360 10908
rect 20296 10848 20360 10852
rect 20376 10908 20440 10912
rect 20376 10852 20380 10908
rect 20380 10852 20436 10908
rect 20436 10852 20440 10908
rect 20376 10848 20440 10852
rect 20456 10908 20520 10912
rect 20456 10852 20460 10908
rect 20460 10852 20516 10908
rect 20516 10852 20520 10908
rect 20456 10848 20520 10852
rect 39480 10908 39544 10912
rect 39480 10852 39484 10908
rect 39484 10852 39540 10908
rect 39540 10852 39544 10908
rect 39480 10848 39544 10852
rect 39560 10908 39624 10912
rect 39560 10852 39564 10908
rect 39564 10852 39620 10908
rect 39620 10852 39624 10908
rect 39560 10848 39624 10852
rect 39640 10908 39704 10912
rect 39640 10852 39644 10908
rect 39644 10852 39700 10908
rect 39700 10852 39704 10908
rect 39640 10848 39704 10852
rect 39720 10908 39784 10912
rect 39720 10852 39724 10908
rect 39724 10852 39780 10908
rect 39780 10852 39784 10908
rect 39720 10848 39784 10852
rect 10584 10364 10648 10368
rect 10584 10308 10588 10364
rect 10588 10308 10644 10364
rect 10644 10308 10648 10364
rect 10584 10304 10648 10308
rect 10664 10364 10728 10368
rect 10664 10308 10668 10364
rect 10668 10308 10724 10364
rect 10724 10308 10728 10364
rect 10664 10304 10728 10308
rect 10744 10364 10808 10368
rect 10744 10308 10748 10364
rect 10748 10308 10804 10364
rect 10804 10308 10808 10364
rect 10744 10304 10808 10308
rect 10824 10364 10888 10368
rect 10824 10308 10828 10364
rect 10828 10308 10884 10364
rect 10884 10308 10888 10364
rect 10824 10304 10888 10308
rect 29848 10364 29912 10368
rect 29848 10308 29852 10364
rect 29852 10308 29908 10364
rect 29908 10308 29912 10364
rect 29848 10304 29912 10308
rect 29928 10364 29992 10368
rect 29928 10308 29932 10364
rect 29932 10308 29988 10364
rect 29988 10308 29992 10364
rect 29928 10304 29992 10308
rect 30008 10364 30072 10368
rect 30008 10308 30012 10364
rect 30012 10308 30068 10364
rect 30068 10308 30072 10364
rect 30008 10304 30072 10308
rect 30088 10364 30152 10368
rect 30088 10308 30092 10364
rect 30092 10308 30148 10364
rect 30148 10308 30152 10364
rect 30088 10304 30152 10308
rect 49112 10364 49176 10368
rect 49112 10308 49116 10364
rect 49116 10308 49172 10364
rect 49172 10308 49176 10364
rect 49112 10304 49176 10308
rect 49192 10364 49256 10368
rect 49192 10308 49196 10364
rect 49196 10308 49252 10364
rect 49252 10308 49256 10364
rect 49192 10304 49256 10308
rect 49272 10364 49336 10368
rect 49272 10308 49276 10364
rect 49276 10308 49332 10364
rect 49332 10308 49336 10364
rect 49272 10304 49336 10308
rect 49352 10364 49416 10368
rect 49352 10308 49356 10364
rect 49356 10308 49412 10364
rect 49412 10308 49416 10364
rect 49352 10304 49416 10308
rect 20216 9820 20280 9824
rect 20216 9764 20220 9820
rect 20220 9764 20276 9820
rect 20276 9764 20280 9820
rect 20216 9760 20280 9764
rect 20296 9820 20360 9824
rect 20296 9764 20300 9820
rect 20300 9764 20356 9820
rect 20356 9764 20360 9820
rect 20296 9760 20360 9764
rect 20376 9820 20440 9824
rect 20376 9764 20380 9820
rect 20380 9764 20436 9820
rect 20436 9764 20440 9820
rect 20376 9760 20440 9764
rect 20456 9820 20520 9824
rect 20456 9764 20460 9820
rect 20460 9764 20516 9820
rect 20516 9764 20520 9820
rect 20456 9760 20520 9764
rect 39480 9820 39544 9824
rect 39480 9764 39484 9820
rect 39484 9764 39540 9820
rect 39540 9764 39544 9820
rect 39480 9760 39544 9764
rect 39560 9820 39624 9824
rect 39560 9764 39564 9820
rect 39564 9764 39620 9820
rect 39620 9764 39624 9820
rect 39560 9760 39624 9764
rect 39640 9820 39704 9824
rect 39640 9764 39644 9820
rect 39644 9764 39700 9820
rect 39700 9764 39704 9820
rect 39640 9760 39704 9764
rect 39720 9820 39784 9824
rect 39720 9764 39724 9820
rect 39724 9764 39780 9820
rect 39780 9764 39784 9820
rect 39720 9760 39784 9764
rect 10584 9276 10648 9280
rect 10584 9220 10588 9276
rect 10588 9220 10644 9276
rect 10644 9220 10648 9276
rect 10584 9216 10648 9220
rect 10664 9276 10728 9280
rect 10664 9220 10668 9276
rect 10668 9220 10724 9276
rect 10724 9220 10728 9276
rect 10664 9216 10728 9220
rect 10744 9276 10808 9280
rect 10744 9220 10748 9276
rect 10748 9220 10804 9276
rect 10804 9220 10808 9276
rect 10744 9216 10808 9220
rect 10824 9276 10888 9280
rect 10824 9220 10828 9276
rect 10828 9220 10884 9276
rect 10884 9220 10888 9276
rect 10824 9216 10888 9220
rect 29848 9276 29912 9280
rect 29848 9220 29852 9276
rect 29852 9220 29908 9276
rect 29908 9220 29912 9276
rect 29848 9216 29912 9220
rect 29928 9276 29992 9280
rect 29928 9220 29932 9276
rect 29932 9220 29988 9276
rect 29988 9220 29992 9276
rect 29928 9216 29992 9220
rect 30008 9276 30072 9280
rect 30008 9220 30012 9276
rect 30012 9220 30068 9276
rect 30068 9220 30072 9276
rect 30008 9216 30072 9220
rect 30088 9276 30152 9280
rect 30088 9220 30092 9276
rect 30092 9220 30148 9276
rect 30148 9220 30152 9276
rect 30088 9216 30152 9220
rect 49112 9276 49176 9280
rect 49112 9220 49116 9276
rect 49116 9220 49172 9276
rect 49172 9220 49176 9276
rect 49112 9216 49176 9220
rect 49192 9276 49256 9280
rect 49192 9220 49196 9276
rect 49196 9220 49252 9276
rect 49252 9220 49256 9276
rect 49192 9216 49256 9220
rect 49272 9276 49336 9280
rect 49272 9220 49276 9276
rect 49276 9220 49332 9276
rect 49332 9220 49336 9276
rect 49272 9216 49336 9220
rect 49352 9276 49416 9280
rect 49352 9220 49356 9276
rect 49356 9220 49412 9276
rect 49412 9220 49416 9276
rect 49352 9216 49416 9220
rect 20216 8732 20280 8736
rect 20216 8676 20220 8732
rect 20220 8676 20276 8732
rect 20276 8676 20280 8732
rect 20216 8672 20280 8676
rect 20296 8732 20360 8736
rect 20296 8676 20300 8732
rect 20300 8676 20356 8732
rect 20356 8676 20360 8732
rect 20296 8672 20360 8676
rect 20376 8732 20440 8736
rect 20376 8676 20380 8732
rect 20380 8676 20436 8732
rect 20436 8676 20440 8732
rect 20376 8672 20440 8676
rect 20456 8732 20520 8736
rect 20456 8676 20460 8732
rect 20460 8676 20516 8732
rect 20516 8676 20520 8732
rect 20456 8672 20520 8676
rect 39480 8732 39544 8736
rect 39480 8676 39484 8732
rect 39484 8676 39540 8732
rect 39540 8676 39544 8732
rect 39480 8672 39544 8676
rect 39560 8732 39624 8736
rect 39560 8676 39564 8732
rect 39564 8676 39620 8732
rect 39620 8676 39624 8732
rect 39560 8672 39624 8676
rect 39640 8732 39704 8736
rect 39640 8676 39644 8732
rect 39644 8676 39700 8732
rect 39700 8676 39704 8732
rect 39640 8672 39704 8676
rect 39720 8732 39784 8736
rect 39720 8676 39724 8732
rect 39724 8676 39780 8732
rect 39780 8676 39784 8732
rect 39720 8672 39784 8676
rect 10584 8188 10648 8192
rect 10584 8132 10588 8188
rect 10588 8132 10644 8188
rect 10644 8132 10648 8188
rect 10584 8128 10648 8132
rect 10664 8188 10728 8192
rect 10664 8132 10668 8188
rect 10668 8132 10724 8188
rect 10724 8132 10728 8188
rect 10664 8128 10728 8132
rect 10744 8188 10808 8192
rect 10744 8132 10748 8188
rect 10748 8132 10804 8188
rect 10804 8132 10808 8188
rect 10744 8128 10808 8132
rect 10824 8188 10888 8192
rect 10824 8132 10828 8188
rect 10828 8132 10884 8188
rect 10884 8132 10888 8188
rect 10824 8128 10888 8132
rect 29848 8188 29912 8192
rect 29848 8132 29852 8188
rect 29852 8132 29908 8188
rect 29908 8132 29912 8188
rect 29848 8128 29912 8132
rect 29928 8188 29992 8192
rect 29928 8132 29932 8188
rect 29932 8132 29988 8188
rect 29988 8132 29992 8188
rect 29928 8128 29992 8132
rect 30008 8188 30072 8192
rect 30008 8132 30012 8188
rect 30012 8132 30068 8188
rect 30068 8132 30072 8188
rect 30008 8128 30072 8132
rect 30088 8188 30152 8192
rect 30088 8132 30092 8188
rect 30092 8132 30148 8188
rect 30148 8132 30152 8188
rect 30088 8128 30152 8132
rect 49112 8188 49176 8192
rect 49112 8132 49116 8188
rect 49116 8132 49172 8188
rect 49172 8132 49176 8188
rect 49112 8128 49176 8132
rect 49192 8188 49256 8192
rect 49192 8132 49196 8188
rect 49196 8132 49252 8188
rect 49252 8132 49256 8188
rect 49192 8128 49256 8132
rect 49272 8188 49336 8192
rect 49272 8132 49276 8188
rect 49276 8132 49332 8188
rect 49332 8132 49336 8188
rect 49272 8128 49336 8132
rect 49352 8188 49416 8192
rect 49352 8132 49356 8188
rect 49356 8132 49412 8188
rect 49412 8132 49416 8188
rect 49352 8128 49416 8132
rect 20216 7644 20280 7648
rect 20216 7588 20220 7644
rect 20220 7588 20276 7644
rect 20276 7588 20280 7644
rect 20216 7584 20280 7588
rect 20296 7644 20360 7648
rect 20296 7588 20300 7644
rect 20300 7588 20356 7644
rect 20356 7588 20360 7644
rect 20296 7584 20360 7588
rect 20376 7644 20440 7648
rect 20376 7588 20380 7644
rect 20380 7588 20436 7644
rect 20436 7588 20440 7644
rect 20376 7584 20440 7588
rect 20456 7644 20520 7648
rect 20456 7588 20460 7644
rect 20460 7588 20516 7644
rect 20516 7588 20520 7644
rect 20456 7584 20520 7588
rect 39480 7644 39544 7648
rect 39480 7588 39484 7644
rect 39484 7588 39540 7644
rect 39540 7588 39544 7644
rect 39480 7584 39544 7588
rect 39560 7644 39624 7648
rect 39560 7588 39564 7644
rect 39564 7588 39620 7644
rect 39620 7588 39624 7644
rect 39560 7584 39624 7588
rect 39640 7644 39704 7648
rect 39640 7588 39644 7644
rect 39644 7588 39700 7644
rect 39700 7588 39704 7644
rect 39640 7584 39704 7588
rect 39720 7644 39784 7648
rect 39720 7588 39724 7644
rect 39724 7588 39780 7644
rect 39780 7588 39784 7644
rect 39720 7584 39784 7588
rect 10584 7100 10648 7104
rect 10584 7044 10588 7100
rect 10588 7044 10644 7100
rect 10644 7044 10648 7100
rect 10584 7040 10648 7044
rect 10664 7100 10728 7104
rect 10664 7044 10668 7100
rect 10668 7044 10724 7100
rect 10724 7044 10728 7100
rect 10664 7040 10728 7044
rect 10744 7100 10808 7104
rect 10744 7044 10748 7100
rect 10748 7044 10804 7100
rect 10804 7044 10808 7100
rect 10744 7040 10808 7044
rect 10824 7100 10888 7104
rect 10824 7044 10828 7100
rect 10828 7044 10884 7100
rect 10884 7044 10888 7100
rect 10824 7040 10888 7044
rect 29848 7100 29912 7104
rect 29848 7044 29852 7100
rect 29852 7044 29908 7100
rect 29908 7044 29912 7100
rect 29848 7040 29912 7044
rect 29928 7100 29992 7104
rect 29928 7044 29932 7100
rect 29932 7044 29988 7100
rect 29988 7044 29992 7100
rect 29928 7040 29992 7044
rect 30008 7100 30072 7104
rect 30008 7044 30012 7100
rect 30012 7044 30068 7100
rect 30068 7044 30072 7100
rect 30008 7040 30072 7044
rect 30088 7100 30152 7104
rect 30088 7044 30092 7100
rect 30092 7044 30148 7100
rect 30148 7044 30152 7100
rect 30088 7040 30152 7044
rect 49112 7100 49176 7104
rect 49112 7044 49116 7100
rect 49116 7044 49172 7100
rect 49172 7044 49176 7100
rect 49112 7040 49176 7044
rect 49192 7100 49256 7104
rect 49192 7044 49196 7100
rect 49196 7044 49252 7100
rect 49252 7044 49256 7100
rect 49192 7040 49256 7044
rect 49272 7100 49336 7104
rect 49272 7044 49276 7100
rect 49276 7044 49332 7100
rect 49332 7044 49336 7100
rect 49272 7040 49336 7044
rect 49352 7100 49416 7104
rect 49352 7044 49356 7100
rect 49356 7044 49412 7100
rect 49412 7044 49416 7100
rect 49352 7040 49416 7044
rect 20216 6556 20280 6560
rect 20216 6500 20220 6556
rect 20220 6500 20276 6556
rect 20276 6500 20280 6556
rect 20216 6496 20280 6500
rect 20296 6556 20360 6560
rect 20296 6500 20300 6556
rect 20300 6500 20356 6556
rect 20356 6500 20360 6556
rect 20296 6496 20360 6500
rect 20376 6556 20440 6560
rect 20376 6500 20380 6556
rect 20380 6500 20436 6556
rect 20436 6500 20440 6556
rect 20376 6496 20440 6500
rect 20456 6556 20520 6560
rect 20456 6500 20460 6556
rect 20460 6500 20516 6556
rect 20516 6500 20520 6556
rect 20456 6496 20520 6500
rect 39480 6556 39544 6560
rect 39480 6500 39484 6556
rect 39484 6500 39540 6556
rect 39540 6500 39544 6556
rect 39480 6496 39544 6500
rect 39560 6556 39624 6560
rect 39560 6500 39564 6556
rect 39564 6500 39620 6556
rect 39620 6500 39624 6556
rect 39560 6496 39624 6500
rect 39640 6556 39704 6560
rect 39640 6500 39644 6556
rect 39644 6500 39700 6556
rect 39700 6500 39704 6556
rect 39640 6496 39704 6500
rect 39720 6556 39784 6560
rect 39720 6500 39724 6556
rect 39724 6500 39780 6556
rect 39780 6500 39784 6556
rect 39720 6496 39784 6500
rect 10584 6012 10648 6016
rect 10584 5956 10588 6012
rect 10588 5956 10644 6012
rect 10644 5956 10648 6012
rect 10584 5952 10648 5956
rect 10664 6012 10728 6016
rect 10664 5956 10668 6012
rect 10668 5956 10724 6012
rect 10724 5956 10728 6012
rect 10664 5952 10728 5956
rect 10744 6012 10808 6016
rect 10744 5956 10748 6012
rect 10748 5956 10804 6012
rect 10804 5956 10808 6012
rect 10744 5952 10808 5956
rect 10824 6012 10888 6016
rect 10824 5956 10828 6012
rect 10828 5956 10884 6012
rect 10884 5956 10888 6012
rect 10824 5952 10888 5956
rect 29848 6012 29912 6016
rect 29848 5956 29852 6012
rect 29852 5956 29908 6012
rect 29908 5956 29912 6012
rect 29848 5952 29912 5956
rect 29928 6012 29992 6016
rect 29928 5956 29932 6012
rect 29932 5956 29988 6012
rect 29988 5956 29992 6012
rect 29928 5952 29992 5956
rect 30008 6012 30072 6016
rect 30008 5956 30012 6012
rect 30012 5956 30068 6012
rect 30068 5956 30072 6012
rect 30008 5952 30072 5956
rect 30088 6012 30152 6016
rect 30088 5956 30092 6012
rect 30092 5956 30148 6012
rect 30148 5956 30152 6012
rect 30088 5952 30152 5956
rect 49112 6012 49176 6016
rect 49112 5956 49116 6012
rect 49116 5956 49172 6012
rect 49172 5956 49176 6012
rect 49112 5952 49176 5956
rect 49192 6012 49256 6016
rect 49192 5956 49196 6012
rect 49196 5956 49252 6012
rect 49252 5956 49256 6012
rect 49192 5952 49256 5956
rect 49272 6012 49336 6016
rect 49272 5956 49276 6012
rect 49276 5956 49332 6012
rect 49332 5956 49336 6012
rect 49272 5952 49336 5956
rect 49352 6012 49416 6016
rect 49352 5956 49356 6012
rect 49356 5956 49412 6012
rect 49412 5956 49416 6012
rect 49352 5952 49416 5956
rect 20216 5468 20280 5472
rect 20216 5412 20220 5468
rect 20220 5412 20276 5468
rect 20276 5412 20280 5468
rect 20216 5408 20280 5412
rect 20296 5468 20360 5472
rect 20296 5412 20300 5468
rect 20300 5412 20356 5468
rect 20356 5412 20360 5468
rect 20296 5408 20360 5412
rect 20376 5468 20440 5472
rect 20376 5412 20380 5468
rect 20380 5412 20436 5468
rect 20436 5412 20440 5468
rect 20376 5408 20440 5412
rect 20456 5468 20520 5472
rect 20456 5412 20460 5468
rect 20460 5412 20516 5468
rect 20516 5412 20520 5468
rect 20456 5408 20520 5412
rect 39480 5468 39544 5472
rect 39480 5412 39484 5468
rect 39484 5412 39540 5468
rect 39540 5412 39544 5468
rect 39480 5408 39544 5412
rect 39560 5468 39624 5472
rect 39560 5412 39564 5468
rect 39564 5412 39620 5468
rect 39620 5412 39624 5468
rect 39560 5408 39624 5412
rect 39640 5468 39704 5472
rect 39640 5412 39644 5468
rect 39644 5412 39700 5468
rect 39700 5412 39704 5468
rect 39640 5408 39704 5412
rect 39720 5468 39784 5472
rect 39720 5412 39724 5468
rect 39724 5412 39780 5468
rect 39780 5412 39784 5468
rect 39720 5408 39784 5412
rect 10584 4924 10648 4928
rect 10584 4868 10588 4924
rect 10588 4868 10644 4924
rect 10644 4868 10648 4924
rect 10584 4864 10648 4868
rect 10664 4924 10728 4928
rect 10664 4868 10668 4924
rect 10668 4868 10724 4924
rect 10724 4868 10728 4924
rect 10664 4864 10728 4868
rect 10744 4924 10808 4928
rect 10744 4868 10748 4924
rect 10748 4868 10804 4924
rect 10804 4868 10808 4924
rect 10744 4864 10808 4868
rect 10824 4924 10888 4928
rect 10824 4868 10828 4924
rect 10828 4868 10884 4924
rect 10884 4868 10888 4924
rect 10824 4864 10888 4868
rect 29848 4924 29912 4928
rect 29848 4868 29852 4924
rect 29852 4868 29908 4924
rect 29908 4868 29912 4924
rect 29848 4864 29912 4868
rect 29928 4924 29992 4928
rect 29928 4868 29932 4924
rect 29932 4868 29988 4924
rect 29988 4868 29992 4924
rect 29928 4864 29992 4868
rect 30008 4924 30072 4928
rect 30008 4868 30012 4924
rect 30012 4868 30068 4924
rect 30068 4868 30072 4924
rect 30008 4864 30072 4868
rect 30088 4924 30152 4928
rect 30088 4868 30092 4924
rect 30092 4868 30148 4924
rect 30148 4868 30152 4924
rect 30088 4864 30152 4868
rect 49112 4924 49176 4928
rect 49112 4868 49116 4924
rect 49116 4868 49172 4924
rect 49172 4868 49176 4924
rect 49112 4864 49176 4868
rect 49192 4924 49256 4928
rect 49192 4868 49196 4924
rect 49196 4868 49252 4924
rect 49252 4868 49256 4924
rect 49192 4864 49256 4868
rect 49272 4924 49336 4928
rect 49272 4868 49276 4924
rect 49276 4868 49332 4924
rect 49332 4868 49336 4924
rect 49272 4864 49336 4868
rect 49352 4924 49416 4928
rect 49352 4868 49356 4924
rect 49356 4868 49412 4924
rect 49412 4868 49416 4924
rect 49352 4864 49416 4868
rect 20216 4380 20280 4384
rect 20216 4324 20220 4380
rect 20220 4324 20276 4380
rect 20276 4324 20280 4380
rect 20216 4320 20280 4324
rect 20296 4380 20360 4384
rect 20296 4324 20300 4380
rect 20300 4324 20356 4380
rect 20356 4324 20360 4380
rect 20296 4320 20360 4324
rect 20376 4380 20440 4384
rect 20376 4324 20380 4380
rect 20380 4324 20436 4380
rect 20436 4324 20440 4380
rect 20376 4320 20440 4324
rect 20456 4380 20520 4384
rect 20456 4324 20460 4380
rect 20460 4324 20516 4380
rect 20516 4324 20520 4380
rect 20456 4320 20520 4324
rect 39480 4380 39544 4384
rect 39480 4324 39484 4380
rect 39484 4324 39540 4380
rect 39540 4324 39544 4380
rect 39480 4320 39544 4324
rect 39560 4380 39624 4384
rect 39560 4324 39564 4380
rect 39564 4324 39620 4380
rect 39620 4324 39624 4380
rect 39560 4320 39624 4324
rect 39640 4380 39704 4384
rect 39640 4324 39644 4380
rect 39644 4324 39700 4380
rect 39700 4324 39704 4380
rect 39640 4320 39704 4324
rect 39720 4380 39784 4384
rect 39720 4324 39724 4380
rect 39724 4324 39780 4380
rect 39780 4324 39784 4380
rect 39720 4320 39784 4324
rect 10584 3836 10648 3840
rect 10584 3780 10588 3836
rect 10588 3780 10644 3836
rect 10644 3780 10648 3836
rect 10584 3776 10648 3780
rect 10664 3836 10728 3840
rect 10664 3780 10668 3836
rect 10668 3780 10724 3836
rect 10724 3780 10728 3836
rect 10664 3776 10728 3780
rect 10744 3836 10808 3840
rect 10744 3780 10748 3836
rect 10748 3780 10804 3836
rect 10804 3780 10808 3836
rect 10744 3776 10808 3780
rect 10824 3836 10888 3840
rect 10824 3780 10828 3836
rect 10828 3780 10884 3836
rect 10884 3780 10888 3836
rect 10824 3776 10888 3780
rect 29848 3836 29912 3840
rect 29848 3780 29852 3836
rect 29852 3780 29908 3836
rect 29908 3780 29912 3836
rect 29848 3776 29912 3780
rect 29928 3836 29992 3840
rect 29928 3780 29932 3836
rect 29932 3780 29988 3836
rect 29988 3780 29992 3836
rect 29928 3776 29992 3780
rect 30008 3836 30072 3840
rect 30008 3780 30012 3836
rect 30012 3780 30068 3836
rect 30068 3780 30072 3836
rect 30008 3776 30072 3780
rect 30088 3836 30152 3840
rect 30088 3780 30092 3836
rect 30092 3780 30148 3836
rect 30148 3780 30152 3836
rect 30088 3776 30152 3780
rect 49112 3836 49176 3840
rect 49112 3780 49116 3836
rect 49116 3780 49172 3836
rect 49172 3780 49176 3836
rect 49112 3776 49176 3780
rect 49192 3836 49256 3840
rect 49192 3780 49196 3836
rect 49196 3780 49252 3836
rect 49252 3780 49256 3836
rect 49192 3776 49256 3780
rect 49272 3836 49336 3840
rect 49272 3780 49276 3836
rect 49276 3780 49332 3836
rect 49332 3780 49336 3836
rect 49272 3776 49336 3780
rect 49352 3836 49416 3840
rect 49352 3780 49356 3836
rect 49356 3780 49412 3836
rect 49412 3780 49416 3836
rect 49352 3776 49416 3780
rect 20216 3292 20280 3296
rect 20216 3236 20220 3292
rect 20220 3236 20276 3292
rect 20276 3236 20280 3292
rect 20216 3232 20280 3236
rect 20296 3292 20360 3296
rect 20296 3236 20300 3292
rect 20300 3236 20356 3292
rect 20356 3236 20360 3292
rect 20296 3232 20360 3236
rect 20376 3292 20440 3296
rect 20376 3236 20380 3292
rect 20380 3236 20436 3292
rect 20436 3236 20440 3292
rect 20376 3232 20440 3236
rect 20456 3292 20520 3296
rect 20456 3236 20460 3292
rect 20460 3236 20516 3292
rect 20516 3236 20520 3292
rect 20456 3232 20520 3236
rect 39480 3292 39544 3296
rect 39480 3236 39484 3292
rect 39484 3236 39540 3292
rect 39540 3236 39544 3292
rect 39480 3232 39544 3236
rect 39560 3292 39624 3296
rect 39560 3236 39564 3292
rect 39564 3236 39620 3292
rect 39620 3236 39624 3292
rect 39560 3232 39624 3236
rect 39640 3292 39704 3296
rect 39640 3236 39644 3292
rect 39644 3236 39700 3292
rect 39700 3236 39704 3292
rect 39640 3232 39704 3236
rect 39720 3292 39784 3296
rect 39720 3236 39724 3292
rect 39724 3236 39780 3292
rect 39780 3236 39784 3292
rect 39720 3232 39784 3236
rect 10584 2748 10648 2752
rect 10584 2692 10588 2748
rect 10588 2692 10644 2748
rect 10644 2692 10648 2748
rect 10584 2688 10648 2692
rect 10664 2748 10728 2752
rect 10664 2692 10668 2748
rect 10668 2692 10724 2748
rect 10724 2692 10728 2748
rect 10664 2688 10728 2692
rect 10744 2748 10808 2752
rect 10744 2692 10748 2748
rect 10748 2692 10804 2748
rect 10804 2692 10808 2748
rect 10744 2688 10808 2692
rect 10824 2748 10888 2752
rect 10824 2692 10828 2748
rect 10828 2692 10884 2748
rect 10884 2692 10888 2748
rect 10824 2688 10888 2692
rect 29848 2748 29912 2752
rect 29848 2692 29852 2748
rect 29852 2692 29908 2748
rect 29908 2692 29912 2748
rect 29848 2688 29912 2692
rect 29928 2748 29992 2752
rect 29928 2692 29932 2748
rect 29932 2692 29988 2748
rect 29988 2692 29992 2748
rect 29928 2688 29992 2692
rect 30008 2748 30072 2752
rect 30008 2692 30012 2748
rect 30012 2692 30068 2748
rect 30068 2692 30072 2748
rect 30008 2688 30072 2692
rect 30088 2748 30152 2752
rect 30088 2692 30092 2748
rect 30092 2692 30148 2748
rect 30148 2692 30152 2748
rect 30088 2688 30152 2692
rect 49112 2748 49176 2752
rect 49112 2692 49116 2748
rect 49116 2692 49172 2748
rect 49172 2692 49176 2748
rect 49112 2688 49176 2692
rect 49192 2748 49256 2752
rect 49192 2692 49196 2748
rect 49196 2692 49252 2748
rect 49252 2692 49256 2748
rect 49192 2688 49256 2692
rect 49272 2748 49336 2752
rect 49272 2692 49276 2748
rect 49276 2692 49332 2748
rect 49332 2692 49336 2748
rect 49272 2688 49336 2692
rect 49352 2748 49416 2752
rect 49352 2692 49356 2748
rect 49356 2692 49412 2748
rect 49412 2692 49416 2748
rect 49352 2688 49416 2692
rect 20216 2204 20280 2208
rect 20216 2148 20220 2204
rect 20220 2148 20276 2204
rect 20276 2148 20280 2204
rect 20216 2144 20280 2148
rect 20296 2204 20360 2208
rect 20296 2148 20300 2204
rect 20300 2148 20356 2204
rect 20356 2148 20360 2204
rect 20296 2144 20360 2148
rect 20376 2204 20440 2208
rect 20376 2148 20380 2204
rect 20380 2148 20436 2204
rect 20436 2148 20440 2204
rect 20376 2144 20440 2148
rect 20456 2204 20520 2208
rect 20456 2148 20460 2204
rect 20460 2148 20516 2204
rect 20516 2148 20520 2204
rect 20456 2144 20520 2148
rect 39480 2204 39544 2208
rect 39480 2148 39484 2204
rect 39484 2148 39540 2204
rect 39540 2148 39544 2204
rect 39480 2144 39544 2148
rect 39560 2204 39624 2208
rect 39560 2148 39564 2204
rect 39564 2148 39620 2204
rect 39620 2148 39624 2204
rect 39560 2144 39624 2148
rect 39640 2204 39704 2208
rect 39640 2148 39644 2204
rect 39644 2148 39700 2204
rect 39700 2148 39704 2204
rect 39640 2144 39704 2148
rect 39720 2204 39784 2208
rect 39720 2148 39724 2204
rect 39724 2148 39780 2204
rect 39780 2148 39784 2204
rect 39720 2144 39784 2148
<< metal4 >>
rect 10576 19072 10896 19632
rect 10576 19008 10584 19072
rect 10648 19008 10664 19072
rect 10728 19008 10744 19072
rect 10808 19008 10824 19072
rect 10888 19008 10896 19072
rect 10576 17984 10896 19008
rect 10576 17920 10584 17984
rect 10648 17920 10664 17984
rect 10728 17920 10744 17984
rect 10808 17920 10824 17984
rect 10888 17920 10896 17984
rect 10576 16896 10896 17920
rect 10576 16832 10584 16896
rect 10648 16832 10664 16896
rect 10728 16832 10744 16896
rect 10808 16832 10824 16896
rect 10888 16832 10896 16896
rect 10576 15808 10896 16832
rect 10576 15744 10584 15808
rect 10648 15744 10664 15808
rect 10728 15744 10744 15808
rect 10808 15744 10824 15808
rect 10888 15744 10896 15808
rect 10576 14720 10896 15744
rect 10576 14656 10584 14720
rect 10648 14656 10664 14720
rect 10728 14656 10744 14720
rect 10808 14656 10824 14720
rect 10888 14656 10896 14720
rect 10576 13632 10896 14656
rect 10576 13568 10584 13632
rect 10648 13568 10664 13632
rect 10728 13568 10744 13632
rect 10808 13568 10824 13632
rect 10888 13568 10896 13632
rect 10576 12544 10896 13568
rect 10576 12480 10584 12544
rect 10648 12480 10664 12544
rect 10728 12480 10744 12544
rect 10808 12480 10824 12544
rect 10888 12480 10896 12544
rect 10576 11456 10896 12480
rect 10576 11392 10584 11456
rect 10648 11392 10664 11456
rect 10728 11392 10744 11456
rect 10808 11392 10824 11456
rect 10888 11392 10896 11456
rect 10576 10368 10896 11392
rect 10576 10304 10584 10368
rect 10648 10304 10664 10368
rect 10728 10304 10744 10368
rect 10808 10304 10824 10368
rect 10888 10304 10896 10368
rect 10576 9280 10896 10304
rect 10576 9216 10584 9280
rect 10648 9216 10664 9280
rect 10728 9216 10744 9280
rect 10808 9216 10824 9280
rect 10888 9216 10896 9280
rect 10576 8192 10896 9216
rect 10576 8128 10584 8192
rect 10648 8128 10664 8192
rect 10728 8128 10744 8192
rect 10808 8128 10824 8192
rect 10888 8128 10896 8192
rect 10576 7104 10896 8128
rect 10576 7040 10584 7104
rect 10648 7040 10664 7104
rect 10728 7040 10744 7104
rect 10808 7040 10824 7104
rect 10888 7040 10896 7104
rect 10576 6016 10896 7040
rect 10576 5952 10584 6016
rect 10648 5952 10664 6016
rect 10728 5952 10744 6016
rect 10808 5952 10824 6016
rect 10888 5952 10896 6016
rect 10576 4928 10896 5952
rect 10576 4864 10584 4928
rect 10648 4864 10664 4928
rect 10728 4864 10744 4928
rect 10808 4864 10824 4928
rect 10888 4864 10896 4928
rect 10576 3840 10896 4864
rect 10576 3776 10584 3840
rect 10648 3776 10664 3840
rect 10728 3776 10744 3840
rect 10808 3776 10824 3840
rect 10888 3776 10896 3840
rect 10576 2752 10896 3776
rect 10576 2688 10584 2752
rect 10648 2688 10664 2752
rect 10728 2688 10744 2752
rect 10808 2688 10824 2752
rect 10888 2688 10896 2752
rect 10576 2128 10896 2688
rect 20208 19616 20528 19632
rect 20208 19552 20216 19616
rect 20280 19552 20296 19616
rect 20360 19552 20376 19616
rect 20440 19552 20456 19616
rect 20520 19552 20528 19616
rect 20208 18528 20528 19552
rect 20208 18464 20216 18528
rect 20280 18464 20296 18528
rect 20360 18464 20376 18528
rect 20440 18464 20456 18528
rect 20520 18464 20528 18528
rect 20208 17440 20528 18464
rect 20208 17376 20216 17440
rect 20280 17376 20296 17440
rect 20360 17376 20376 17440
rect 20440 17376 20456 17440
rect 20520 17376 20528 17440
rect 20208 16352 20528 17376
rect 20208 16288 20216 16352
rect 20280 16288 20296 16352
rect 20360 16288 20376 16352
rect 20440 16288 20456 16352
rect 20520 16288 20528 16352
rect 20208 15264 20528 16288
rect 20208 15200 20216 15264
rect 20280 15200 20296 15264
rect 20360 15200 20376 15264
rect 20440 15200 20456 15264
rect 20520 15200 20528 15264
rect 20208 14176 20528 15200
rect 20208 14112 20216 14176
rect 20280 14112 20296 14176
rect 20360 14112 20376 14176
rect 20440 14112 20456 14176
rect 20520 14112 20528 14176
rect 20208 13088 20528 14112
rect 20208 13024 20216 13088
rect 20280 13024 20296 13088
rect 20360 13024 20376 13088
rect 20440 13024 20456 13088
rect 20520 13024 20528 13088
rect 20208 12000 20528 13024
rect 20208 11936 20216 12000
rect 20280 11936 20296 12000
rect 20360 11936 20376 12000
rect 20440 11936 20456 12000
rect 20520 11936 20528 12000
rect 20208 10912 20528 11936
rect 20208 10848 20216 10912
rect 20280 10848 20296 10912
rect 20360 10848 20376 10912
rect 20440 10848 20456 10912
rect 20520 10848 20528 10912
rect 20208 9824 20528 10848
rect 20208 9760 20216 9824
rect 20280 9760 20296 9824
rect 20360 9760 20376 9824
rect 20440 9760 20456 9824
rect 20520 9760 20528 9824
rect 20208 8736 20528 9760
rect 20208 8672 20216 8736
rect 20280 8672 20296 8736
rect 20360 8672 20376 8736
rect 20440 8672 20456 8736
rect 20520 8672 20528 8736
rect 20208 7648 20528 8672
rect 20208 7584 20216 7648
rect 20280 7584 20296 7648
rect 20360 7584 20376 7648
rect 20440 7584 20456 7648
rect 20520 7584 20528 7648
rect 20208 6560 20528 7584
rect 20208 6496 20216 6560
rect 20280 6496 20296 6560
rect 20360 6496 20376 6560
rect 20440 6496 20456 6560
rect 20520 6496 20528 6560
rect 20208 5472 20528 6496
rect 20208 5408 20216 5472
rect 20280 5408 20296 5472
rect 20360 5408 20376 5472
rect 20440 5408 20456 5472
rect 20520 5408 20528 5472
rect 20208 4384 20528 5408
rect 20208 4320 20216 4384
rect 20280 4320 20296 4384
rect 20360 4320 20376 4384
rect 20440 4320 20456 4384
rect 20520 4320 20528 4384
rect 20208 3296 20528 4320
rect 20208 3232 20216 3296
rect 20280 3232 20296 3296
rect 20360 3232 20376 3296
rect 20440 3232 20456 3296
rect 20520 3232 20528 3296
rect 20208 2208 20528 3232
rect 20208 2144 20216 2208
rect 20280 2144 20296 2208
rect 20360 2144 20376 2208
rect 20440 2144 20456 2208
rect 20520 2144 20528 2208
rect 20208 2128 20528 2144
rect 29840 19072 30160 19632
rect 29840 19008 29848 19072
rect 29912 19008 29928 19072
rect 29992 19008 30008 19072
rect 30072 19008 30088 19072
rect 30152 19008 30160 19072
rect 29840 17984 30160 19008
rect 29840 17920 29848 17984
rect 29912 17920 29928 17984
rect 29992 17920 30008 17984
rect 30072 17920 30088 17984
rect 30152 17920 30160 17984
rect 29840 16896 30160 17920
rect 29840 16832 29848 16896
rect 29912 16832 29928 16896
rect 29992 16832 30008 16896
rect 30072 16832 30088 16896
rect 30152 16832 30160 16896
rect 29840 15808 30160 16832
rect 29840 15744 29848 15808
rect 29912 15744 29928 15808
rect 29992 15744 30008 15808
rect 30072 15744 30088 15808
rect 30152 15744 30160 15808
rect 29840 14720 30160 15744
rect 29840 14656 29848 14720
rect 29912 14656 29928 14720
rect 29992 14656 30008 14720
rect 30072 14656 30088 14720
rect 30152 14656 30160 14720
rect 29840 13632 30160 14656
rect 29840 13568 29848 13632
rect 29912 13568 29928 13632
rect 29992 13568 30008 13632
rect 30072 13568 30088 13632
rect 30152 13568 30160 13632
rect 29840 12544 30160 13568
rect 29840 12480 29848 12544
rect 29912 12480 29928 12544
rect 29992 12480 30008 12544
rect 30072 12480 30088 12544
rect 30152 12480 30160 12544
rect 29840 11456 30160 12480
rect 29840 11392 29848 11456
rect 29912 11392 29928 11456
rect 29992 11392 30008 11456
rect 30072 11392 30088 11456
rect 30152 11392 30160 11456
rect 29840 10368 30160 11392
rect 29840 10304 29848 10368
rect 29912 10304 29928 10368
rect 29992 10304 30008 10368
rect 30072 10304 30088 10368
rect 30152 10304 30160 10368
rect 29840 9280 30160 10304
rect 29840 9216 29848 9280
rect 29912 9216 29928 9280
rect 29992 9216 30008 9280
rect 30072 9216 30088 9280
rect 30152 9216 30160 9280
rect 29840 8192 30160 9216
rect 29840 8128 29848 8192
rect 29912 8128 29928 8192
rect 29992 8128 30008 8192
rect 30072 8128 30088 8192
rect 30152 8128 30160 8192
rect 29840 7104 30160 8128
rect 29840 7040 29848 7104
rect 29912 7040 29928 7104
rect 29992 7040 30008 7104
rect 30072 7040 30088 7104
rect 30152 7040 30160 7104
rect 29840 6016 30160 7040
rect 29840 5952 29848 6016
rect 29912 5952 29928 6016
rect 29992 5952 30008 6016
rect 30072 5952 30088 6016
rect 30152 5952 30160 6016
rect 29840 4928 30160 5952
rect 29840 4864 29848 4928
rect 29912 4864 29928 4928
rect 29992 4864 30008 4928
rect 30072 4864 30088 4928
rect 30152 4864 30160 4928
rect 29840 3840 30160 4864
rect 29840 3776 29848 3840
rect 29912 3776 29928 3840
rect 29992 3776 30008 3840
rect 30072 3776 30088 3840
rect 30152 3776 30160 3840
rect 29840 2752 30160 3776
rect 29840 2688 29848 2752
rect 29912 2688 29928 2752
rect 29992 2688 30008 2752
rect 30072 2688 30088 2752
rect 30152 2688 30160 2752
rect 29840 2128 30160 2688
rect 39472 19616 39792 19632
rect 39472 19552 39480 19616
rect 39544 19552 39560 19616
rect 39624 19552 39640 19616
rect 39704 19552 39720 19616
rect 39784 19552 39792 19616
rect 39472 18528 39792 19552
rect 39472 18464 39480 18528
rect 39544 18464 39560 18528
rect 39624 18464 39640 18528
rect 39704 18464 39720 18528
rect 39784 18464 39792 18528
rect 39472 17440 39792 18464
rect 39472 17376 39480 17440
rect 39544 17376 39560 17440
rect 39624 17376 39640 17440
rect 39704 17376 39720 17440
rect 39784 17376 39792 17440
rect 39472 16352 39792 17376
rect 39472 16288 39480 16352
rect 39544 16288 39560 16352
rect 39624 16288 39640 16352
rect 39704 16288 39720 16352
rect 39784 16288 39792 16352
rect 39472 15264 39792 16288
rect 39472 15200 39480 15264
rect 39544 15200 39560 15264
rect 39624 15200 39640 15264
rect 39704 15200 39720 15264
rect 39784 15200 39792 15264
rect 39472 14176 39792 15200
rect 39472 14112 39480 14176
rect 39544 14112 39560 14176
rect 39624 14112 39640 14176
rect 39704 14112 39720 14176
rect 39784 14112 39792 14176
rect 39472 13088 39792 14112
rect 39472 13024 39480 13088
rect 39544 13024 39560 13088
rect 39624 13024 39640 13088
rect 39704 13024 39720 13088
rect 39784 13024 39792 13088
rect 39472 12000 39792 13024
rect 39472 11936 39480 12000
rect 39544 11936 39560 12000
rect 39624 11936 39640 12000
rect 39704 11936 39720 12000
rect 39784 11936 39792 12000
rect 39472 10912 39792 11936
rect 39472 10848 39480 10912
rect 39544 10848 39560 10912
rect 39624 10848 39640 10912
rect 39704 10848 39720 10912
rect 39784 10848 39792 10912
rect 39472 9824 39792 10848
rect 39472 9760 39480 9824
rect 39544 9760 39560 9824
rect 39624 9760 39640 9824
rect 39704 9760 39720 9824
rect 39784 9760 39792 9824
rect 39472 8736 39792 9760
rect 39472 8672 39480 8736
rect 39544 8672 39560 8736
rect 39624 8672 39640 8736
rect 39704 8672 39720 8736
rect 39784 8672 39792 8736
rect 39472 7648 39792 8672
rect 39472 7584 39480 7648
rect 39544 7584 39560 7648
rect 39624 7584 39640 7648
rect 39704 7584 39720 7648
rect 39784 7584 39792 7648
rect 39472 6560 39792 7584
rect 39472 6496 39480 6560
rect 39544 6496 39560 6560
rect 39624 6496 39640 6560
rect 39704 6496 39720 6560
rect 39784 6496 39792 6560
rect 39472 5472 39792 6496
rect 39472 5408 39480 5472
rect 39544 5408 39560 5472
rect 39624 5408 39640 5472
rect 39704 5408 39720 5472
rect 39784 5408 39792 5472
rect 39472 4384 39792 5408
rect 39472 4320 39480 4384
rect 39544 4320 39560 4384
rect 39624 4320 39640 4384
rect 39704 4320 39720 4384
rect 39784 4320 39792 4384
rect 39472 3296 39792 4320
rect 39472 3232 39480 3296
rect 39544 3232 39560 3296
rect 39624 3232 39640 3296
rect 39704 3232 39720 3296
rect 39784 3232 39792 3296
rect 39472 2208 39792 3232
rect 39472 2144 39480 2208
rect 39544 2144 39560 2208
rect 39624 2144 39640 2208
rect 39704 2144 39720 2208
rect 39784 2144 39792 2208
rect 39472 2128 39792 2144
rect 49104 19072 49424 19632
rect 49104 19008 49112 19072
rect 49176 19008 49192 19072
rect 49256 19008 49272 19072
rect 49336 19008 49352 19072
rect 49416 19008 49424 19072
rect 49104 17984 49424 19008
rect 49104 17920 49112 17984
rect 49176 17920 49192 17984
rect 49256 17920 49272 17984
rect 49336 17920 49352 17984
rect 49416 17920 49424 17984
rect 49104 16896 49424 17920
rect 49104 16832 49112 16896
rect 49176 16832 49192 16896
rect 49256 16832 49272 16896
rect 49336 16832 49352 16896
rect 49416 16832 49424 16896
rect 49104 15808 49424 16832
rect 49104 15744 49112 15808
rect 49176 15744 49192 15808
rect 49256 15744 49272 15808
rect 49336 15744 49352 15808
rect 49416 15744 49424 15808
rect 49104 14720 49424 15744
rect 49104 14656 49112 14720
rect 49176 14656 49192 14720
rect 49256 14656 49272 14720
rect 49336 14656 49352 14720
rect 49416 14656 49424 14720
rect 49104 13632 49424 14656
rect 49104 13568 49112 13632
rect 49176 13568 49192 13632
rect 49256 13568 49272 13632
rect 49336 13568 49352 13632
rect 49416 13568 49424 13632
rect 49104 12544 49424 13568
rect 49104 12480 49112 12544
rect 49176 12480 49192 12544
rect 49256 12480 49272 12544
rect 49336 12480 49352 12544
rect 49416 12480 49424 12544
rect 49104 11456 49424 12480
rect 49104 11392 49112 11456
rect 49176 11392 49192 11456
rect 49256 11392 49272 11456
rect 49336 11392 49352 11456
rect 49416 11392 49424 11456
rect 49104 10368 49424 11392
rect 49104 10304 49112 10368
rect 49176 10304 49192 10368
rect 49256 10304 49272 10368
rect 49336 10304 49352 10368
rect 49416 10304 49424 10368
rect 49104 9280 49424 10304
rect 49104 9216 49112 9280
rect 49176 9216 49192 9280
rect 49256 9216 49272 9280
rect 49336 9216 49352 9280
rect 49416 9216 49424 9280
rect 49104 8192 49424 9216
rect 49104 8128 49112 8192
rect 49176 8128 49192 8192
rect 49256 8128 49272 8192
rect 49336 8128 49352 8192
rect 49416 8128 49424 8192
rect 49104 7104 49424 8128
rect 49104 7040 49112 7104
rect 49176 7040 49192 7104
rect 49256 7040 49272 7104
rect 49336 7040 49352 7104
rect 49416 7040 49424 7104
rect 49104 6016 49424 7040
rect 49104 5952 49112 6016
rect 49176 5952 49192 6016
rect 49256 5952 49272 6016
rect 49336 5952 49352 6016
rect 49416 5952 49424 6016
rect 49104 4928 49424 5952
rect 49104 4864 49112 4928
rect 49176 4864 49192 4928
rect 49256 4864 49272 4928
rect 49336 4864 49352 4928
rect 49416 4864 49424 4928
rect 49104 3840 49424 4864
rect 49104 3776 49112 3840
rect 49176 3776 49192 3840
rect 49256 3776 49272 3840
rect 49336 3776 49352 3840
rect 49416 3776 49424 3840
rect 49104 2752 49424 3776
rect 49104 2688 49112 2752
rect 49176 2688 49192 2752
rect 49256 2688 49272 2752
rect 49336 2688 49352 2752
rect 49416 2688 49424 2752
rect 49104 2128 49424 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 57408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 57408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 57408 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1644511149
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44
timestamp 1644511149
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1644511149
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1644511149
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1644511149
transform 1 0 9200 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1644511149
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_132 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_154 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_172
timestamp 1644511149
transform 1 0 16928 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_180
timestamp 1644511149
transform 1 0 17664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_185
timestamp 1644511149
transform 1 0 18124 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_200
timestamp 1644511149
transform 1 0 19504 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_212
timestamp 1644511149
transform 1 0 20608 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216
timestamp 1644511149
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_231
timestamp 1644511149
transform 1 0 22356 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_243
timestamp 1644511149
transform 1 0 23460 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1644511149
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_262
timestamp 1644511149
transform 1 0 25208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_274
timestamp 1644511149
transform 1 0 26312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_284
timestamp 1644511149
transform 1 0 27232 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_312
timestamp 1644511149
transform 1 0 29808 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_320
timestamp 1644511149
transform 1 0 30544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_325
timestamp 1644511149
transform 1 0 31004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_340
timestamp 1644511149
transform 1 0 32384 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_352
timestamp 1644511149
transform 1 0 33488 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_356
timestamp 1644511149
transform 1 0 33856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_371
timestamp 1644511149
transform 1 0 35236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_383
timestamp 1644511149
transform 1 0 36340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_387
timestamp 1644511149
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_402
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_414
timestamp 1644511149
transform 1 0 39192 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_424
timestamp 1644511149
transform 1 0 40112 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_452
timestamp 1644511149
transform 1 0 42688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_460
timestamp 1644511149
transform 1 0 43424 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_464
timestamp 1644511149
transform 1 0 43792 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_480
timestamp 1644511149
transform 1 0 45264 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_495
timestamp 1644511149
transform 1 0 46644 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1644511149
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_518
timestamp 1644511149
transform 1 0 48760 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1644511149
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_549
timestamp 1644511149
transform 1 0 51612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1644511149
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_571
timestamp 1644511149
transform 1 0 53636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_577
timestamp 1644511149
transform 1 0 54188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_584
timestamp 1644511149
transform 1 0 54832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_599
timestamp 1644511149
transform 1 0 56212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_605
timestamp 1644511149
transform 1 0 56764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_612
timestamp 1644511149
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_617
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_14
timestamp 1644511149
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1644511149
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32
timestamp 1644511149
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_36
timestamp 1644511149
transform 1 0 4416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1644511149
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_50
timestamp 1644511149
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_63
timestamp 1644511149
transform 1 0 6900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_72
timestamp 1644511149
transform 1 0 7728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_79
timestamp 1644511149
transform 1 0 8372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 1644511149
transform 1 0 8924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1644511149
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_98
timestamp 1644511149
transform 1 0 10120 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1644511149
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_117
timestamp 1644511149
transform 1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_124
timestamp 1644511149
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp 1644511149
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_140
timestamp 1644511149
transform 1 0 13984 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_152
timestamp 1644511149
transform 1 0 15088 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1644511149
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_429
timestamp 1644511149
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1644511149
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_461
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_473
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1644511149
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_533
timestamp 1644511149
transform 1 0 50140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_545
timestamp 1644511149
transform 1 0 51244 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_557
timestamp 1644511149
transform 1 0 52348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_569
timestamp 1644511149
transform 1 0 53452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_580
timestamp 1644511149
transform 1 0 54464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_588
timestamp 1644511149
transform 1 0 55200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_597
timestamp 1644511149
transform 1 0 56028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_611
timestamp 1644511149
transform 1 0 57316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_617
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_35
timestamp 1644511149
transform 1 0 4324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_39
timestamp 1644511149
transform 1 0 4692 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1644511149
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_54
timestamp 1644511149
transform 1 0 6072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_58
timestamp 1644511149
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1644511149
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75
timestamp 1644511149
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_90
timestamp 1644511149
transform 1 0 9384 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1644511149
transform 1 0 10488 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_107
timestamp 1644511149
transform 1 0 10948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_114
timestamp 1644511149
transform 1 0 11592 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_126
timestamp 1644511149
transform 1 0 12696 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1644511149
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_489
timestamp 1644511149
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_501
timestamp 1644511149
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_513
timestamp 1644511149
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_597
timestamp 1644511149
transform 1 0 56028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_607
timestamp 1644511149
transform 1 0 56948 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1644511149
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1644511149
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_30
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1644511149
transform 1 0 5152 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_67
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_593
timestamp 1644511149
transform 1 0 55660 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_602
timestamp 1644511149
transform 1 0 56488 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_612
timestamp 1644511149
transform 1 0 57408 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_607
timestamp 1644511149
transform 1 0 56948 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_621
timestamp 1644511149
transform 1 0 58236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_605
timestamp 1644511149
transform 1 0 56764 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_612
timestamp 1644511149
transform 1 0 57408 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_611
timestamp 1644511149
transform 1 0 57316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_621
timestamp 1644511149
transform 1 0 58236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1644511149
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_173
timestamp 1644511149
transform 1 0 17020 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_185
timestamp 1644511149
transform 1 0 18124 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_190
timestamp 1644511149
transform 1 0 18584 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1644511149
transform 1 0 19688 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_214
timestamp 1644511149
transform 1 0 20792 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1644511149
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1644511149
transform 1 0 58236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_161
timestamp 1644511149
transform 1 0 15916 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_171
timestamp 1644511149
transform 1 0 16836 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_187
timestamp 1644511149
transform 1 0 18308 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_205
timestamp 1644511149
transform 1 0 19964 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_217
timestamp 1644511149
transform 1 0 21068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_229
timestamp 1644511149
transform 1 0 22172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_241
timestamp 1644511149
transform 1 0 23276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1644511149
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_621
timestamp 1644511149
transform 1 0 58236 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_89
timestamp 1644511149
transform 1 0 9292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_96
timestamp 1644511149
transform 1 0 9936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1644511149
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_203
timestamp 1644511149
transform 1 0 19780 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1644511149
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1644511149
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_621
timestamp 1644511149
transform 1 0 58236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1644511149
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp 1644511149
transform 1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_100
timestamp 1644511149
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_108
timestamp 1644511149
transform 1 0 11040 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_116
timestamp 1644511149
transform 1 0 11776 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1644511149
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1644511149
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_207
timestamp 1644511149
transform 1 0 20148 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1644511149
transform 1 0 20700 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_218
timestamp 1644511149
transform 1 0 21160 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_230
timestamp 1644511149
transform 1 0 22264 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_242
timestamp 1644511149
transform 1 0 23368 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1644511149
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_615
timestamp 1644511149
transform 1 0 57684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_621
timestamp 1644511149
transform 1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1644511149
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1644511149
transform 1 0 9752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1644511149
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_133
timestamp 1644511149
transform 1 0 13340 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_231
timestamp 1644511149
transform 1 0 22356 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_236
timestamp 1644511149
transform 1 0 22816 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_614
timestamp 1644511149
transform 1 0 57592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_621
timestamp 1644511149
transform 1 0 58236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_106
timestamp 1644511149
transform 1 0 10856 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_118
timestamp 1644511149
transform 1 0 11960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_122
timestamp 1644511149
transform 1 0 12328 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1644511149
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1644511149
transform 1 0 14352 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_156
timestamp 1644511149
transform 1 0 15456 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_168
timestamp 1644511149
transform 1 0 16560 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_180
timestamp 1644511149
transform 1 0 17664 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1644511149
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_238
timestamp 1644511149
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1644511149
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_257
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_269
timestamp 1644511149
transform 1 0 25852 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_279
timestamp 1644511149
transform 1 0 26772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_292
timestamp 1644511149
transform 1 0 27968 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1644511149
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1644511149
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_264
timestamp 1644511149
transform 1 0 25392 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_272
timestamp 1644511149
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_290
timestamp 1644511149
transform 1 0 27784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_302
timestamp 1644511149
transform 1 0 28888 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_314
timestamp 1644511149
transform 1 0 29992 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_326
timestamp 1644511149
transform 1 0 31096 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_334
timestamp 1644511149
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_621
timestamp 1644511149
transform 1 0 58236 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_283
timestamp 1644511149
transform 1 0 27140 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_295
timestamp 1644511149
transform 1 0 28244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_615
timestamp 1644511149
transform 1 0 57684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_621
timestamp 1644511149
transform 1 0 58236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_605
timestamp 1644511149
transform 1 0 56764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_612
timestamp 1644511149
transform 1 0 57408 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1644511149
transform 1 0 58236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_319
timestamp 1644511149
transform 1 0 30452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_327
timestamp 1644511149
transform 1 0 31188 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_339
timestamp 1644511149
transform 1 0 32292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_351
timestamp 1644511149
transform 1 0 33396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_427
timestamp 1644511149
transform 1 0 40388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_439
timestamp 1644511149
transform 1 0 41492 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_451
timestamp 1644511149
transform 1 0 42596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_463
timestamp 1644511149
transform 1 0 43700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_621
timestamp 1644511149
transform 1 0 58236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_330
timestamp 1644511149
transform 1 0 31464 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_346
timestamp 1644511149
transform 1 0 32936 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_354
timestamp 1644511149
transform 1 0 33672 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_621
timestamp 1644511149
transform 1 0 58236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_325
timestamp 1644511149
transform 1 0 31004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_330
timestamp 1644511149
transform 1 0 31464 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_338
timestamp 1644511149
transform 1 0 32200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_349
timestamp 1644511149
transform 1 0 33212 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 1644511149
transform 1 0 34132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_374
timestamp 1644511149
transform 1 0 35512 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_386
timestamp 1644511149
transform 1 0 36616 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_398
timestamp 1644511149
transform 1 0 37720 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_406
timestamp 1644511149
transform 1 0 38456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_412
timestamp 1644511149
transform 1 0 39008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_621
timestamp 1644511149
transform 1 0 58236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_401
timestamp 1644511149
transform 1 0 37996 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_406
timestamp 1644511149
transform 1 0 38456 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_418
timestamp 1644511149
transform 1 0 39560 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_430
timestamp 1644511149
transform 1 0 40664 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_442
timestamp 1644511149
transform 1 0 41768 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_614
timestamp 1644511149
transform 1 0 57592 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_621
timestamp 1644511149
transform 1 0 58236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_403
timestamp 1644511149
transform 1 0 38180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_415
timestamp 1644511149
transform 1 0 39284 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_621
timestamp 1644511149
transform 1 0 58236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_401
timestamp 1644511149
transform 1 0 37996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_413
timestamp 1644511149
transform 1 0 39100 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_425
timestamp 1644511149
transform 1 0 40204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_437
timestamp 1644511149
transform 1 0 41308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1644511149
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_621
timestamp 1644511149
transform 1 0 58236 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_404
timestamp 1644511149
transform 1 0 38272 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_416
timestamp 1644511149
transform 1 0 39376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_431
timestamp 1644511149
transform 1 0 40756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_444
timestamp 1644511149
transform 1 0 41952 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_456
timestamp 1644511149
transform 1 0 43056 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_468
timestamp 1644511149
transform 1 0 44160 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1644511149
transform 1 0 58236 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_420
timestamp 1644511149
transform 1 0 39744 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_432
timestamp 1644511149
transform 1 0 40848 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_444
timestamp 1644511149
transform 1 0 41952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_459
timestamp 1644511149
transform 1 0 43332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_471
timestamp 1644511149
transform 1 0 44436 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_483
timestamp 1644511149
transform 1 0 45540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_495
timestamp 1644511149
transform 1 0 46644 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_621
timestamp 1644511149
transform 1 0 58236 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_448
timestamp 1644511149
transform 1 0 42320 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_460
timestamp 1644511149
transform 1 0 43424 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_472
timestamp 1644511149
transform 1 0 44528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_621
timestamp 1644511149
transform 1 0 58236 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_469
timestamp 1644511149
transform 1 0 44252 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_612
timestamp 1644511149
transform 1 0 57408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1644511149
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_461
timestamp 1644511149
transform 1 0 43516 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_471
timestamp 1644511149
transform 1 0 44436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_486
timestamp 1644511149
transform 1 0 45816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_493
timestamp 1644511149
transform 1 0 46460 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_505
timestamp 1644511149
transform 1 0 47564 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_517
timestamp 1644511149
transform 1 0 48668 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_529
timestamp 1644511149
transform 1 0 49772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_606
timestamp 1644511149
transform 1 0 56856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_621
timestamp 1644511149
transform 1 0 58236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_479
timestamp 1644511149
transform 1 0 45172 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_487
timestamp 1644511149
transform 1 0 45908 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_514
timestamp 1644511149
transform 1 0 48392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_526
timestamp 1644511149
transform 1 0 49496 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_538
timestamp 1644511149
transform 1 0 50600 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_550
timestamp 1644511149
transform 1 0 51704 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_558
timestamp 1644511149
transform 1 0 52440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_604
timestamp 1644511149
transform 1 0 56672 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_612
timestamp 1644511149
transform 1 0 57408 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1644511149
transform 1 0 58236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_495
timestamp 1644511149
transform 1 0 46644 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_499
timestamp 1644511149
transform 1 0 47012 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_507
timestamp 1644511149
transform 1 0 47748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_512
timestamp 1644511149
transform 1 0 48208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_536
timestamp 1644511149
transform 1 0 50416 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_548
timestamp 1644511149
transform 1 0 51520 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_560
timestamp 1644511149
transform 1 0 52624 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_572
timestamp 1644511149
transform 1 0 53728 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_584
timestamp 1644511149
transform 1 0 54832 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_597
timestamp 1644511149
transform 1 0 56028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_605
timestamp 1644511149
transform 1 0 56764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_618
timestamp 1644511149
transform 1 0 57960 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_624
timestamp 1644511149
transform 1 0 58512 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_547
timestamp 1644511149
transform 1 0 51428 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_551
timestamp 1644511149
transform 1 0 51796 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_564
timestamp 1644511149
transform 1 0 52992 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_584
timestamp 1644511149
transform 1 0 54832 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_591
timestamp 1644511149
transform 1 0 55476 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_599
timestamp 1644511149
transform 1 0 56212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_612
timestamp 1644511149
transform 1 0 57408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_621
timestamp 1644511149
transform 1 0 58236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_539
timestamp 1644511149
transform 1 0 50692 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_549
timestamp 1644511149
transform 1 0 51612 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_562
timestamp 1644511149
transform 1 0 52808 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_575
timestamp 1644511149
transform 1 0 54004 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_584
timestamp 1644511149
transform 1 0 54832 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_598
timestamp 1644511149
transform 1 0 56120 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_611
timestamp 1644511149
transform 1 0 57316 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_621
timestamp 1644511149
transform 1 0 58236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_7
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_33
timestamp 1644511149
transform 1 0 4140 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_41
timestamp 1644511149
transform 1 0 4876 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_46
timestamp 1644511149
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1644511149
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_62
timestamp 1644511149
transform 1 0 6808 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_70
timestamp 1644511149
transform 1 0 7544 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_77
timestamp 1644511149
transform 1 0 8188 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_83
timestamp 1644511149
transform 1 0 8740 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_85
timestamp 1644511149
transform 1 0 8924 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_101
timestamp 1644511149
transform 1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_119
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_124
timestamp 1644511149
transform 1 0 12512 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_136
timestamp 1644511149
transform 1 0 13616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_145
timestamp 1644511149
transform 1 0 14444 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_154
timestamp 1644511149
transform 1 0 15272 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1644511149
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_180
timestamp 1644511149
transform 1 0 17664 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_185
timestamp 1644511149
transform 1 0 18124 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_200
timestamp 1644511149
transform 1 0 19504 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_212
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_231
timestamp 1644511149
transform 1 0 22356 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_243
timestamp 1644511149
transform 1 0 23460 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_247
timestamp 1644511149
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_251
timestamp 1644511149
transform 1 0 24196 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_253
timestamp 1644511149
transform 1 0 24380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_262
timestamp 1644511149
transform 1 0 25208 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1644511149
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_284
timestamp 1644511149
transform 1 0 27232 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_312
timestamp 1644511149
transform 1 0 29808 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_320
timestamp 1644511149
transform 1 0 30544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_325
timestamp 1644511149
transform 1 0 31004 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1644511149
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_340
timestamp 1644511149
transform 1 0 32384 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_352
timestamp 1644511149
transform 1 0 33488 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_356
timestamp 1644511149
transform 1 0 33856 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_365
timestamp 1644511149
transform 1 0 34684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_371
timestamp 1644511149
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_383
timestamp 1644511149
transform 1 0 36340 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1644511149
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_402
timestamp 1644511149
transform 1 0 38088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_414
timestamp 1644511149
transform 1 0 39192 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_424
timestamp 1644511149
transform 1 0 40112 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_433
timestamp 1644511149
transform 1 0 40940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1644511149
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_452
timestamp 1644511149
transform 1 0 42688 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_460
timestamp 1644511149
transform 1 0 43424 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_464
timestamp 1644511149
transform 1 0 43792 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_480
timestamp 1644511149
transform 1 0 45264 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_495
timestamp 1644511149
transform 1 0 46644 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_511
timestamp 1644511149
transform 1 0 48116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_526
timestamp 1644511149
transform 1 0 49496 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_533
timestamp 1644511149
transform 1 0 50140 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_542
timestamp 1644511149
transform 1 0 50968 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_550
timestamp 1644511149
transform 1 0 51704 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_556
timestamp 1644511149
transform 1 0 52256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_565
timestamp 1644511149
transform 1 0 53084 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_569
timestamp 1644511149
transform 1 0 53452 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_576
timestamp 1644511149
transform 1 0 54096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_584
timestamp 1644511149
transform 1 0 54832 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_589
timestamp 1644511149
transform 1 0 55292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_596
timestamp 1644511149
transform 1 0 55936 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_604
timestamp 1644511149
transform 1 0 56672 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_612
timestamp 1644511149
transform 1 0 57408 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_621
timestamp 1644511149
transform 1 0 58236 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 3680 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 13984 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 24288 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 29440 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 34592 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 39744 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 44896 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 50048 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 55200 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _064_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 38640 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _065_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19780 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _066_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _068_
timestamp 1644511149
transform 1 0 16008 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1644511149
transform 1 0 17388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _070_
timestamp 1644511149
transform 1 0 17480 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1644511149
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _072_
timestamp 1644511149
transform 1 0 18952 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1644511149
transform 1 0 19596 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 1644511149
transform 1 0 20148 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1644511149
transform 1 0 20792 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _076_
timestamp 1644511149
transform 1 0 26404 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _077_
timestamp 1644511149
transform 1 0 22172 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1644511149
transform 1 0 22448 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _079_
timestamp 1644511149
transform 1 0 23184 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _081_
timestamp 1644511149
transform 1 0 24564 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1644511149
transform 1 0 25760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _083_
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _084_
timestamp 1644511149
transform 1 0 26772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _085_
timestamp 1644511149
transform 1 0 27140 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _086_
timestamp 1644511149
transform 1 0 27876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _087_
timestamp 1644511149
transform 1 0 30820 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _088_
timestamp 1644511149
transform 1 0 29440 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp 1644511149
transform 1 0 30084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp 1644511149
transform 1 0 30636 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1644511149
transform 1 0 31096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _092_
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _093_
timestamp 1644511149
transform 1 0 32476 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _094_
timestamp 1644511149
transform 1 0 33304 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _095_
timestamp 1644511149
transform 1 0 33948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _096_
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1644511149
transform 1 0 35052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1644511149
transform 1 0 38088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _099_
timestamp 1644511149
transform 1 0 36064 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _100_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _101_
timestamp 1644511149
transform 1 0 37444 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _102_
timestamp 1644511149
transform 1 0 38180 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _103_
timestamp 1644511149
transform 1 0 38916 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _104_
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _105_
timestamp 1644511149
transform 1 0 41124 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _106_
timestamp 1644511149
transform 1 0 41032 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _107_
timestamp 1644511149
transform 1 0 41492 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _108_
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1644511149
transform 1 0 44804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _110_
timestamp 1644511149
transform 1 0 43608 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _111_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44344 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _112_
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1644511149
transform 1 0 46184 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _114_
timestamp 1644511149
transform 1 0 46000 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1644511149
transform 1 0 46736 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _116_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1644511149
transform 1 0 47932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _118_
timestamp 1644511149
transform 1 0 48576 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1644511149
transform 1 0 55660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _121_
timestamp 1644511149
transform 1 0 50784 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1644511149
transform 1 0 51520 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _123_
timestamp 1644511149
transform 1 0 51980 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _125_
timestamp 1644511149
transform 1 0 53176 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _127_
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _129_
timestamp 1644511149
transform 1 0 56488 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1644511149
transform 1 0 55200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _131_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _132_
timestamp 1644511149
transform 1 0 57132 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1644511149
transform 1 0 53176 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 1644511149
transform 1 0 56580 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1644511149
transform 1 0 57224 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1644511149
transform 1 0 6164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _137_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _138_
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _139_
timestamp 1644511149
transform 1 0 3496 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _140_
timestamp 1644511149
transform 1 0 4232 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _141_
timestamp 1644511149
transform 1 0 4508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _142_
timestamp 1644511149
transform 1 0 4784 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _143_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _144_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _145_
timestamp 1644511149
transform 1 0 6808 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _146_
timestamp 1644511149
transform 1 0 7636 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1644511149
transform 1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _148_
timestamp 1644511149
transform 1 0 9384 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1644511149
transform 1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _150_
timestamp 1644511149
transform 1 0 10488 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1644511149
transform 1 0 10580 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _152_
timestamp 1644511149
transform 1 0 12052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1644511149
transform 1 0 12052 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _154_
timestamp 1644511149
transform 1 0 12972 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _156_
timestamp 1644511149
transform 1 0 9384 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _157_
timestamp 1644511149
transform 1 0 9108 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1644511149
transform 1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _159_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _161_
timestamp 1644511149
transform 1 0 2852 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1644511149
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _163_
timestamp 1644511149
transform 1 0 4692 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _165_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _167_
timestamp 1644511149
transform 1 0 7268 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1644511149
transform 1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1644511149
transform 1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _170_
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _172_
timestamp 1644511149
transform 1 0 10488 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1644511149
transform 1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _174_
timestamp 1644511149
transform 1 0 12052 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _175_
timestamp 1644511149
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _176_
timestamp 1644511149
transform 1 0 12880 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _177_
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _178_
timestamp 1644511149
transform 1 0 9568 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _179_
timestamp 1644511149
transform 1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 56856 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1644511149
transform 1 0 56856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 55476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1644511149
transform 1 0 55476 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1644511149
transform 1 0 55936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1644511149
transform 1 0 57684 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1644511149
transform 1 0 56856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1644511149
transform 1 0 56764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input11
timestamp 1644511149
transform 1 0 54280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1644511149
transform 1 0 29532 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1644511149
transform 1 0 30728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1644511149
transform 1 0 33580 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1644511149
transform 1 0 34960 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1644511149
transform 1 0 36432 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1644511149
transform 1 0 37812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1644511149
transform 1 0 39836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 40664 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1644511149
transform 1 0 44988 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 46368 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 49220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1644511149
transform 1 0 50692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform 1 0 53544 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1644511149
transform 1 0 54556 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1644511149
transform 1 0 56396 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1644511149
transform 1 0 17848 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1644511149
transform 1 0 56580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1644511149
transform 1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1644511149
transform 1 0 20700 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 22080 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1644511149
transform 1 0 23552 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1644511149
transform 1 0 24932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1644511149
transform 1 0 27784 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 14996 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 33580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 36432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 40664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform 1 0 46368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 47840 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1644511149
transform 1 0 49220 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1644511149
transform 1 0 50692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1644511149
transform 1 0 53544 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1644511149
transform 1 0 56396 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1644511149
transform 1 0 57316 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1644511149
transform 1 0 57316 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1644511149
transform 1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1644511149
transform 1 0 27784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 2116 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 3772 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 4968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 6440 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 7820 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 10672 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 12144 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 2760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 57868 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 57868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 57868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 57868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 57868 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 57868 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 57868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1644511149
transform 1 0 57040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1644511149
transform 1 0 57868 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1644511149
transform 1 0 57040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1644511149
transform 1 0 56304 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1644511149
transform 1 0 55568 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1644511149
transform 1 0 55844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1644511149
transform 1 0 54464 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1644511149
transform 1 0 57868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1644511149
transform 1 0 57868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1644511149
transform 1 0 57868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1644511149
transform 1 0 57040 0 -1 10880
box -38 -48 406 592
<< labels >>
rlabel metal3 s 59200 552 60000 672 6 addr[0]
port 0 nsew signal input
rlabel metal3 s 59200 1096 60000 1216 6 addr[1]
port 1 nsew signal input
rlabel metal3 s 59200 1640 60000 1760 6 addr[2]
port 2 nsew signal input
rlabel metal3 s 59200 2184 60000 2304 6 addr[3]
port 3 nsew signal input
rlabel metal3 s 59200 2592 60000 2712 6 addr[4]
port 4 nsew signal input
rlabel metal3 s 59200 3136 60000 3256 6 addr[5]
port 5 nsew signal input
rlabel metal3 s 59200 3680 60000 3800 6 addr[6]
port 6 nsew signal input
rlabel metal3 s 59200 4224 60000 4344 6 addr[7]
port 7 nsew signal input
rlabel metal3 s 59200 4632 60000 4752 6 addr[8]
port 8 nsew signal input
rlabel metal3 s 59200 5176 60000 5296 6 addr[9]
port 9 nsew signal input
rlabel metal2 s 2042 21200 2098 22000 6 addr_mem0[0]
port 10 nsew signal tristate
rlabel metal2 s 3514 21200 3570 22000 6 addr_mem0[1]
port 11 nsew signal tristate
rlabel metal2 s 4894 21200 4950 22000 6 addr_mem0[2]
port 12 nsew signal tristate
rlabel metal2 s 6366 21200 6422 22000 6 addr_mem0[3]
port 13 nsew signal tristate
rlabel metal2 s 7746 21200 7802 22000 6 addr_mem0[4]
port 14 nsew signal tristate
rlabel metal2 s 9218 21200 9274 22000 6 addr_mem0[5]
port 15 nsew signal tristate
rlabel metal2 s 10598 21200 10654 22000 6 addr_mem0[6]
port 16 nsew signal tristate
rlabel metal2 s 12070 21200 12126 22000 6 addr_mem0[7]
port 17 nsew signal tristate
rlabel metal2 s 13450 21200 13506 22000 6 addr_mem0[8]
port 18 nsew signal tristate
rlabel metal2 s 2042 0 2098 800 6 addr_mem1[0]
port 19 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 addr_mem1[1]
port 20 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 addr_mem1[2]
port 21 nsew signal tristate
rlabel metal2 s 6366 0 6422 800 6 addr_mem1[3]
port 22 nsew signal tristate
rlabel metal2 s 7746 0 7802 800 6 addr_mem1[4]
port 23 nsew signal tristate
rlabel metal2 s 9218 0 9274 800 6 addr_mem1[5]
port 24 nsew signal tristate
rlabel metal2 s 10598 0 10654 800 6 addr_mem1[6]
port 25 nsew signal tristate
rlabel metal2 s 12070 0 12126 800 6 addr_mem1[7]
port 26 nsew signal tristate
rlabel metal2 s 13450 0 13506 800 6 addr_mem1[8]
port 27 nsew signal tristate
rlabel metal3 s 59200 144 60000 264 6 csb
port 28 nsew signal input
rlabel metal2 s 662 21200 718 22000 6 csb_mem0
port 29 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 csb_mem1
port 30 nsew signal tristate
rlabel metal3 s 59200 5720 60000 5840 6 dout[0]
port 31 nsew signal tristate
rlabel metal3 s 59200 10888 60000 11008 6 dout[10]
port 32 nsew signal tristate
rlabel metal3 s 59200 11296 60000 11416 6 dout[11]
port 33 nsew signal tristate
rlabel metal3 s 59200 11840 60000 11960 6 dout[12]
port 34 nsew signal tristate
rlabel metal3 s 59200 12384 60000 12504 6 dout[13]
port 35 nsew signal tristate
rlabel metal3 s 59200 12928 60000 13048 6 dout[14]
port 36 nsew signal tristate
rlabel metal3 s 59200 13336 60000 13456 6 dout[15]
port 37 nsew signal tristate
rlabel metal3 s 59200 13880 60000 14000 6 dout[16]
port 38 nsew signal tristate
rlabel metal3 s 59200 14424 60000 14544 6 dout[17]
port 39 nsew signal tristate
rlabel metal3 s 59200 14968 60000 15088 6 dout[18]
port 40 nsew signal tristate
rlabel metal3 s 59200 15512 60000 15632 6 dout[19]
port 41 nsew signal tristate
rlabel metal3 s 59200 6264 60000 6384 6 dout[1]
port 42 nsew signal tristate
rlabel metal3 s 59200 15920 60000 16040 6 dout[20]
port 43 nsew signal tristate
rlabel metal3 s 59200 16464 60000 16584 6 dout[21]
port 44 nsew signal tristate
rlabel metal3 s 59200 17008 60000 17128 6 dout[22]
port 45 nsew signal tristate
rlabel metal3 s 59200 17552 60000 17672 6 dout[23]
port 46 nsew signal tristate
rlabel metal3 s 59200 17960 60000 18080 6 dout[24]
port 47 nsew signal tristate
rlabel metal3 s 59200 18504 60000 18624 6 dout[25]
port 48 nsew signal tristate
rlabel metal3 s 59200 19048 60000 19168 6 dout[26]
port 49 nsew signal tristate
rlabel metal3 s 59200 19592 60000 19712 6 dout[27]
port 50 nsew signal tristate
rlabel metal3 s 59200 20000 60000 20120 6 dout[28]
port 51 nsew signal tristate
rlabel metal3 s 59200 20544 60000 20664 6 dout[29]
port 52 nsew signal tristate
rlabel metal3 s 59200 6672 60000 6792 6 dout[2]
port 53 nsew signal tristate
rlabel metal3 s 59200 21088 60000 21208 6 dout[30]
port 54 nsew signal tristate
rlabel metal3 s 59200 21632 60000 21752 6 dout[31]
port 55 nsew signal tristate
rlabel metal3 s 59200 7216 60000 7336 6 dout[3]
port 56 nsew signal tristate
rlabel metal3 s 59200 7760 60000 7880 6 dout[4]
port 57 nsew signal tristate
rlabel metal3 s 59200 8304 60000 8424 6 dout[5]
port 58 nsew signal tristate
rlabel metal3 s 59200 8848 60000 8968 6 dout[6]
port 59 nsew signal tristate
rlabel metal3 s 59200 9256 60000 9376 6 dout[7]
port 60 nsew signal tristate
rlabel metal3 s 59200 9800 60000 9920 6 dout[8]
port 61 nsew signal tristate
rlabel metal3 s 59200 10344 60000 10464 6 dout[9]
port 62 nsew signal tristate
rlabel metal2 s 14922 21200 14978 22000 6 dout_mem0[0]
port 63 nsew signal input
rlabel metal2 s 29182 21200 29238 22000 6 dout_mem0[10]
port 64 nsew signal input
rlabel metal2 s 30654 21200 30710 22000 6 dout_mem0[11]
port 65 nsew signal input
rlabel metal2 s 32034 21200 32090 22000 6 dout_mem0[12]
port 66 nsew signal input
rlabel metal2 s 33506 21200 33562 22000 6 dout_mem0[13]
port 67 nsew signal input
rlabel metal2 s 34886 21200 34942 22000 6 dout_mem0[14]
port 68 nsew signal input
rlabel metal2 s 36358 21200 36414 22000 6 dout_mem0[15]
port 69 nsew signal input
rlabel metal2 s 37738 21200 37794 22000 6 dout_mem0[16]
port 70 nsew signal input
rlabel metal2 s 39210 21200 39266 22000 6 dout_mem0[17]
port 71 nsew signal input
rlabel metal2 s 40590 21200 40646 22000 6 dout_mem0[18]
port 72 nsew signal input
rlabel metal2 s 42062 21200 42118 22000 6 dout_mem0[19]
port 73 nsew signal input
rlabel metal2 s 16302 21200 16358 22000 6 dout_mem0[1]
port 74 nsew signal input
rlabel metal2 s 43442 21200 43498 22000 6 dout_mem0[20]
port 75 nsew signal input
rlabel metal2 s 44914 21200 44970 22000 6 dout_mem0[21]
port 76 nsew signal input
rlabel metal2 s 46294 21200 46350 22000 6 dout_mem0[22]
port 77 nsew signal input
rlabel metal2 s 47766 21200 47822 22000 6 dout_mem0[23]
port 78 nsew signal input
rlabel metal2 s 49146 21200 49202 22000 6 dout_mem0[24]
port 79 nsew signal input
rlabel metal2 s 50618 21200 50674 22000 6 dout_mem0[25]
port 80 nsew signal input
rlabel metal2 s 51998 21200 52054 22000 6 dout_mem0[26]
port 81 nsew signal input
rlabel metal2 s 53470 21200 53526 22000 6 dout_mem0[27]
port 82 nsew signal input
rlabel metal2 s 54850 21200 54906 22000 6 dout_mem0[28]
port 83 nsew signal input
rlabel metal2 s 56322 21200 56378 22000 6 dout_mem0[29]
port 84 nsew signal input
rlabel metal2 s 17774 21200 17830 22000 6 dout_mem0[2]
port 85 nsew signal input
rlabel metal2 s 57702 21200 57758 22000 6 dout_mem0[30]
port 86 nsew signal input
rlabel metal2 s 59174 21200 59230 22000 6 dout_mem0[31]
port 87 nsew signal input
rlabel metal2 s 19154 21200 19210 22000 6 dout_mem0[3]
port 88 nsew signal input
rlabel metal2 s 20626 21200 20682 22000 6 dout_mem0[4]
port 89 nsew signal input
rlabel metal2 s 22006 21200 22062 22000 6 dout_mem0[5]
port 90 nsew signal input
rlabel metal2 s 23478 21200 23534 22000 6 dout_mem0[6]
port 91 nsew signal input
rlabel metal2 s 24858 21200 24914 22000 6 dout_mem0[7]
port 92 nsew signal input
rlabel metal2 s 26330 21200 26386 22000 6 dout_mem0[8]
port 93 nsew signal input
rlabel metal2 s 27710 21200 27766 22000 6 dout_mem0[9]
port 94 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 dout_mem1[0]
port 95 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 dout_mem1[10]
port 96 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 dout_mem1[11]
port 97 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 dout_mem1[12]
port 98 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 dout_mem1[13]
port 99 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 dout_mem1[14]
port 100 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 dout_mem1[15]
port 101 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 dout_mem1[16]
port 102 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 dout_mem1[17]
port 103 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 dout_mem1[18]
port 104 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 dout_mem1[19]
port 105 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 dout_mem1[1]
port 106 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 dout_mem1[20]
port 107 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 dout_mem1[21]
port 108 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 dout_mem1[22]
port 109 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 dout_mem1[23]
port 110 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 dout_mem1[24]
port 111 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 dout_mem1[25]
port 112 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 dout_mem1[26]
port 113 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 dout_mem1[27]
port 114 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 dout_mem1[28]
port 115 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 dout_mem1[29]
port 116 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 dout_mem1[2]
port 117 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 dout_mem1[30]
port 118 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 dout_mem1[31]
port 119 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 dout_mem1[3]
port 120 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 dout_mem1[4]
port 121 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 dout_mem1[5]
port 122 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 dout_mem1[6]
port 123 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 dout_mem1[7]
port 124 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 dout_mem1[8]
port 125 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 dout_mem1[9]
port 126 nsew signal input
rlabel metal4 s 10576 2128 10896 19632 6 vccd1
port 127 nsew power input
rlabel metal4 s 29840 2128 30160 19632 6 vccd1
port 127 nsew power input
rlabel metal4 s 49104 2128 49424 19632 6 vccd1
port 127 nsew power input
rlabel metal4 s 20208 2128 20528 19632 6 vssd1
port 128 nsew ground input
rlabel metal4 s 39472 2128 39792 19632 6 vssd1
port 128 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 60000 22000
<< end >>
