VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_memory
  CLASS BLOCK ;
  FOREIGN wb_memory ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 350.000 ;
  PIN addr_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 346.000 22.910 350.000 ;
    END
  END addr_mem0[0]
  PIN addr_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 346.000 41.310 350.000 ;
    END
  END addr_mem0[1]
  PIN addr_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 346.000 59.710 350.000 ;
    END
  END addr_mem0[2]
  PIN addr_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 346.000 78.110 350.000 ;
    END
  END addr_mem0[3]
  PIN addr_mem0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 346.000 96.510 350.000 ;
    END
  END addr_mem0[4]
  PIN addr_mem0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 346.000 110.310 350.000 ;
    END
  END addr_mem0[5]
  PIN addr_mem0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 346.000 124.110 350.000 ;
    END
  END addr_mem0[6]
  PIN addr_mem0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 346.000 137.910 350.000 ;
    END
  END addr_mem0[7]
  PIN addr_mem0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 346.000 151.710 350.000 ;
    END
  END addr_mem0[8]
  PIN addr_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 346.000 386.310 350.000 ;
    END
  END addr_mem1[0]
  PIN addr_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 346.000 404.710 350.000 ;
    END
  END addr_mem1[1]
  PIN addr_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 346.000 423.110 350.000 ;
    END
  END addr_mem1[2]
  PIN addr_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 346.000 441.510 350.000 ;
    END
  END addr_mem1[3]
  PIN addr_mem1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 346.000 459.910 350.000 ;
    END
  END addr_mem1[4]
  PIN addr_mem1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 346.000 473.710 350.000 ;
    END
  END addr_mem1[5]
  PIN addr_mem1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 346.000 487.510 350.000 ;
    END
  END addr_mem1[6]
  PIN addr_mem1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 346.000 501.310 350.000 ;
    END
  END addr_mem1[7]
  PIN addr_mem1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 346.000 515.110 350.000 ;
    END
  END addr_mem1[8]
  PIN csb_mem0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 346.000 13.710 350.000 ;
    END
  END csb_mem0
  PIN csb_mem1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 346.000 377.110 350.000 ;
    END
  END csb_mem1
  PIN din_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 346.000 27.510 350.000 ;
    END
  END din_mem0[0]
  PIN din_mem0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 346.000 174.710 350.000 ;
    END
  END din_mem0[10]
  PIN din_mem0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 346.000 183.910 350.000 ;
    END
  END din_mem0[11]
  PIN din_mem0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 346.000 193.110 350.000 ;
    END
  END din_mem0[12]
  PIN din_mem0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 346.000 202.310 350.000 ;
    END
  END din_mem0[13]
  PIN din_mem0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 346.000 211.510 350.000 ;
    END
  END din_mem0[14]
  PIN din_mem0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 346.000 220.710 350.000 ;
    END
  END din_mem0[15]
  PIN din_mem0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 346.000 229.910 350.000 ;
    END
  END din_mem0[16]
  PIN din_mem0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 346.000 239.110 350.000 ;
    END
  END din_mem0[17]
  PIN din_mem0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 346.000 248.310 350.000 ;
    END
  END din_mem0[18]
  PIN din_mem0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 346.000 257.510 350.000 ;
    END
  END din_mem0[19]
  PIN din_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 346.000 45.910 350.000 ;
    END
  END din_mem0[1]
  PIN din_mem0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 346.000 266.710 350.000 ;
    END
  END din_mem0[20]
  PIN din_mem0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 346.000 275.910 350.000 ;
    END
  END din_mem0[21]
  PIN din_mem0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 346.000 285.110 350.000 ;
    END
  END din_mem0[22]
  PIN din_mem0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 346.000 294.310 350.000 ;
    END
  END din_mem0[23]
  PIN din_mem0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 346.000 303.510 350.000 ;
    END
  END din_mem0[24]
  PIN din_mem0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 346.000 312.710 350.000 ;
    END
  END din_mem0[25]
  PIN din_mem0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 346.000 321.910 350.000 ;
    END
  END din_mem0[26]
  PIN din_mem0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 346.000 331.110 350.000 ;
    END
  END din_mem0[27]
  PIN din_mem0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 346.000 340.310 350.000 ;
    END
  END din_mem0[28]
  PIN din_mem0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 346.000 349.510 350.000 ;
    END
  END din_mem0[29]
  PIN din_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 346.000 64.310 350.000 ;
    END
  END din_mem0[2]
  PIN din_mem0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 346.000 358.710 350.000 ;
    END
  END din_mem0[30]
  PIN din_mem0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 346.000 367.910 350.000 ;
    END
  END din_mem0[31]
  PIN din_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 346.000 82.710 350.000 ;
    END
  END din_mem0[3]
  PIN din_mem0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 346.000 101.110 350.000 ;
    END
  END din_mem0[4]
  PIN din_mem0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 346.000 114.910 350.000 ;
    END
  END din_mem0[5]
  PIN din_mem0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 346.000 128.710 350.000 ;
    END
  END din_mem0[6]
  PIN din_mem0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 346.000 142.510 350.000 ;
    END
  END din_mem0[7]
  PIN din_mem0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 346.000 156.310 350.000 ;
    END
  END din_mem0[8]
  PIN din_mem0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 346.000 165.510 350.000 ;
    END
  END din_mem0[9]
  PIN din_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 346.000 390.910 350.000 ;
    END
  END din_mem1[0]
  PIN din_mem1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 346.000 538.110 350.000 ;
    END
  END din_mem1[10]
  PIN din_mem1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 346.000 547.310 350.000 ;
    END
  END din_mem1[11]
  PIN din_mem1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 346.000 556.510 350.000 ;
    END
  END din_mem1[12]
  PIN din_mem1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 346.000 565.710 350.000 ;
    END
  END din_mem1[13]
  PIN din_mem1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 346.000 574.910 350.000 ;
    END
  END din_mem1[14]
  PIN din_mem1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 346.000 584.110 350.000 ;
    END
  END din_mem1[15]
  PIN din_mem1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 346.000 593.310 350.000 ;
    END
  END din_mem1[16]
  PIN din_mem1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 346.000 602.510 350.000 ;
    END
  END din_mem1[17]
  PIN din_mem1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 346.000 611.710 350.000 ;
    END
  END din_mem1[18]
  PIN din_mem1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 346.000 620.910 350.000 ;
    END
  END din_mem1[19]
  PIN din_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 346.000 409.310 350.000 ;
    END
  END din_mem1[1]
  PIN din_mem1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 346.000 630.110 350.000 ;
    END
  END din_mem1[20]
  PIN din_mem1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 346.000 639.310 350.000 ;
    END
  END din_mem1[21]
  PIN din_mem1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 346.000 648.510 350.000 ;
    END
  END din_mem1[22]
  PIN din_mem1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 346.000 657.710 350.000 ;
    END
  END din_mem1[23]
  PIN din_mem1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 346.000 666.910 350.000 ;
    END
  END din_mem1[24]
  PIN din_mem1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 346.000 676.110 350.000 ;
    END
  END din_mem1[25]
  PIN din_mem1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 346.000 685.310 350.000 ;
    END
  END din_mem1[26]
  PIN din_mem1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 346.000 694.510 350.000 ;
    END
  END din_mem1[27]
  PIN din_mem1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 346.000 703.710 350.000 ;
    END
  END din_mem1[28]
  PIN din_mem1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 346.000 712.910 350.000 ;
    END
  END din_mem1[29]
  PIN din_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 346.000 427.710 350.000 ;
    END
  END din_mem1[2]
  PIN din_mem1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 346.000 722.110 350.000 ;
    END
  END din_mem1[30]
  PIN din_mem1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 346.000 731.310 350.000 ;
    END
  END din_mem1[31]
  PIN din_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 346.000 446.110 350.000 ;
    END
  END din_mem1[3]
  PIN din_mem1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 346.000 464.510 350.000 ;
    END
  END din_mem1[4]
  PIN din_mem1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 346.000 478.310 350.000 ;
    END
  END din_mem1[5]
  PIN din_mem1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 346.000 492.110 350.000 ;
    END
  END din_mem1[6]
  PIN din_mem1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 346.000 505.910 350.000 ;
    END
  END din_mem1[7]
  PIN din_mem1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 346.000 519.710 350.000 ;
    END
  END din_mem1[8]
  PIN din_mem1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 346.000 528.910 350.000 ;
    END
  END din_mem1[9]
  PIN dout_mem0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 346.000 32.110 350.000 ;
    END
  END dout_mem0[0]
  PIN dout_mem0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 346.000 179.310 350.000 ;
    END
  END dout_mem0[10]
  PIN dout_mem0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 346.000 188.510 350.000 ;
    END
  END dout_mem0[11]
  PIN dout_mem0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 346.000 197.710 350.000 ;
    END
  END dout_mem0[12]
  PIN dout_mem0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 346.000 206.910 350.000 ;
    END
  END dout_mem0[13]
  PIN dout_mem0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 346.000 216.110 350.000 ;
    END
  END dout_mem0[14]
  PIN dout_mem0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 346.000 225.310 350.000 ;
    END
  END dout_mem0[15]
  PIN dout_mem0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 346.000 234.510 350.000 ;
    END
  END dout_mem0[16]
  PIN dout_mem0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 346.000 243.710 350.000 ;
    END
  END dout_mem0[17]
  PIN dout_mem0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 346.000 252.910 350.000 ;
    END
  END dout_mem0[18]
  PIN dout_mem0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 346.000 262.110 350.000 ;
    END
  END dout_mem0[19]
  PIN dout_mem0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 346.000 50.510 350.000 ;
    END
  END dout_mem0[1]
  PIN dout_mem0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 346.000 271.310 350.000 ;
    END
  END dout_mem0[20]
  PIN dout_mem0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 346.000 280.510 350.000 ;
    END
  END dout_mem0[21]
  PIN dout_mem0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 346.000 289.710 350.000 ;
    END
  END dout_mem0[22]
  PIN dout_mem0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 346.000 298.910 350.000 ;
    END
  END dout_mem0[23]
  PIN dout_mem0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 346.000 308.110 350.000 ;
    END
  END dout_mem0[24]
  PIN dout_mem0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 346.000 317.310 350.000 ;
    END
  END dout_mem0[25]
  PIN dout_mem0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 346.000 326.510 350.000 ;
    END
  END dout_mem0[26]
  PIN dout_mem0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 346.000 335.710 350.000 ;
    END
  END dout_mem0[27]
  PIN dout_mem0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 346.000 344.910 350.000 ;
    END
  END dout_mem0[28]
  PIN dout_mem0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 346.000 354.110 350.000 ;
    END
  END dout_mem0[29]
  PIN dout_mem0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 346.000 68.910 350.000 ;
    END
  END dout_mem0[2]
  PIN dout_mem0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 346.000 363.310 350.000 ;
    END
  END dout_mem0[30]
  PIN dout_mem0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 346.000 372.510 350.000 ;
    END
  END dout_mem0[31]
  PIN dout_mem0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 346.000 87.310 350.000 ;
    END
  END dout_mem0[3]
  PIN dout_mem0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 346.000 105.710 350.000 ;
    END
  END dout_mem0[4]
  PIN dout_mem0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 346.000 119.510 350.000 ;
    END
  END dout_mem0[5]
  PIN dout_mem0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 346.000 133.310 350.000 ;
    END
  END dout_mem0[6]
  PIN dout_mem0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 346.000 147.110 350.000 ;
    END
  END dout_mem0[7]
  PIN dout_mem0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 346.000 160.910 350.000 ;
    END
  END dout_mem0[8]
  PIN dout_mem0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 346.000 170.110 350.000 ;
    END
  END dout_mem0[9]
  PIN dout_mem1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 346.000 395.510 350.000 ;
    END
  END dout_mem1[0]
  PIN dout_mem1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 346.000 542.710 350.000 ;
    END
  END dout_mem1[10]
  PIN dout_mem1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 346.000 551.910 350.000 ;
    END
  END dout_mem1[11]
  PIN dout_mem1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 346.000 561.110 350.000 ;
    END
  END dout_mem1[12]
  PIN dout_mem1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 346.000 570.310 350.000 ;
    END
  END dout_mem1[13]
  PIN dout_mem1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 346.000 579.510 350.000 ;
    END
  END dout_mem1[14]
  PIN dout_mem1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 346.000 588.710 350.000 ;
    END
  END dout_mem1[15]
  PIN dout_mem1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 346.000 597.910 350.000 ;
    END
  END dout_mem1[16]
  PIN dout_mem1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 346.000 607.110 350.000 ;
    END
  END dout_mem1[17]
  PIN dout_mem1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 346.000 616.310 350.000 ;
    END
  END dout_mem1[18]
  PIN dout_mem1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 346.000 625.510 350.000 ;
    END
  END dout_mem1[19]
  PIN dout_mem1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 346.000 413.910 350.000 ;
    END
  END dout_mem1[1]
  PIN dout_mem1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 346.000 634.710 350.000 ;
    END
  END dout_mem1[20]
  PIN dout_mem1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 346.000 643.910 350.000 ;
    END
  END dout_mem1[21]
  PIN dout_mem1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 346.000 653.110 350.000 ;
    END
  END dout_mem1[22]
  PIN dout_mem1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 346.000 662.310 350.000 ;
    END
  END dout_mem1[23]
  PIN dout_mem1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 346.000 671.510 350.000 ;
    END
  END dout_mem1[24]
  PIN dout_mem1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 346.000 680.710 350.000 ;
    END
  END dout_mem1[25]
  PIN dout_mem1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 346.000 689.910 350.000 ;
    END
  END dout_mem1[26]
  PIN dout_mem1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 346.000 699.110 350.000 ;
    END
  END dout_mem1[27]
  PIN dout_mem1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 346.000 708.310 350.000 ;
    END
  END dout_mem1[28]
  PIN dout_mem1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 346.000 717.510 350.000 ;
    END
  END dout_mem1[29]
  PIN dout_mem1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 346.000 432.310 350.000 ;
    END
  END dout_mem1[2]
  PIN dout_mem1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 346.000 726.710 350.000 ;
    END
  END dout_mem1[30]
  PIN dout_mem1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 346.000 735.910 350.000 ;
    END
  END dout_mem1[31]
  PIN dout_mem1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.430 346.000 450.710 350.000 ;
    END
  END dout_mem1[3]
  PIN dout_mem1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.830 346.000 469.110 350.000 ;
    END
  END dout_mem1[4]
  PIN dout_mem1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 346.000 482.910 350.000 ;
    END
  END dout_mem1[5]
  PIN dout_mem1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 346.000 496.710 350.000 ;
    END
  END dout_mem1[6]
  PIN dout_mem1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 346.000 510.510 350.000 ;
    END
  END dout_mem1[7]
  PIN dout_mem1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 346.000 524.310 350.000 ;
    END
  END dout_mem1[8]
  PIN dout_mem1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 346.000 533.510 350.000 ;
    END
  END dout_mem1[9]
  PIN io_wbs_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END io_wbs_ack
  PIN io_wbs_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END io_wbs_adr[0]
  PIN io_wbs_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END io_wbs_adr[10]
  PIN io_wbs_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END io_wbs_adr[11]
  PIN io_wbs_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END io_wbs_adr[12]
  PIN io_wbs_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END io_wbs_adr[13]
  PIN io_wbs_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END io_wbs_adr[14]
  PIN io_wbs_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END io_wbs_adr[15]
  PIN io_wbs_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END io_wbs_adr[16]
  PIN io_wbs_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END io_wbs_adr[17]
  PIN io_wbs_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END io_wbs_adr[18]
  PIN io_wbs_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END io_wbs_adr[19]
  PIN io_wbs_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END io_wbs_adr[1]
  PIN io_wbs_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END io_wbs_adr[20]
  PIN io_wbs_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END io_wbs_adr[21]
  PIN io_wbs_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END io_wbs_adr[22]
  PIN io_wbs_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END io_wbs_adr[23]
  PIN io_wbs_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END io_wbs_adr[24]
  PIN io_wbs_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END io_wbs_adr[25]
  PIN io_wbs_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END io_wbs_adr[26]
  PIN io_wbs_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END io_wbs_adr[27]
  PIN io_wbs_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END io_wbs_adr[28]
  PIN io_wbs_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END io_wbs_adr[29]
  PIN io_wbs_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END io_wbs_adr[2]
  PIN io_wbs_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END io_wbs_adr[30]
  PIN io_wbs_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END io_wbs_adr[31]
  PIN io_wbs_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END io_wbs_adr[3]
  PIN io_wbs_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_wbs_adr[4]
  PIN io_wbs_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END io_wbs_adr[5]
  PIN io_wbs_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END io_wbs_adr[6]
  PIN io_wbs_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END io_wbs_adr[7]
  PIN io_wbs_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END io_wbs_adr[8]
  PIN io_wbs_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END io_wbs_adr[9]
  PIN io_wbs_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END io_wbs_clk
  PIN io_wbs_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END io_wbs_cyc
  PIN io_wbs_datrd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END io_wbs_datrd[0]
  PIN io_wbs_datrd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END io_wbs_datrd[10]
  PIN io_wbs_datrd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END io_wbs_datrd[11]
  PIN io_wbs_datrd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END io_wbs_datrd[12]
  PIN io_wbs_datrd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END io_wbs_datrd[13]
  PIN io_wbs_datrd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END io_wbs_datrd[14]
  PIN io_wbs_datrd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END io_wbs_datrd[15]
  PIN io_wbs_datrd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END io_wbs_datrd[16]
  PIN io_wbs_datrd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END io_wbs_datrd[17]
  PIN io_wbs_datrd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END io_wbs_datrd[18]
  PIN io_wbs_datrd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END io_wbs_datrd[19]
  PIN io_wbs_datrd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END io_wbs_datrd[1]
  PIN io_wbs_datrd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END io_wbs_datrd[20]
  PIN io_wbs_datrd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END io_wbs_datrd[21]
  PIN io_wbs_datrd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END io_wbs_datrd[22]
  PIN io_wbs_datrd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END io_wbs_datrd[23]
  PIN io_wbs_datrd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END io_wbs_datrd[24]
  PIN io_wbs_datrd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 0.000 606.190 4.000 ;
    END
  END io_wbs_datrd[25]
  PIN io_wbs_datrd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END io_wbs_datrd[26]
  PIN io_wbs_datrd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END io_wbs_datrd[27]
  PIN io_wbs_datrd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END io_wbs_datrd[28]
  PIN io_wbs_datrd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END io_wbs_datrd[29]
  PIN io_wbs_datrd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END io_wbs_datrd[2]
  PIN io_wbs_datrd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END io_wbs_datrd[30]
  PIN io_wbs_datrd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END io_wbs_datrd[31]
  PIN io_wbs_datrd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END io_wbs_datrd[3]
  PIN io_wbs_datrd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END io_wbs_datrd[4]
  PIN io_wbs_datrd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END io_wbs_datrd[5]
  PIN io_wbs_datrd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END io_wbs_datrd[6]
  PIN io_wbs_datrd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END io_wbs_datrd[7]
  PIN io_wbs_datrd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END io_wbs_datrd[8]
  PIN io_wbs_datrd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END io_wbs_datrd[9]
  PIN io_wbs_datwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END io_wbs_datwr[0]
  PIN io_wbs_datwr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END io_wbs_datwr[10]
  PIN io_wbs_datwr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END io_wbs_datwr[11]
  PIN io_wbs_datwr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END io_wbs_datwr[12]
  PIN io_wbs_datwr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END io_wbs_datwr[13]
  PIN io_wbs_datwr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END io_wbs_datwr[14]
  PIN io_wbs_datwr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END io_wbs_datwr[15]
  PIN io_wbs_datwr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END io_wbs_datwr[16]
  PIN io_wbs_datwr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END io_wbs_datwr[17]
  PIN io_wbs_datwr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END io_wbs_datwr[18]
  PIN io_wbs_datwr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END io_wbs_datwr[19]
  PIN io_wbs_datwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END io_wbs_datwr[1]
  PIN io_wbs_datwr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END io_wbs_datwr[20]
  PIN io_wbs_datwr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END io_wbs_datwr[21]
  PIN io_wbs_datwr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END io_wbs_datwr[22]
  PIN io_wbs_datwr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END io_wbs_datwr[23]
  PIN io_wbs_datwr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END io_wbs_datwr[24]
  PIN io_wbs_datwr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END io_wbs_datwr[25]
  PIN io_wbs_datwr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END io_wbs_datwr[26]
  PIN io_wbs_datwr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.210 0.000 654.490 4.000 ;
    END
  END io_wbs_datwr[27]
  PIN io_wbs_datwr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END io_wbs_datwr[28]
  PIN io_wbs_datwr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END io_wbs_datwr[29]
  PIN io_wbs_datwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END io_wbs_datwr[2]
  PIN io_wbs_datwr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END io_wbs_datwr[30]
  PIN io_wbs_datwr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 0.000 737.290 4.000 ;
    END
  END io_wbs_datwr[31]
  PIN io_wbs_datwr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END io_wbs_datwr[3]
  PIN io_wbs_datwr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END io_wbs_datwr[4]
  PIN io_wbs_datwr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END io_wbs_datwr[5]
  PIN io_wbs_datwr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 4.000 ;
    END
  END io_wbs_datwr[6]
  PIN io_wbs_datwr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END io_wbs_datwr[7]
  PIN io_wbs_datwr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END io_wbs_datwr[8]
  PIN io_wbs_datwr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END io_wbs_datwr[9]
  PIN io_wbs_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END io_wbs_rst
  PIN io_wbs_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END io_wbs_sel[0]
  PIN io_wbs_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END io_wbs_sel[1]
  PIN io_wbs_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END io_wbs_sel[2]
  PIN io_wbs_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END io_wbs_sel[3]
  PIN io_wbs_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END io_wbs_stb
  PIN io_wbs_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END io_wbs_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 337.520 ;
    END
  END vssd1
  PIN web_mem0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 346.000 18.310 350.000 ;
    END
  END web_mem0
  PIN web_mem1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 346.000 381.710 350.000 ;
    END
  END web_mem1
  PIN wmask_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 346.000 36.710 350.000 ;
    END
  END wmask_mem0[0]
  PIN wmask_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 346.000 55.110 350.000 ;
    END
  END wmask_mem0[1]
  PIN wmask_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 346.000 73.510 350.000 ;
    END
  END wmask_mem0[2]
  PIN wmask_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 346.000 91.910 350.000 ;
    END
  END wmask_mem0[3]
  PIN wmask_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 346.000 400.110 350.000 ;
    END
  END wmask_mem1[0]
  PIN wmask_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 346.000 418.510 350.000 ;
    END
  END wmask_mem1[1]
  PIN wmask_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 346.000 436.910 350.000 ;
    END
  END wmask_mem1[2]
  PIN wmask_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 346.000 455.310 350.000 ;
    END
  END wmask_mem1[3]
  OBS
      LAYER nwell ;
        RECT 5.330 333.145 744.470 335.975 ;
        RECT 5.330 327.705 744.470 330.535 ;
        RECT 5.330 322.265 744.470 325.095 ;
        RECT 5.330 316.825 744.470 319.655 ;
        RECT 5.330 311.385 744.470 314.215 ;
        RECT 5.330 305.945 744.470 308.775 ;
        RECT 5.330 300.505 744.470 303.335 ;
        RECT 5.330 295.065 744.470 297.895 ;
        RECT 5.330 289.625 744.470 292.455 ;
        RECT 5.330 284.185 744.470 287.015 ;
        RECT 5.330 278.745 744.470 281.575 ;
        RECT 5.330 273.305 744.470 276.135 ;
        RECT 5.330 267.865 744.470 270.695 ;
        RECT 5.330 262.425 744.470 265.255 ;
        RECT 5.330 256.985 744.470 259.815 ;
        RECT 5.330 251.545 744.470 254.375 ;
        RECT 5.330 246.105 744.470 248.935 ;
        RECT 5.330 240.665 744.470 243.495 ;
        RECT 5.330 235.225 744.470 238.055 ;
        RECT 5.330 229.785 744.470 232.615 ;
        RECT 5.330 224.345 744.470 227.175 ;
        RECT 5.330 218.905 744.470 221.735 ;
        RECT 5.330 213.465 744.470 216.295 ;
        RECT 5.330 208.025 744.470 210.855 ;
        RECT 5.330 202.585 744.470 205.415 ;
        RECT 5.330 197.145 744.470 199.975 ;
        RECT 5.330 191.705 744.470 194.535 ;
        RECT 5.330 186.265 744.470 189.095 ;
        RECT 5.330 180.825 744.470 183.655 ;
        RECT 5.330 175.385 744.470 178.215 ;
        RECT 5.330 169.945 744.470 172.775 ;
        RECT 5.330 164.505 744.470 167.335 ;
        RECT 5.330 159.065 744.470 161.895 ;
        RECT 5.330 153.625 744.470 156.455 ;
        RECT 5.330 148.185 744.470 151.015 ;
        RECT 5.330 142.745 744.470 145.575 ;
        RECT 5.330 137.305 744.470 140.135 ;
        RECT 5.330 131.865 744.470 134.695 ;
        RECT 5.330 126.425 744.470 129.255 ;
        RECT 5.330 120.985 744.470 123.815 ;
        RECT 5.330 115.545 744.470 118.375 ;
        RECT 5.330 110.105 744.470 112.935 ;
        RECT 5.330 104.665 744.470 107.495 ;
        RECT 5.330 99.225 744.470 102.055 ;
        RECT 5.330 93.785 744.470 96.615 ;
        RECT 5.330 88.345 744.470 91.175 ;
        RECT 5.330 82.905 744.470 85.735 ;
        RECT 5.330 77.465 744.470 80.295 ;
        RECT 5.330 72.025 744.470 74.855 ;
        RECT 5.330 66.585 744.470 69.415 ;
        RECT 5.330 61.145 744.470 63.975 ;
        RECT 5.330 55.705 744.470 58.535 ;
        RECT 5.330 50.265 744.470 53.095 ;
        RECT 5.330 44.825 744.470 47.655 ;
        RECT 5.330 39.385 744.470 42.215 ;
        RECT 5.330 33.945 744.470 36.775 ;
        RECT 5.330 28.505 744.470 31.335 ;
        RECT 5.330 23.065 744.470 25.895 ;
        RECT 5.330 17.625 744.470 20.455 ;
        RECT 5.330 12.185 744.470 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 744.280 337.365 ;
      LAYER met1 ;
        RECT 5.520 8.540 744.280 348.460 ;
      LAYER met2 ;
        RECT 12.520 345.720 13.150 348.490 ;
        RECT 13.990 345.720 17.750 348.490 ;
        RECT 18.590 345.720 22.350 348.490 ;
        RECT 23.190 345.720 26.950 348.490 ;
        RECT 27.790 345.720 31.550 348.490 ;
        RECT 32.390 345.720 36.150 348.490 ;
        RECT 36.990 345.720 40.750 348.490 ;
        RECT 41.590 345.720 45.350 348.490 ;
        RECT 46.190 345.720 49.950 348.490 ;
        RECT 50.790 345.720 54.550 348.490 ;
        RECT 55.390 345.720 59.150 348.490 ;
        RECT 59.990 345.720 63.750 348.490 ;
        RECT 64.590 345.720 68.350 348.490 ;
        RECT 69.190 345.720 72.950 348.490 ;
        RECT 73.790 345.720 77.550 348.490 ;
        RECT 78.390 345.720 82.150 348.490 ;
        RECT 82.990 345.720 86.750 348.490 ;
        RECT 87.590 345.720 91.350 348.490 ;
        RECT 92.190 345.720 95.950 348.490 ;
        RECT 96.790 345.720 100.550 348.490 ;
        RECT 101.390 345.720 105.150 348.490 ;
        RECT 105.990 345.720 109.750 348.490 ;
        RECT 110.590 345.720 114.350 348.490 ;
        RECT 115.190 345.720 118.950 348.490 ;
        RECT 119.790 345.720 123.550 348.490 ;
        RECT 124.390 345.720 128.150 348.490 ;
        RECT 128.990 345.720 132.750 348.490 ;
        RECT 133.590 345.720 137.350 348.490 ;
        RECT 138.190 345.720 141.950 348.490 ;
        RECT 142.790 345.720 146.550 348.490 ;
        RECT 147.390 345.720 151.150 348.490 ;
        RECT 151.990 345.720 155.750 348.490 ;
        RECT 156.590 345.720 160.350 348.490 ;
        RECT 161.190 345.720 164.950 348.490 ;
        RECT 165.790 345.720 169.550 348.490 ;
        RECT 170.390 345.720 174.150 348.490 ;
        RECT 174.990 345.720 178.750 348.490 ;
        RECT 179.590 345.720 183.350 348.490 ;
        RECT 184.190 345.720 187.950 348.490 ;
        RECT 188.790 345.720 192.550 348.490 ;
        RECT 193.390 345.720 197.150 348.490 ;
        RECT 197.990 345.720 201.750 348.490 ;
        RECT 202.590 345.720 206.350 348.490 ;
        RECT 207.190 345.720 210.950 348.490 ;
        RECT 211.790 345.720 215.550 348.490 ;
        RECT 216.390 345.720 220.150 348.490 ;
        RECT 220.990 345.720 224.750 348.490 ;
        RECT 225.590 345.720 229.350 348.490 ;
        RECT 230.190 345.720 233.950 348.490 ;
        RECT 234.790 345.720 238.550 348.490 ;
        RECT 239.390 345.720 243.150 348.490 ;
        RECT 243.990 345.720 247.750 348.490 ;
        RECT 248.590 345.720 252.350 348.490 ;
        RECT 253.190 345.720 256.950 348.490 ;
        RECT 257.790 345.720 261.550 348.490 ;
        RECT 262.390 345.720 266.150 348.490 ;
        RECT 266.990 345.720 270.750 348.490 ;
        RECT 271.590 345.720 275.350 348.490 ;
        RECT 276.190 345.720 279.950 348.490 ;
        RECT 280.790 345.720 284.550 348.490 ;
        RECT 285.390 345.720 289.150 348.490 ;
        RECT 289.990 345.720 293.750 348.490 ;
        RECT 294.590 345.720 298.350 348.490 ;
        RECT 299.190 345.720 302.950 348.490 ;
        RECT 303.790 345.720 307.550 348.490 ;
        RECT 308.390 345.720 312.150 348.490 ;
        RECT 312.990 345.720 316.750 348.490 ;
        RECT 317.590 345.720 321.350 348.490 ;
        RECT 322.190 345.720 325.950 348.490 ;
        RECT 326.790 345.720 330.550 348.490 ;
        RECT 331.390 345.720 335.150 348.490 ;
        RECT 335.990 345.720 339.750 348.490 ;
        RECT 340.590 345.720 344.350 348.490 ;
        RECT 345.190 345.720 348.950 348.490 ;
        RECT 349.790 345.720 353.550 348.490 ;
        RECT 354.390 345.720 358.150 348.490 ;
        RECT 358.990 345.720 362.750 348.490 ;
        RECT 363.590 345.720 367.350 348.490 ;
        RECT 368.190 345.720 371.950 348.490 ;
        RECT 372.790 345.720 376.550 348.490 ;
        RECT 377.390 345.720 381.150 348.490 ;
        RECT 381.990 345.720 385.750 348.490 ;
        RECT 386.590 345.720 390.350 348.490 ;
        RECT 391.190 345.720 394.950 348.490 ;
        RECT 395.790 345.720 399.550 348.490 ;
        RECT 400.390 345.720 404.150 348.490 ;
        RECT 404.990 345.720 408.750 348.490 ;
        RECT 409.590 345.720 413.350 348.490 ;
        RECT 414.190 345.720 417.950 348.490 ;
        RECT 418.790 345.720 422.550 348.490 ;
        RECT 423.390 345.720 427.150 348.490 ;
        RECT 427.990 345.720 431.750 348.490 ;
        RECT 432.590 345.720 436.350 348.490 ;
        RECT 437.190 345.720 440.950 348.490 ;
        RECT 441.790 345.720 445.550 348.490 ;
        RECT 446.390 345.720 450.150 348.490 ;
        RECT 450.990 345.720 454.750 348.490 ;
        RECT 455.590 345.720 459.350 348.490 ;
        RECT 460.190 345.720 463.950 348.490 ;
        RECT 464.790 345.720 468.550 348.490 ;
        RECT 469.390 345.720 473.150 348.490 ;
        RECT 473.990 345.720 477.750 348.490 ;
        RECT 478.590 345.720 482.350 348.490 ;
        RECT 483.190 345.720 486.950 348.490 ;
        RECT 487.790 345.720 491.550 348.490 ;
        RECT 492.390 345.720 496.150 348.490 ;
        RECT 496.990 345.720 500.750 348.490 ;
        RECT 501.590 345.720 505.350 348.490 ;
        RECT 506.190 345.720 509.950 348.490 ;
        RECT 510.790 345.720 514.550 348.490 ;
        RECT 515.390 345.720 519.150 348.490 ;
        RECT 519.990 345.720 523.750 348.490 ;
        RECT 524.590 345.720 528.350 348.490 ;
        RECT 529.190 345.720 532.950 348.490 ;
        RECT 533.790 345.720 537.550 348.490 ;
        RECT 538.390 345.720 542.150 348.490 ;
        RECT 542.990 345.720 546.750 348.490 ;
        RECT 547.590 345.720 551.350 348.490 ;
        RECT 552.190 345.720 555.950 348.490 ;
        RECT 556.790 345.720 560.550 348.490 ;
        RECT 561.390 345.720 565.150 348.490 ;
        RECT 565.990 345.720 569.750 348.490 ;
        RECT 570.590 345.720 574.350 348.490 ;
        RECT 575.190 345.720 578.950 348.490 ;
        RECT 579.790 345.720 583.550 348.490 ;
        RECT 584.390 345.720 588.150 348.490 ;
        RECT 588.990 345.720 592.750 348.490 ;
        RECT 593.590 345.720 597.350 348.490 ;
        RECT 598.190 345.720 601.950 348.490 ;
        RECT 602.790 345.720 606.550 348.490 ;
        RECT 607.390 345.720 611.150 348.490 ;
        RECT 611.990 345.720 615.750 348.490 ;
        RECT 616.590 345.720 620.350 348.490 ;
        RECT 621.190 345.720 624.950 348.490 ;
        RECT 625.790 345.720 629.550 348.490 ;
        RECT 630.390 345.720 634.150 348.490 ;
        RECT 634.990 345.720 638.750 348.490 ;
        RECT 639.590 345.720 643.350 348.490 ;
        RECT 644.190 345.720 647.950 348.490 ;
        RECT 648.790 345.720 652.550 348.490 ;
        RECT 653.390 345.720 657.150 348.490 ;
        RECT 657.990 345.720 661.750 348.490 ;
        RECT 662.590 345.720 666.350 348.490 ;
        RECT 667.190 345.720 670.950 348.490 ;
        RECT 671.790 345.720 675.550 348.490 ;
        RECT 676.390 345.720 680.150 348.490 ;
        RECT 680.990 345.720 684.750 348.490 ;
        RECT 685.590 345.720 689.350 348.490 ;
        RECT 690.190 345.720 693.950 348.490 ;
        RECT 694.790 345.720 698.550 348.490 ;
        RECT 699.390 345.720 703.150 348.490 ;
        RECT 703.990 345.720 707.750 348.490 ;
        RECT 708.590 345.720 712.350 348.490 ;
        RECT 713.190 345.720 716.950 348.490 ;
        RECT 717.790 345.720 721.550 348.490 ;
        RECT 722.390 345.720 726.150 348.490 ;
        RECT 726.990 345.720 730.750 348.490 ;
        RECT 731.590 345.720 735.350 348.490 ;
        RECT 736.190 345.720 737.290 348.490 ;
        RECT 12.520 4.280 737.290 345.720 ;
        RECT 13.070 3.670 19.130 4.280 ;
        RECT 19.970 3.670 26.030 4.280 ;
        RECT 26.870 3.670 32.930 4.280 ;
        RECT 33.770 3.670 39.830 4.280 ;
        RECT 40.670 3.670 46.730 4.280 ;
        RECT 47.570 3.670 53.630 4.280 ;
        RECT 54.470 3.670 60.530 4.280 ;
        RECT 61.370 3.670 67.430 4.280 ;
        RECT 68.270 3.670 74.330 4.280 ;
        RECT 75.170 3.670 81.230 4.280 ;
        RECT 82.070 3.670 88.130 4.280 ;
        RECT 88.970 3.670 95.030 4.280 ;
        RECT 95.870 3.670 101.930 4.280 ;
        RECT 102.770 3.670 108.830 4.280 ;
        RECT 109.670 3.670 115.730 4.280 ;
        RECT 116.570 3.670 122.630 4.280 ;
        RECT 123.470 3.670 129.530 4.280 ;
        RECT 130.370 3.670 136.430 4.280 ;
        RECT 137.270 3.670 143.330 4.280 ;
        RECT 144.170 3.670 150.230 4.280 ;
        RECT 151.070 3.670 157.130 4.280 ;
        RECT 157.970 3.670 164.030 4.280 ;
        RECT 164.870 3.670 170.930 4.280 ;
        RECT 171.770 3.670 177.830 4.280 ;
        RECT 178.670 3.670 184.730 4.280 ;
        RECT 185.570 3.670 191.630 4.280 ;
        RECT 192.470 3.670 198.530 4.280 ;
        RECT 199.370 3.670 205.430 4.280 ;
        RECT 206.270 3.670 212.330 4.280 ;
        RECT 213.170 3.670 219.230 4.280 ;
        RECT 220.070 3.670 226.130 4.280 ;
        RECT 226.970 3.670 233.030 4.280 ;
        RECT 233.870 3.670 239.930 4.280 ;
        RECT 240.770 3.670 246.830 4.280 ;
        RECT 247.670 3.670 253.730 4.280 ;
        RECT 254.570 3.670 260.630 4.280 ;
        RECT 261.470 3.670 267.530 4.280 ;
        RECT 268.370 3.670 274.430 4.280 ;
        RECT 275.270 3.670 281.330 4.280 ;
        RECT 282.170 3.670 288.230 4.280 ;
        RECT 289.070 3.670 295.130 4.280 ;
        RECT 295.970 3.670 302.030 4.280 ;
        RECT 302.870 3.670 308.930 4.280 ;
        RECT 309.770 3.670 315.830 4.280 ;
        RECT 316.670 3.670 322.730 4.280 ;
        RECT 323.570 3.670 329.630 4.280 ;
        RECT 330.470 3.670 336.530 4.280 ;
        RECT 337.370 3.670 343.430 4.280 ;
        RECT 344.270 3.670 350.330 4.280 ;
        RECT 351.170 3.670 357.230 4.280 ;
        RECT 358.070 3.670 364.130 4.280 ;
        RECT 364.970 3.670 371.030 4.280 ;
        RECT 371.870 3.670 377.930 4.280 ;
        RECT 378.770 3.670 384.830 4.280 ;
        RECT 385.670 3.670 391.730 4.280 ;
        RECT 392.570 3.670 398.630 4.280 ;
        RECT 399.470 3.670 405.530 4.280 ;
        RECT 406.370 3.670 412.430 4.280 ;
        RECT 413.270 3.670 419.330 4.280 ;
        RECT 420.170 3.670 426.230 4.280 ;
        RECT 427.070 3.670 433.130 4.280 ;
        RECT 433.970 3.670 440.030 4.280 ;
        RECT 440.870 3.670 446.930 4.280 ;
        RECT 447.770 3.670 453.830 4.280 ;
        RECT 454.670 3.670 460.730 4.280 ;
        RECT 461.570 3.670 467.630 4.280 ;
        RECT 468.470 3.670 474.530 4.280 ;
        RECT 475.370 3.670 481.430 4.280 ;
        RECT 482.270 3.670 488.330 4.280 ;
        RECT 489.170 3.670 495.230 4.280 ;
        RECT 496.070 3.670 502.130 4.280 ;
        RECT 502.970 3.670 509.030 4.280 ;
        RECT 509.870 3.670 515.930 4.280 ;
        RECT 516.770 3.670 522.830 4.280 ;
        RECT 523.670 3.670 529.730 4.280 ;
        RECT 530.570 3.670 536.630 4.280 ;
        RECT 537.470 3.670 543.530 4.280 ;
        RECT 544.370 3.670 550.430 4.280 ;
        RECT 551.270 3.670 557.330 4.280 ;
        RECT 558.170 3.670 564.230 4.280 ;
        RECT 565.070 3.670 571.130 4.280 ;
        RECT 571.970 3.670 578.030 4.280 ;
        RECT 578.870 3.670 584.930 4.280 ;
        RECT 585.770 3.670 591.830 4.280 ;
        RECT 592.670 3.670 598.730 4.280 ;
        RECT 599.570 3.670 605.630 4.280 ;
        RECT 606.470 3.670 612.530 4.280 ;
        RECT 613.370 3.670 619.430 4.280 ;
        RECT 620.270 3.670 626.330 4.280 ;
        RECT 627.170 3.670 633.230 4.280 ;
        RECT 634.070 3.670 640.130 4.280 ;
        RECT 640.970 3.670 647.030 4.280 ;
        RECT 647.870 3.670 653.930 4.280 ;
        RECT 654.770 3.670 660.830 4.280 ;
        RECT 661.670 3.670 667.730 4.280 ;
        RECT 668.570 3.670 674.630 4.280 ;
        RECT 675.470 3.670 681.530 4.280 ;
        RECT 682.370 3.670 688.430 4.280 ;
        RECT 689.270 3.670 695.330 4.280 ;
        RECT 696.170 3.670 702.230 4.280 ;
        RECT 703.070 3.670 709.130 4.280 ;
        RECT 709.970 3.670 716.030 4.280 ;
        RECT 716.870 3.670 722.930 4.280 ;
        RECT 723.770 3.670 729.830 4.280 ;
        RECT 730.670 3.670 736.730 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 737.315 339.145 ;
  END
END wb_memory
END LIBRARY

