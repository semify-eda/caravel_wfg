magic
tech sky130A
magscale 1 2
timestamp 1657004107
<< obsli1 >>
rect 1104 2159 58880 19601
<< obsm1 >>
rect 658 2128 59234 19848
<< metal2 >>
rect 662 21200 718 22000
rect 2042 21200 2098 22000
rect 3514 21200 3570 22000
rect 4894 21200 4950 22000
rect 6366 21200 6422 22000
rect 7746 21200 7802 22000
rect 9218 21200 9274 22000
rect 10598 21200 10654 22000
rect 12070 21200 12126 22000
rect 13450 21200 13506 22000
rect 14922 21200 14978 22000
rect 16302 21200 16358 22000
rect 17774 21200 17830 22000
rect 19154 21200 19210 22000
rect 20626 21200 20682 22000
rect 22006 21200 22062 22000
rect 23478 21200 23534 22000
rect 24858 21200 24914 22000
rect 26330 21200 26386 22000
rect 27710 21200 27766 22000
rect 29182 21200 29238 22000
rect 30654 21200 30710 22000
rect 32034 21200 32090 22000
rect 33506 21200 33562 22000
rect 34886 21200 34942 22000
rect 36358 21200 36414 22000
rect 37738 21200 37794 22000
rect 39210 21200 39266 22000
rect 40590 21200 40646 22000
rect 42062 21200 42118 22000
rect 43442 21200 43498 22000
rect 44914 21200 44970 22000
rect 46294 21200 46350 22000
rect 47766 21200 47822 22000
rect 49146 21200 49202 22000
rect 50618 21200 50674 22000
rect 51998 21200 52054 22000
rect 53470 21200 53526 22000
rect 54850 21200 54906 22000
rect 56322 21200 56378 22000
rect 57702 21200 57758 22000
rect 59174 21200 59230 22000
rect 662 0 718 800
rect 2042 0 2098 800
rect 3514 0 3570 800
rect 4894 0 4950 800
rect 6366 0 6422 800
rect 7746 0 7802 800
rect 9218 0 9274 800
rect 10598 0 10654 800
rect 12070 0 12126 800
rect 13450 0 13506 800
rect 14922 0 14978 800
rect 16302 0 16358 800
rect 17774 0 17830 800
rect 19154 0 19210 800
rect 20626 0 20682 800
rect 22006 0 22062 800
rect 23478 0 23534 800
rect 24858 0 24914 800
rect 26330 0 26386 800
rect 27710 0 27766 800
rect 29182 0 29238 800
rect 30654 0 30710 800
rect 32034 0 32090 800
rect 33506 0 33562 800
rect 34886 0 34942 800
rect 36358 0 36414 800
rect 37738 0 37794 800
rect 39210 0 39266 800
rect 40590 0 40646 800
rect 42062 0 42118 800
rect 43442 0 43498 800
rect 44914 0 44970 800
rect 46294 0 46350 800
rect 47766 0 47822 800
rect 49146 0 49202 800
rect 50618 0 50674 800
rect 51998 0 52054 800
rect 53470 0 53526 800
rect 54850 0 54906 800
rect 56322 0 56378 800
rect 57702 0 57758 800
rect 59174 0 59230 800
<< obsm2 >>
rect 774 21144 1986 21729
rect 2154 21144 3458 21729
rect 3626 21144 4838 21729
rect 5006 21144 6310 21729
rect 6478 21144 7690 21729
rect 7858 21144 9162 21729
rect 9330 21144 10542 21729
rect 10710 21144 12014 21729
rect 12182 21144 13394 21729
rect 13562 21144 14866 21729
rect 15034 21144 16246 21729
rect 16414 21144 17718 21729
rect 17886 21144 19098 21729
rect 19266 21144 20570 21729
rect 20738 21144 21950 21729
rect 22118 21144 23422 21729
rect 23590 21144 24802 21729
rect 24970 21144 26274 21729
rect 26442 21144 27654 21729
rect 27822 21144 29126 21729
rect 29294 21144 30598 21729
rect 30766 21144 31978 21729
rect 32146 21144 33450 21729
rect 33618 21144 34830 21729
rect 34998 21144 36302 21729
rect 36470 21144 37682 21729
rect 37850 21144 39154 21729
rect 39322 21144 40534 21729
rect 40702 21144 42006 21729
rect 42174 21144 43386 21729
rect 43554 21144 44858 21729
rect 45026 21144 46238 21729
rect 46406 21144 47710 21729
rect 47878 21144 49090 21729
rect 49258 21144 50562 21729
rect 50730 21144 51942 21729
rect 52110 21144 53414 21729
rect 53582 21144 54794 21729
rect 54962 21144 56266 21729
rect 56434 21144 57646 21729
rect 57814 21144 59118 21729
rect 664 856 59228 21144
rect 774 54 1986 856
rect 2154 54 3458 856
rect 3626 54 4838 856
rect 5006 54 6310 856
rect 6478 54 7690 856
rect 7858 54 9162 856
rect 9330 54 10542 856
rect 10710 54 12014 856
rect 12182 54 13394 856
rect 13562 54 14866 856
rect 15034 54 16246 856
rect 16414 54 17718 856
rect 17886 54 19098 856
rect 19266 54 20570 856
rect 20738 54 21950 856
rect 22118 54 23422 856
rect 23590 54 24802 856
rect 24970 54 26274 856
rect 26442 54 27654 856
rect 27822 54 29126 856
rect 29294 54 30598 856
rect 30766 54 31978 856
rect 32146 54 33450 856
rect 33618 54 34830 856
rect 34998 54 36302 856
rect 36470 54 37682 856
rect 37850 54 39154 856
rect 39322 54 40534 856
rect 40702 54 42006 856
rect 42174 54 43386 856
rect 43554 54 44858 856
rect 45026 54 46238 856
rect 46406 54 47710 856
rect 47878 54 49090 856
rect 49258 54 50562 856
rect 50730 54 51942 856
rect 52110 54 53414 856
rect 53582 54 54794 856
rect 54962 54 56266 856
rect 56434 54 57646 856
rect 57814 54 59118 856
<< metal3 >>
rect 59200 21632 60000 21752
rect 59200 21088 60000 21208
rect 59200 20544 60000 20664
rect 59200 20000 60000 20120
rect 59200 19592 60000 19712
rect 59200 19048 60000 19168
rect 59200 18504 60000 18624
rect 59200 17960 60000 18080
rect 59200 17552 60000 17672
rect 59200 17008 60000 17128
rect 59200 16464 60000 16584
rect 59200 15920 60000 16040
rect 59200 15512 60000 15632
rect 59200 14968 60000 15088
rect 59200 14424 60000 14544
rect 59200 13880 60000 14000
rect 59200 13336 60000 13456
rect 59200 12928 60000 13048
rect 59200 12384 60000 12504
rect 59200 11840 60000 11960
rect 59200 11296 60000 11416
rect 59200 10888 60000 11008
rect 59200 10344 60000 10464
rect 59200 9800 60000 9920
rect 59200 9256 60000 9376
rect 59200 8848 60000 8968
rect 59200 8304 60000 8424
rect 59200 7760 60000 7880
rect 59200 7216 60000 7336
rect 59200 6672 60000 6792
rect 59200 6264 60000 6384
rect 59200 5720 60000 5840
rect 59200 5176 60000 5296
rect 59200 4632 60000 4752
rect 59200 4224 60000 4344
rect 59200 3680 60000 3800
rect 59200 3136 60000 3256
rect 59200 2592 60000 2712
rect 59200 2184 60000 2304
rect 59200 1640 60000 1760
rect 59200 1096 60000 1216
rect 59200 552 60000 672
rect 59200 144 60000 264
<< obsm3 >>
rect 10576 21552 59120 21725
rect 10576 21288 59200 21552
rect 10576 21008 59120 21288
rect 10576 20744 59200 21008
rect 10576 20464 59120 20744
rect 10576 20200 59200 20464
rect 10576 19920 59120 20200
rect 10576 19792 59200 19920
rect 10576 19512 59120 19792
rect 10576 19248 59200 19512
rect 10576 18968 59120 19248
rect 10576 18704 59200 18968
rect 10576 18424 59120 18704
rect 10576 18160 59200 18424
rect 10576 17880 59120 18160
rect 10576 17752 59200 17880
rect 10576 17472 59120 17752
rect 10576 17208 59200 17472
rect 10576 16928 59120 17208
rect 10576 16664 59200 16928
rect 10576 16384 59120 16664
rect 10576 16120 59200 16384
rect 10576 15840 59120 16120
rect 10576 15712 59200 15840
rect 10576 15432 59120 15712
rect 10576 15168 59200 15432
rect 10576 14888 59120 15168
rect 10576 14624 59200 14888
rect 10576 14344 59120 14624
rect 10576 14080 59200 14344
rect 10576 13800 59120 14080
rect 10576 13536 59200 13800
rect 10576 13256 59120 13536
rect 10576 13128 59200 13256
rect 10576 12848 59120 13128
rect 10576 12584 59200 12848
rect 10576 12304 59120 12584
rect 10576 12040 59200 12304
rect 10576 11760 59120 12040
rect 10576 11496 59200 11760
rect 10576 11216 59120 11496
rect 10576 11088 59200 11216
rect 10576 10808 59120 11088
rect 10576 10544 59200 10808
rect 10576 10264 59120 10544
rect 10576 10000 59200 10264
rect 10576 9720 59120 10000
rect 10576 9456 59200 9720
rect 10576 9176 59120 9456
rect 10576 9048 59200 9176
rect 10576 8768 59120 9048
rect 10576 8504 59200 8768
rect 10576 8224 59120 8504
rect 10576 7960 59200 8224
rect 10576 7680 59120 7960
rect 10576 7416 59200 7680
rect 10576 7136 59120 7416
rect 10576 6872 59200 7136
rect 10576 6592 59120 6872
rect 10576 6464 59200 6592
rect 10576 6184 59120 6464
rect 10576 5920 59200 6184
rect 10576 5640 59120 5920
rect 10576 5376 59200 5640
rect 10576 5096 59120 5376
rect 10576 4832 59200 5096
rect 10576 4552 59120 4832
rect 10576 4424 59200 4552
rect 10576 4144 59120 4424
rect 10576 3880 59200 4144
rect 10576 3600 59120 3880
rect 10576 3336 59200 3600
rect 10576 3056 59120 3336
rect 10576 2792 59200 3056
rect 10576 2512 59120 2792
rect 10576 2384 59200 2512
rect 10576 2104 59120 2384
rect 10576 1840 59200 2104
rect 10576 1560 59120 1840
rect 10576 1296 59200 1560
rect 10576 1016 59120 1296
rect 10576 752 59200 1016
rect 10576 472 59120 752
rect 10576 344 59200 472
rect 10576 171 59120 344
<< metal4 >>
rect 10576 2128 10896 19632
rect 20208 2128 20528 19632
rect 29840 2128 30160 19632
rect 39472 2128 39792 19632
rect 49104 2128 49424 19632
<< labels >>
rlabel metal3 s 59200 552 60000 672 6 addr[0]
port 1 nsew signal input
rlabel metal3 s 59200 1096 60000 1216 6 addr[1]
port 2 nsew signal input
rlabel metal3 s 59200 1640 60000 1760 6 addr[2]
port 3 nsew signal input
rlabel metal3 s 59200 2184 60000 2304 6 addr[3]
port 4 nsew signal input
rlabel metal3 s 59200 2592 60000 2712 6 addr[4]
port 5 nsew signal input
rlabel metal3 s 59200 3136 60000 3256 6 addr[5]
port 6 nsew signal input
rlabel metal3 s 59200 3680 60000 3800 6 addr[6]
port 7 nsew signal input
rlabel metal3 s 59200 4224 60000 4344 6 addr[7]
port 8 nsew signal input
rlabel metal3 s 59200 4632 60000 4752 6 addr[8]
port 9 nsew signal input
rlabel metal3 s 59200 5176 60000 5296 6 addr[9]
port 10 nsew signal input
rlabel metal2 s 2042 21200 2098 22000 6 addr_mem0[0]
port 11 nsew signal output
rlabel metal2 s 3514 21200 3570 22000 6 addr_mem0[1]
port 12 nsew signal output
rlabel metal2 s 4894 21200 4950 22000 6 addr_mem0[2]
port 13 nsew signal output
rlabel metal2 s 6366 21200 6422 22000 6 addr_mem0[3]
port 14 nsew signal output
rlabel metal2 s 7746 21200 7802 22000 6 addr_mem0[4]
port 15 nsew signal output
rlabel metal2 s 9218 21200 9274 22000 6 addr_mem0[5]
port 16 nsew signal output
rlabel metal2 s 10598 21200 10654 22000 6 addr_mem0[6]
port 17 nsew signal output
rlabel metal2 s 12070 21200 12126 22000 6 addr_mem0[7]
port 18 nsew signal output
rlabel metal2 s 13450 21200 13506 22000 6 addr_mem0[8]
port 19 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 addr_mem1[0]
port 20 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 addr_mem1[1]
port 21 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 addr_mem1[2]
port 22 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 addr_mem1[3]
port 23 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 addr_mem1[4]
port 24 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 addr_mem1[5]
port 25 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 addr_mem1[6]
port 26 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 addr_mem1[7]
port 27 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 addr_mem1[8]
port 28 nsew signal output
rlabel metal3 s 59200 144 60000 264 6 csb
port 29 nsew signal input
rlabel metal2 s 662 21200 718 22000 6 csb_mem0
port 30 nsew signal output
rlabel metal2 s 662 0 718 800 6 csb_mem1
port 31 nsew signal output
rlabel metal3 s 59200 5720 60000 5840 6 dout[0]
port 32 nsew signal output
rlabel metal3 s 59200 10888 60000 11008 6 dout[10]
port 33 nsew signal output
rlabel metal3 s 59200 11296 60000 11416 6 dout[11]
port 34 nsew signal output
rlabel metal3 s 59200 11840 60000 11960 6 dout[12]
port 35 nsew signal output
rlabel metal3 s 59200 12384 60000 12504 6 dout[13]
port 36 nsew signal output
rlabel metal3 s 59200 12928 60000 13048 6 dout[14]
port 37 nsew signal output
rlabel metal3 s 59200 13336 60000 13456 6 dout[15]
port 38 nsew signal output
rlabel metal3 s 59200 13880 60000 14000 6 dout[16]
port 39 nsew signal output
rlabel metal3 s 59200 14424 60000 14544 6 dout[17]
port 40 nsew signal output
rlabel metal3 s 59200 14968 60000 15088 6 dout[18]
port 41 nsew signal output
rlabel metal3 s 59200 15512 60000 15632 6 dout[19]
port 42 nsew signal output
rlabel metal3 s 59200 6264 60000 6384 6 dout[1]
port 43 nsew signal output
rlabel metal3 s 59200 15920 60000 16040 6 dout[20]
port 44 nsew signal output
rlabel metal3 s 59200 16464 60000 16584 6 dout[21]
port 45 nsew signal output
rlabel metal3 s 59200 17008 60000 17128 6 dout[22]
port 46 nsew signal output
rlabel metal3 s 59200 17552 60000 17672 6 dout[23]
port 47 nsew signal output
rlabel metal3 s 59200 17960 60000 18080 6 dout[24]
port 48 nsew signal output
rlabel metal3 s 59200 18504 60000 18624 6 dout[25]
port 49 nsew signal output
rlabel metal3 s 59200 19048 60000 19168 6 dout[26]
port 50 nsew signal output
rlabel metal3 s 59200 19592 60000 19712 6 dout[27]
port 51 nsew signal output
rlabel metal3 s 59200 20000 60000 20120 6 dout[28]
port 52 nsew signal output
rlabel metal3 s 59200 20544 60000 20664 6 dout[29]
port 53 nsew signal output
rlabel metal3 s 59200 6672 60000 6792 6 dout[2]
port 54 nsew signal output
rlabel metal3 s 59200 21088 60000 21208 6 dout[30]
port 55 nsew signal output
rlabel metal3 s 59200 21632 60000 21752 6 dout[31]
port 56 nsew signal output
rlabel metal3 s 59200 7216 60000 7336 6 dout[3]
port 57 nsew signal output
rlabel metal3 s 59200 7760 60000 7880 6 dout[4]
port 58 nsew signal output
rlabel metal3 s 59200 8304 60000 8424 6 dout[5]
port 59 nsew signal output
rlabel metal3 s 59200 8848 60000 8968 6 dout[6]
port 60 nsew signal output
rlabel metal3 s 59200 9256 60000 9376 6 dout[7]
port 61 nsew signal output
rlabel metal3 s 59200 9800 60000 9920 6 dout[8]
port 62 nsew signal output
rlabel metal3 s 59200 10344 60000 10464 6 dout[9]
port 63 nsew signal output
rlabel metal2 s 14922 21200 14978 22000 6 dout_mem0[0]
port 64 nsew signal input
rlabel metal2 s 29182 21200 29238 22000 6 dout_mem0[10]
port 65 nsew signal input
rlabel metal2 s 30654 21200 30710 22000 6 dout_mem0[11]
port 66 nsew signal input
rlabel metal2 s 32034 21200 32090 22000 6 dout_mem0[12]
port 67 nsew signal input
rlabel metal2 s 33506 21200 33562 22000 6 dout_mem0[13]
port 68 nsew signal input
rlabel metal2 s 34886 21200 34942 22000 6 dout_mem0[14]
port 69 nsew signal input
rlabel metal2 s 36358 21200 36414 22000 6 dout_mem0[15]
port 70 nsew signal input
rlabel metal2 s 37738 21200 37794 22000 6 dout_mem0[16]
port 71 nsew signal input
rlabel metal2 s 39210 21200 39266 22000 6 dout_mem0[17]
port 72 nsew signal input
rlabel metal2 s 40590 21200 40646 22000 6 dout_mem0[18]
port 73 nsew signal input
rlabel metal2 s 42062 21200 42118 22000 6 dout_mem0[19]
port 74 nsew signal input
rlabel metal2 s 16302 21200 16358 22000 6 dout_mem0[1]
port 75 nsew signal input
rlabel metal2 s 43442 21200 43498 22000 6 dout_mem0[20]
port 76 nsew signal input
rlabel metal2 s 44914 21200 44970 22000 6 dout_mem0[21]
port 77 nsew signal input
rlabel metal2 s 46294 21200 46350 22000 6 dout_mem0[22]
port 78 nsew signal input
rlabel metal2 s 47766 21200 47822 22000 6 dout_mem0[23]
port 79 nsew signal input
rlabel metal2 s 49146 21200 49202 22000 6 dout_mem0[24]
port 80 nsew signal input
rlabel metal2 s 50618 21200 50674 22000 6 dout_mem0[25]
port 81 nsew signal input
rlabel metal2 s 51998 21200 52054 22000 6 dout_mem0[26]
port 82 nsew signal input
rlabel metal2 s 53470 21200 53526 22000 6 dout_mem0[27]
port 83 nsew signal input
rlabel metal2 s 54850 21200 54906 22000 6 dout_mem0[28]
port 84 nsew signal input
rlabel metal2 s 56322 21200 56378 22000 6 dout_mem0[29]
port 85 nsew signal input
rlabel metal2 s 17774 21200 17830 22000 6 dout_mem0[2]
port 86 nsew signal input
rlabel metal2 s 57702 21200 57758 22000 6 dout_mem0[30]
port 87 nsew signal input
rlabel metal2 s 59174 21200 59230 22000 6 dout_mem0[31]
port 88 nsew signal input
rlabel metal2 s 19154 21200 19210 22000 6 dout_mem0[3]
port 89 nsew signal input
rlabel metal2 s 20626 21200 20682 22000 6 dout_mem0[4]
port 90 nsew signal input
rlabel metal2 s 22006 21200 22062 22000 6 dout_mem0[5]
port 91 nsew signal input
rlabel metal2 s 23478 21200 23534 22000 6 dout_mem0[6]
port 92 nsew signal input
rlabel metal2 s 24858 21200 24914 22000 6 dout_mem0[7]
port 93 nsew signal input
rlabel metal2 s 26330 21200 26386 22000 6 dout_mem0[8]
port 94 nsew signal input
rlabel metal2 s 27710 21200 27766 22000 6 dout_mem0[9]
port 95 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 dout_mem1[0]
port 96 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 dout_mem1[10]
port 97 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 dout_mem1[11]
port 98 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 dout_mem1[12]
port 99 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 dout_mem1[13]
port 100 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 dout_mem1[14]
port 101 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 dout_mem1[15]
port 102 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 dout_mem1[16]
port 103 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 dout_mem1[17]
port 104 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 dout_mem1[18]
port 105 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 dout_mem1[19]
port 106 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 dout_mem1[1]
port 107 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 dout_mem1[20]
port 108 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 dout_mem1[21]
port 109 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 dout_mem1[22]
port 110 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 dout_mem1[23]
port 111 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 dout_mem1[24]
port 112 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 dout_mem1[25]
port 113 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 dout_mem1[26]
port 114 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 dout_mem1[27]
port 115 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 dout_mem1[28]
port 116 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 dout_mem1[29]
port 117 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 dout_mem1[2]
port 118 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 dout_mem1[30]
port 119 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 dout_mem1[31]
port 120 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 dout_mem1[3]
port 121 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 dout_mem1[4]
port 122 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 dout_mem1[5]
port 123 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 dout_mem1[6]
port 124 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 dout_mem1[7]
port 125 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 dout_mem1[8]
port 126 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 dout_mem1[9]
port 127 nsew signal input
rlabel metal4 s 10576 2128 10896 19632 6 vccd1
port 128 nsew power input
rlabel metal4 s 29840 2128 30160 19632 6 vccd1
port 128 nsew power input
rlabel metal4 s 49104 2128 49424 19632 6 vccd1
port 128 nsew power input
rlabel metal4 s 20208 2128 20528 19632 6 vssd1
port 129 nsew ground input
rlabel metal4 s 39472 2128 39792 19632 6 vssd1
port 129 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 60000 22000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 741482
string GDS_FILE /home/leo/Dokumente/caravel_workspace/caravel_wfg/openlane/merge_memory/runs/merge_memory/results/finishing/merge_memory.magic.gds
string GDS_START 72906
<< end >>

