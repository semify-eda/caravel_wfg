magic
tech sky130A
magscale 1 2
timestamp 1657184941
<< viali >>
rect 117329 37417 117363 37451
rect 118065 37417 118099 37451
rect 117145 37213 117179 37247
rect 117881 37213 117915 37247
rect 117329 36873 117363 36907
rect 117145 36737 117179 36771
rect 117881 36737 117915 36771
rect 118065 36601 118099 36635
rect 117881 36125 117915 36159
rect 118065 35989 118099 36023
rect 117881 35037 117915 35071
rect 118065 34901 118099 34935
rect 117881 33949 117915 33983
rect 118065 33813 118099 33847
rect 117881 33473 117915 33507
rect 118065 33269 118099 33303
rect 117881 32385 117915 32419
rect 118065 32181 118099 32215
rect 117881 31297 117915 31331
rect 118065 31093 118099 31127
rect 117881 30209 117915 30243
rect 118065 30073 118099 30107
rect 117881 29597 117915 29631
rect 118065 29461 118099 29495
rect 117881 28509 117915 28543
rect 118065 28373 118099 28407
rect 117881 27421 117915 27455
rect 118065 27285 118099 27319
rect 117881 26945 117915 26979
rect 118065 26741 118099 26775
rect 117513 25857 117547 25891
rect 117881 25857 117915 25891
rect 118065 25653 118099 25687
rect 117513 24769 117547 24803
rect 117881 24769 117915 24803
rect 118065 24565 118099 24599
rect 117513 23681 117547 23715
rect 117881 23681 117915 23715
rect 118065 23545 118099 23579
rect 117513 23069 117547 23103
rect 117881 23069 117915 23103
rect 118065 22933 118099 22967
rect 117881 21981 117915 22015
rect 117513 21845 117547 21879
rect 118065 21845 118099 21879
rect 117513 20893 117547 20927
rect 117881 20893 117915 20927
rect 118065 20757 118099 20791
rect 117513 20417 117547 20451
rect 117881 20417 117915 20451
rect 118065 20213 118099 20247
rect 117881 19329 117915 19363
rect 117513 19125 117547 19159
rect 118065 19125 118099 19159
rect 117881 18241 117915 18275
rect 117513 18037 117547 18071
rect 118065 18037 118099 18071
rect 117513 17629 117547 17663
rect 117881 17629 117915 17663
rect 118065 17493 118099 17527
rect 117881 16541 117915 16575
rect 117513 16405 117547 16439
rect 118065 16405 118099 16439
rect 117513 15453 117547 15487
rect 117881 15453 117915 15487
rect 118065 15317 118099 15351
rect 117513 14365 117547 14399
rect 117881 14365 117915 14399
rect 118065 14229 118099 14263
rect 117513 13889 117547 13923
rect 117881 13889 117915 13923
rect 118065 13685 118099 13719
rect 89453 12937 89487 12971
rect 89269 12801 89303 12835
rect 117513 12801 117547 12835
rect 117881 12801 117915 12835
rect 118065 12597 118099 12631
rect 117881 11713 117915 11747
rect 118065 11577 118099 11611
rect 117513 11509 117547 11543
rect 118065 11237 118099 11271
rect 117513 11101 117547 11135
rect 117881 11101 117915 11135
rect 76113 10217 76147 10251
rect 75929 10013 75963 10047
rect 117789 9945 117823 9979
rect 117881 9877 117915 9911
rect 117789 8857 117823 8891
rect 117881 8789 117915 8823
rect 117789 7769 117823 7803
rect 117881 7701 117915 7735
rect 117789 7361 117823 7395
rect 117881 7157 117915 7191
rect 91017 6409 91051 6443
rect 88809 6273 88843 6307
rect 90833 6273 90867 6307
rect 117789 6273 117823 6307
rect 88993 6069 89027 6103
rect 117881 6069 117915 6103
rect 117973 5661 118007 5695
rect 117789 5525 117823 5559
rect 117789 5185 117823 5219
rect 117881 4981 117915 5015
rect 116409 4777 116443 4811
rect 116225 4573 116259 4607
rect 117789 4505 117823 4539
rect 117881 4437 117915 4471
rect 97825 4233 97859 4267
rect 100677 4233 100711 4267
rect 117789 4165 117823 4199
rect 98009 4097 98043 4131
rect 100861 4097 100895 4131
rect 115121 4097 115155 4131
rect 115857 4097 115891 4131
rect 116593 4097 116627 4131
rect 117973 3961 118007 3995
rect 114937 3893 114971 3927
rect 116041 3893 116075 3927
rect 116777 3893 116811 3927
rect 117881 3689 117915 3723
rect 99021 3621 99055 3655
rect 106013 3621 106047 3655
rect 114937 3621 114971 3655
rect 115765 3621 115799 3655
rect 116409 3553 116443 3587
rect 63141 3485 63175 3519
rect 68385 3485 68419 3519
rect 68845 3485 68879 3519
rect 76573 3485 76607 3519
rect 82277 3485 82311 3519
rect 83749 3485 83783 3519
rect 85129 3485 85163 3519
rect 86601 3485 86635 3519
rect 87981 3485 88015 3519
rect 91753 3485 91787 3519
rect 92213 3485 92247 3519
rect 96721 3485 96755 3519
rect 97917 3485 97951 3519
rect 99665 3485 99699 3519
rect 100401 3485 100435 3519
rect 105829 3485 105863 3519
rect 107025 3485 107059 3519
rect 112269 3485 112303 3519
rect 114753 3485 114787 3519
rect 115121 3485 115155 3519
rect 116133 3485 116167 3519
rect 116225 3485 116259 3519
rect 98837 3417 98871 3451
rect 117789 3417 117823 3451
rect 62957 3349 62991 3383
rect 68661 3349 68695 3383
rect 76389 3349 76423 3383
rect 82093 3349 82127 3383
rect 83565 3349 83599 3383
rect 84945 3349 84979 3383
rect 86417 3349 86451 3383
rect 87797 3349 87831 3383
rect 91569 3349 91603 3383
rect 92397 3349 92431 3383
rect 96537 3349 96571 3383
rect 98101 3349 98135 3383
rect 99849 3349 99883 3383
rect 100585 3349 100619 3383
rect 106841 3349 106875 3383
rect 112085 3349 112119 3383
rect 115305 3349 115339 3383
rect 65809 3145 65843 3179
rect 76665 3145 76699 3179
rect 78689 3145 78723 3179
rect 79609 3145 79643 3179
rect 81725 3145 81759 3179
rect 82829 3145 82863 3179
rect 85221 3145 85255 3179
rect 86693 3145 86727 3179
rect 92673 3145 92707 3179
rect 95985 3145 96019 3179
rect 96721 3145 96755 3179
rect 99113 3145 99147 3179
rect 99573 3145 99607 3179
rect 101045 3145 101079 3179
rect 102425 3145 102459 3179
rect 104449 3145 104483 3179
rect 106105 3145 106139 3179
rect 107025 3145 107059 3179
rect 108497 3145 108531 3179
rect 110797 3145 110831 3179
rect 111901 3145 111935 3179
rect 115121 3145 115155 3179
rect 115489 3145 115523 3179
rect 115857 3145 115891 3179
rect 116317 3145 116351 3179
rect 117053 3145 117087 3179
rect 87521 3077 87555 3111
rect 88901 3077 88935 3111
rect 109785 3077 109819 3111
rect 110429 3077 110463 3111
rect 116869 3077 116903 3111
rect 55413 3009 55447 3043
rect 59277 3009 59311 3043
rect 60289 3009 60323 3043
rect 60749 3009 60783 3043
rect 61669 3009 61703 3043
rect 63601 3009 63635 3043
rect 64889 3009 64923 3043
rect 65993 3009 66027 3043
rect 66269 3009 66303 3043
rect 66913 3009 66947 3043
rect 67373 3009 67407 3043
rect 68201 3009 68235 3043
rect 69121 3009 69155 3043
rect 70225 3009 70259 3043
rect 70685 3009 70719 3043
rect 71697 3009 71731 3043
rect 72157 3009 72191 3043
rect 73537 3009 73571 3043
rect 75193 3009 75227 3043
rect 76573 3009 76607 3043
rect 77953 3009 77987 3043
rect 78597 3009 78631 3043
rect 79517 3009 79551 3043
rect 80897 3009 80931 3043
rect 81633 3009 81667 3043
rect 82553 3009 82587 3043
rect 83749 3009 83783 3043
rect 85129 3009 85163 3043
rect 86601 3009 86635 3043
rect 89729 3009 89763 3043
rect 90925 3009 90959 3043
rect 92581 3009 92615 3043
rect 95157 3009 95191 3043
rect 95801 3009 95835 3043
rect 96537 3009 96571 3043
rect 97641 3009 97675 3043
rect 98285 3009 98319 3043
rect 99481 3009 99515 3043
rect 100125 3009 100159 3043
rect 100401 3009 100435 3043
rect 101229 3009 101263 3043
rect 102241 3009 102275 3043
rect 103161 3009 103195 3043
rect 104265 3009 104299 3043
rect 105001 3009 105035 3043
rect 105369 3009 105403 3043
rect 106013 3009 106047 3043
rect 106841 3009 106875 3043
rect 107853 3009 107887 3043
rect 108313 3009 108347 3043
rect 109877 3009 109911 3043
rect 110613 3009 110647 3043
rect 111717 3009 111751 3043
rect 112545 3009 112579 3043
rect 113741 3009 113775 3043
rect 116225 3009 116259 3043
rect 117237 3009 117271 3043
rect 117789 3009 117823 3043
rect 65533 2941 65567 2975
rect 84025 2941 84059 2975
rect 89085 2941 89119 2975
rect 92765 2941 92799 2975
rect 93225 2941 93259 2975
rect 99757 2941 99791 2975
rect 106197 2941 106231 2975
rect 109969 2941 110003 2975
rect 116409 2941 116443 2975
rect 60105 2873 60139 2907
rect 67189 2873 67223 2907
rect 70041 2873 70075 2907
rect 71513 2873 71547 2907
rect 105645 2873 105679 2907
rect 109417 2873 109451 2907
rect 55689 2805 55723 2839
rect 59461 2805 59495 2839
rect 60933 2805 60967 2839
rect 61485 2805 61519 2839
rect 63785 2805 63819 2839
rect 65073 2805 65107 2839
rect 66453 2805 66487 2839
rect 68385 2805 68419 2839
rect 69305 2805 69339 2839
rect 69673 2805 69707 2839
rect 70869 2805 70903 2839
rect 72341 2805 72375 2839
rect 73353 2805 73387 2839
rect 75009 2805 75043 2839
rect 77769 2805 77803 2839
rect 80713 2805 80747 2839
rect 87613 2805 87647 2839
rect 89545 2805 89579 2839
rect 90741 2805 90775 2839
rect 91477 2805 91511 2839
rect 91845 2805 91879 2839
rect 92213 2805 92247 2839
rect 94973 2805 95007 2839
rect 97733 2805 97767 2839
rect 98469 2805 98503 2839
rect 100493 2805 100527 2839
rect 102977 2805 103011 2839
rect 104817 2805 104851 2839
rect 107669 2805 107703 2839
rect 112637 2805 112671 2839
rect 113557 2805 113591 2839
rect 117881 2805 117915 2839
rect 56149 2601 56183 2635
rect 56793 2601 56827 2635
rect 57161 2601 57195 2635
rect 58265 2601 58299 2635
rect 59645 2601 59679 2635
rect 64153 2601 64187 2635
rect 64705 2601 64739 2635
rect 65165 2601 65199 2635
rect 74641 2601 74675 2635
rect 75929 2601 75963 2635
rect 77217 2601 77251 2635
rect 78689 2601 78723 2635
rect 81081 2601 81115 2635
rect 82645 2601 82679 2635
rect 83657 2601 83691 2635
rect 84853 2601 84887 2635
rect 86233 2601 86267 2635
rect 87521 2601 87555 2635
rect 88809 2601 88843 2635
rect 90097 2601 90131 2635
rect 91569 2601 91603 2635
rect 93133 2601 93167 2635
rect 93961 2601 93995 2635
rect 95065 2601 95099 2635
rect 96537 2601 96571 2635
rect 100309 2601 100343 2635
rect 101689 2601 101723 2635
rect 102885 2601 102919 2635
rect 105093 2601 105127 2635
rect 107301 2601 107335 2635
rect 111073 2601 111107 2635
rect 111993 2601 112027 2635
rect 114937 2601 114971 2635
rect 17049 2533 17083 2567
rect 22569 2533 22603 2567
rect 97733 2533 97767 2567
rect 99113 2533 99147 2567
rect 109417 2533 109451 2567
rect 113281 2533 113315 2567
rect 75101 2465 75135 2499
rect 75285 2465 75319 2499
rect 76573 2465 76607 2499
rect 77861 2465 77895 2499
rect 79241 2465 79275 2499
rect 81541 2465 81575 2499
rect 81725 2465 81759 2499
rect 83197 2465 83231 2499
rect 84117 2465 84151 2499
rect 84209 2465 84243 2499
rect 85313 2465 85347 2499
rect 85497 2465 85531 2499
rect 86693 2465 86727 2499
rect 86785 2465 86819 2499
rect 87981 2465 88015 2499
rect 88165 2465 88199 2499
rect 89269 2465 89303 2499
rect 89361 2465 89395 2499
rect 90557 2465 90591 2499
rect 90741 2465 90775 2499
rect 92029 2465 92063 2499
rect 92213 2465 92247 2499
rect 95525 2465 95559 2499
rect 95709 2465 95743 2499
rect 96997 2465 97031 2499
rect 97181 2465 97215 2499
rect 98193 2465 98227 2499
rect 98377 2465 98411 2499
rect 99665 2465 99699 2499
rect 100769 2465 100803 2499
rect 100861 2465 100895 2499
rect 102333 2465 102367 2499
rect 103529 2465 103563 2499
rect 105553 2465 105587 2499
rect 105645 2465 105679 2499
rect 107761 2465 107795 2499
rect 107853 2465 107887 2499
rect 108865 2465 108899 2499
rect 109969 2465 110003 2499
rect 112453 2465 112487 2499
rect 112637 2465 112671 2499
rect 113741 2465 113775 2499
rect 113833 2465 113867 2499
rect 115397 2465 115431 2499
rect 115489 2465 115523 2499
rect 117329 2465 117363 2499
rect 1409 2397 1443 2431
rect 2145 2397 2179 2431
rect 3801 2397 3835 2431
rect 4997 2397 5031 2431
rect 6469 2397 6503 2431
rect 7573 2397 7607 2431
rect 7849 2397 7883 2431
rect 9321 2397 9355 2431
rect 10425 2397 10459 2431
rect 10701 2397 10735 2431
rect 12173 2397 12207 2431
rect 14105 2397 14139 2431
rect 22293 2397 22327 2431
rect 61393 2397 61427 2431
rect 62129 2397 62163 2431
rect 63509 2397 63543 2431
rect 64061 2397 64095 2431
rect 64889 2397 64923 2431
rect 65717 2397 65751 2431
rect 66729 2397 66763 2431
rect 68293 2397 68327 2431
rect 69581 2397 69615 2431
rect 72801 2397 72835 2431
rect 73537 2397 73571 2431
rect 80069 2397 80103 2431
rect 83013 2397 83047 2431
rect 85221 2397 85255 2431
rect 92949 2397 92983 2431
rect 94145 2397 94179 2431
rect 99573 2397 99607 2431
rect 102149 2397 102183 2431
rect 104449 2397 104483 2431
rect 105461 2397 105495 2431
rect 110797 2397 110831 2431
rect 111257 2397 111291 2431
rect 116501 2397 116535 2431
rect 117605 2397 117639 2431
rect 9965 2329 9999 2363
rect 15117 2329 15151 2363
rect 15485 2329 15519 2363
rect 16773 2329 16807 2363
rect 17969 2329 18003 2363
rect 18337 2329 18371 2363
rect 19349 2329 19383 2363
rect 20821 2329 20855 2363
rect 22109 2329 22143 2363
rect 24501 2329 24535 2363
rect 25421 2329 25455 2363
rect 27077 2329 27111 2363
rect 27997 2329 28031 2363
rect 29653 2329 29687 2363
rect 30021 2329 30055 2363
rect 30849 2329 30883 2363
rect 32229 2329 32263 2363
rect 32597 2329 32631 2363
rect 33701 2329 33735 2363
rect 35173 2329 35207 2363
rect 37381 2329 37415 2363
rect 38301 2329 38335 2363
rect 39957 2329 39991 2363
rect 40877 2329 40911 2363
rect 42533 2329 42567 2363
rect 43637 2329 43671 2363
rect 45109 2329 45143 2363
rect 46489 2329 46523 2363
rect 46857 2329 46891 2363
rect 47961 2329 47995 2363
rect 49249 2329 49283 2363
rect 50813 2329 50847 2363
rect 51181 2329 51215 2363
rect 52837 2329 52871 2363
rect 53757 2329 53791 2363
rect 54125 2329 54159 2363
rect 56517 2329 56551 2363
rect 57989 2329 58023 2363
rect 59553 2329 59587 2363
rect 61025 2329 61059 2363
rect 63141 2329 63175 2363
rect 71053 2329 71087 2363
rect 72433 2329 72467 2363
rect 76297 2329 76331 2363
rect 79149 2329 79183 2363
rect 99481 2329 99515 2363
rect 100125 2329 100159 2363
rect 108681 2329 108715 2363
rect 113649 2329 113683 2363
rect 115949 2329 115983 2363
rect 116777 2329 116811 2363
rect 1593 2261 1627 2295
rect 2329 2261 2363 2295
rect 3985 2261 4019 2295
rect 5181 2261 5215 2295
rect 6653 2261 6687 2295
rect 7113 2261 7147 2295
rect 8033 2261 8067 2295
rect 9505 2261 9539 2295
rect 10885 2261 10919 2295
rect 12357 2261 12391 2295
rect 14289 2261 14323 2295
rect 19625 2261 19659 2295
rect 20085 2261 20119 2295
rect 20453 2261 20487 2295
rect 21097 2261 21131 2295
rect 24777 2261 24811 2295
rect 25697 2261 25731 2295
rect 27353 2261 27387 2295
rect 28273 2261 28307 2295
rect 31125 2261 31159 2295
rect 32965 2261 32999 2295
rect 33333 2261 33367 2295
rect 33977 2261 34011 2295
rect 34989 2261 35023 2295
rect 35449 2261 35483 2295
rect 37657 2261 37691 2295
rect 38577 2261 38611 2295
rect 40233 2261 40267 2295
rect 41153 2261 41187 2295
rect 42809 2261 42843 2295
rect 43913 2261 43947 2295
rect 45201 2261 45235 2295
rect 48237 2261 48271 2295
rect 49525 2261 49559 2295
rect 53113 2261 53147 2295
rect 55781 2261 55815 2295
rect 62313 2261 62347 2295
rect 65809 2261 65843 2295
rect 66821 2261 66855 2295
rect 67373 2261 67407 2295
rect 68385 2261 68419 2295
rect 68937 2261 68971 2295
rect 69673 2261 69707 2295
rect 70225 2261 70259 2295
rect 71145 2261 71179 2295
rect 73721 2261 73755 2295
rect 75009 2261 75043 2295
rect 76389 2261 76423 2295
rect 77585 2261 77619 2295
rect 77677 2261 77711 2295
rect 79057 2261 79091 2295
rect 79701 2261 79735 2295
rect 79885 2261 79919 2295
rect 80621 2261 80655 2295
rect 81449 2261 81483 2295
rect 82093 2261 82127 2295
rect 82461 2261 82495 2295
rect 83105 2261 83139 2295
rect 84025 2261 84059 2295
rect 86601 2261 86635 2295
rect 87889 2261 87923 2295
rect 89177 2261 89211 2295
rect 90465 2261 90499 2295
rect 91937 2261 91971 2295
rect 95433 2261 95467 2295
rect 96905 2261 96939 2295
rect 98101 2261 98135 2295
rect 100677 2261 100711 2295
rect 102057 2261 102091 2295
rect 103253 2261 103287 2295
rect 103345 2261 103379 2295
rect 104265 2261 104299 2295
rect 107669 2261 107703 2295
rect 108313 2261 108347 2295
rect 109785 2261 109819 2295
rect 109877 2261 109911 2295
rect 110613 2261 110647 2295
rect 111533 2261 111567 2295
rect 112361 2261 112395 2295
rect 115305 2261 115339 2295
rect 116317 2261 116351 2295
<< metal1 >>
rect 1104 37562 118864 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 96374 37562
rect 96426 37510 96438 37562
rect 96490 37510 96502 37562
rect 96554 37510 96566 37562
rect 96618 37510 96630 37562
rect 96682 37510 118864 37562
rect 1104 37488 118864 37510
rect 117222 37408 117228 37460
rect 117280 37448 117286 37460
rect 117317 37451 117375 37457
rect 117317 37448 117329 37451
rect 117280 37420 117329 37448
rect 117280 37408 117286 37420
rect 117317 37417 117329 37420
rect 117363 37417 117375 37451
rect 118050 37448 118056 37460
rect 118011 37420 118056 37448
rect 117317 37411 117375 37417
rect 118050 37408 118056 37420
rect 118108 37408 118114 37460
rect 114922 37204 114928 37256
rect 114980 37244 114986 37256
rect 117133 37247 117191 37253
rect 117133 37244 117145 37247
rect 114980 37216 117145 37244
rect 114980 37204 114986 37216
rect 117133 37213 117145 37216
rect 117179 37213 117191 37247
rect 117133 37207 117191 37213
rect 117590 37204 117596 37256
rect 117648 37244 117654 37256
rect 117869 37247 117927 37253
rect 117869 37244 117881 37247
rect 117648 37216 117881 37244
rect 117648 37204 117654 37216
rect 117869 37213 117881 37216
rect 117915 37213 117927 37247
rect 117869 37207 117927 37213
rect 1104 37018 118864 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 81014 37018
rect 81066 36966 81078 37018
rect 81130 36966 81142 37018
rect 81194 36966 81206 37018
rect 81258 36966 81270 37018
rect 81322 36966 111734 37018
rect 111786 36966 111798 37018
rect 111850 36966 111862 37018
rect 111914 36966 111926 37018
rect 111978 36966 111990 37018
rect 112042 36966 118864 37018
rect 1104 36944 118864 36966
rect 117130 36864 117136 36916
rect 117188 36904 117194 36916
rect 117317 36907 117375 36913
rect 117317 36904 117329 36907
rect 117188 36876 117329 36904
rect 117188 36864 117194 36876
rect 117317 36873 117329 36876
rect 117363 36873 117375 36907
rect 117317 36867 117375 36873
rect 98914 36728 98920 36780
rect 98972 36768 98978 36780
rect 117133 36771 117191 36777
rect 117133 36768 117145 36771
rect 98972 36740 117145 36768
rect 98972 36728 98978 36740
rect 117133 36737 117145 36740
rect 117179 36737 117191 36771
rect 117133 36731 117191 36737
rect 117869 36771 117927 36777
rect 117869 36737 117881 36771
rect 117915 36768 117927 36771
rect 118418 36768 118424 36780
rect 117915 36740 118424 36768
rect 117915 36737 117927 36740
rect 117869 36731 117927 36737
rect 118418 36728 118424 36740
rect 118476 36728 118482 36780
rect 118050 36632 118056 36644
rect 118011 36604 118056 36632
rect 118050 36592 118056 36604
rect 118108 36592 118114 36644
rect 1104 36474 118864 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 96374 36474
rect 96426 36422 96438 36474
rect 96490 36422 96502 36474
rect 96554 36422 96566 36474
rect 96618 36422 96630 36474
rect 96682 36422 118864 36474
rect 1104 36400 118864 36422
rect 117869 36159 117927 36165
rect 117869 36125 117881 36159
rect 117915 36156 117927 36159
rect 118142 36156 118148 36168
rect 117915 36128 118148 36156
rect 117915 36125 117927 36128
rect 117869 36119 117927 36125
rect 118142 36116 118148 36128
rect 118200 36116 118206 36168
rect 118050 36020 118056 36032
rect 118011 35992 118056 36020
rect 118050 35980 118056 35992
rect 118108 35980 118114 36032
rect 1104 35930 118864 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 81014 35930
rect 81066 35878 81078 35930
rect 81130 35878 81142 35930
rect 81194 35878 81206 35930
rect 81258 35878 81270 35930
rect 81322 35878 111734 35930
rect 111786 35878 111798 35930
rect 111850 35878 111862 35930
rect 111914 35878 111926 35930
rect 111978 35878 111990 35930
rect 112042 35878 118864 35930
rect 1104 35856 118864 35878
rect 1104 35386 118864 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 96374 35386
rect 96426 35334 96438 35386
rect 96490 35334 96502 35386
rect 96554 35334 96566 35386
rect 96618 35334 96630 35386
rect 96682 35334 118864 35386
rect 1104 35312 118864 35334
rect 117682 35028 117688 35080
rect 117740 35068 117746 35080
rect 117869 35071 117927 35077
rect 117869 35068 117881 35071
rect 117740 35040 117881 35068
rect 117740 35028 117746 35040
rect 117869 35037 117881 35040
rect 117915 35037 117927 35071
rect 117869 35031 117927 35037
rect 118050 34932 118056 34944
rect 118011 34904 118056 34932
rect 118050 34892 118056 34904
rect 118108 34892 118114 34944
rect 1104 34842 118864 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 81014 34842
rect 81066 34790 81078 34842
rect 81130 34790 81142 34842
rect 81194 34790 81206 34842
rect 81258 34790 81270 34842
rect 81322 34790 111734 34842
rect 111786 34790 111798 34842
rect 111850 34790 111862 34842
rect 111914 34790 111926 34842
rect 111978 34790 111990 34842
rect 112042 34790 118864 34842
rect 1104 34768 118864 34790
rect 1104 34298 118864 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 96374 34298
rect 96426 34246 96438 34298
rect 96490 34246 96502 34298
rect 96554 34246 96566 34298
rect 96618 34246 96630 34298
rect 96682 34246 118864 34298
rect 1104 34224 118864 34246
rect 112162 33940 112168 33992
rect 112220 33980 112226 33992
rect 117869 33983 117927 33989
rect 117869 33980 117881 33983
rect 112220 33952 117881 33980
rect 112220 33940 112226 33952
rect 117869 33949 117881 33952
rect 117915 33949 117927 33983
rect 117869 33943 117927 33949
rect 118050 33844 118056 33856
rect 118011 33816 118056 33844
rect 118050 33804 118056 33816
rect 118108 33804 118114 33856
rect 1104 33754 118864 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 81014 33754
rect 81066 33702 81078 33754
rect 81130 33702 81142 33754
rect 81194 33702 81206 33754
rect 81258 33702 81270 33754
rect 81322 33702 111734 33754
rect 111786 33702 111798 33754
rect 111850 33702 111862 33754
rect 111914 33702 111926 33754
rect 111978 33702 111990 33754
rect 112042 33702 118864 33754
rect 1104 33680 118864 33702
rect 110782 33464 110788 33516
rect 110840 33504 110846 33516
rect 117869 33507 117927 33513
rect 117869 33504 117881 33507
rect 110840 33476 117881 33504
rect 110840 33464 110846 33476
rect 117869 33473 117881 33476
rect 117915 33473 117927 33507
rect 117869 33467 117927 33473
rect 118050 33300 118056 33312
rect 118011 33272 118056 33300
rect 118050 33260 118056 33272
rect 118108 33260 118114 33312
rect 1104 33210 118864 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 96374 33210
rect 96426 33158 96438 33210
rect 96490 33158 96502 33210
rect 96554 33158 96566 33210
rect 96618 33158 96630 33210
rect 96682 33158 118864 33210
rect 1104 33136 118864 33158
rect 1104 32666 118864 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 81014 32666
rect 81066 32614 81078 32666
rect 81130 32614 81142 32666
rect 81194 32614 81206 32666
rect 81258 32614 81270 32666
rect 81322 32614 111734 32666
rect 111786 32614 111798 32666
rect 111850 32614 111862 32666
rect 111914 32614 111926 32666
rect 111978 32614 111990 32666
rect 112042 32614 118864 32666
rect 1104 32592 118864 32614
rect 108482 32376 108488 32428
rect 108540 32416 108546 32428
rect 117869 32419 117927 32425
rect 117869 32416 117881 32419
rect 108540 32388 117881 32416
rect 108540 32376 108546 32388
rect 117869 32385 117881 32388
rect 117915 32385 117927 32419
rect 117869 32379 117927 32385
rect 118050 32212 118056 32224
rect 118011 32184 118056 32212
rect 118050 32172 118056 32184
rect 118108 32172 118114 32224
rect 1104 32122 118864 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 96374 32122
rect 96426 32070 96438 32122
rect 96490 32070 96502 32122
rect 96554 32070 96566 32122
rect 96618 32070 96630 32122
rect 96682 32070 118864 32122
rect 1104 32048 118864 32070
rect 1104 31578 118864 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 81014 31578
rect 81066 31526 81078 31578
rect 81130 31526 81142 31578
rect 81194 31526 81206 31578
rect 81258 31526 81270 31578
rect 81322 31526 111734 31578
rect 111786 31526 111798 31578
rect 111850 31526 111862 31578
rect 111914 31526 111926 31578
rect 111978 31526 111990 31578
rect 112042 31526 118864 31578
rect 1104 31504 118864 31526
rect 107102 31288 107108 31340
rect 107160 31328 107166 31340
rect 117869 31331 117927 31337
rect 117869 31328 117881 31331
rect 107160 31300 117881 31328
rect 107160 31288 107166 31300
rect 117869 31297 117881 31300
rect 117915 31297 117927 31331
rect 117869 31291 117927 31297
rect 118050 31124 118056 31136
rect 118011 31096 118056 31124
rect 118050 31084 118056 31096
rect 118108 31084 118114 31136
rect 1104 31034 118864 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 96374 31034
rect 96426 30982 96438 31034
rect 96490 30982 96502 31034
rect 96554 30982 96566 31034
rect 96618 30982 96630 31034
rect 96682 30982 118864 31034
rect 1104 30960 118864 30982
rect 1104 30490 118864 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 81014 30490
rect 81066 30438 81078 30490
rect 81130 30438 81142 30490
rect 81194 30438 81206 30490
rect 81258 30438 81270 30490
rect 81322 30438 111734 30490
rect 111786 30438 111798 30490
rect 111850 30438 111862 30490
rect 111914 30438 111926 30490
rect 111978 30438 111990 30490
rect 112042 30438 118864 30490
rect 1104 30416 118864 30438
rect 105998 30200 106004 30252
rect 106056 30240 106062 30252
rect 117869 30243 117927 30249
rect 117869 30240 117881 30243
rect 106056 30212 117881 30240
rect 106056 30200 106062 30212
rect 117869 30209 117881 30212
rect 117915 30209 117927 30243
rect 117869 30203 117927 30209
rect 118050 30104 118056 30116
rect 118011 30076 118056 30104
rect 118050 30064 118056 30076
rect 118108 30064 118114 30116
rect 1104 29946 118864 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 96374 29946
rect 96426 29894 96438 29946
rect 96490 29894 96502 29946
rect 96554 29894 96566 29946
rect 96618 29894 96630 29946
rect 96682 29894 118864 29946
rect 1104 29872 118864 29894
rect 104434 29588 104440 29640
rect 104492 29628 104498 29640
rect 117869 29631 117927 29637
rect 117869 29628 117881 29631
rect 104492 29600 117881 29628
rect 104492 29588 104498 29600
rect 117869 29597 117881 29600
rect 117915 29597 117927 29631
rect 117869 29591 117927 29597
rect 118050 29492 118056 29504
rect 118011 29464 118056 29492
rect 118050 29452 118056 29464
rect 118108 29452 118114 29504
rect 1104 29402 118864 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 81014 29402
rect 81066 29350 81078 29402
rect 81130 29350 81142 29402
rect 81194 29350 81206 29402
rect 81258 29350 81270 29402
rect 81322 29350 111734 29402
rect 111786 29350 111798 29402
rect 111850 29350 111862 29402
rect 111914 29350 111926 29402
rect 111978 29350 111990 29402
rect 112042 29350 118864 29402
rect 1104 29328 118864 29350
rect 1104 28858 118864 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 96374 28858
rect 96426 28806 96438 28858
rect 96490 28806 96502 28858
rect 96554 28806 96566 28858
rect 96618 28806 96630 28858
rect 96682 28806 118864 28858
rect 1104 28784 118864 28806
rect 102410 28500 102416 28552
rect 102468 28540 102474 28552
rect 117869 28543 117927 28549
rect 117869 28540 117881 28543
rect 102468 28512 117881 28540
rect 102468 28500 102474 28512
rect 117869 28509 117881 28512
rect 117915 28509 117927 28543
rect 117869 28503 117927 28509
rect 118050 28404 118056 28416
rect 118011 28376 118056 28404
rect 118050 28364 118056 28376
rect 118108 28364 118114 28416
rect 1104 28314 118864 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 81014 28314
rect 81066 28262 81078 28314
rect 81130 28262 81142 28314
rect 81194 28262 81206 28314
rect 81258 28262 81270 28314
rect 81322 28262 111734 28314
rect 111786 28262 111798 28314
rect 111850 28262 111862 28314
rect 111914 28262 111926 28314
rect 111978 28262 111990 28314
rect 112042 28262 118864 28314
rect 1104 28240 118864 28262
rect 1104 27770 118864 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 96374 27770
rect 96426 27718 96438 27770
rect 96490 27718 96502 27770
rect 96554 27718 96566 27770
rect 96618 27718 96630 27770
rect 96682 27718 118864 27770
rect 1104 27696 118864 27718
rect 100570 27412 100576 27464
rect 100628 27452 100634 27464
rect 117869 27455 117927 27461
rect 117869 27452 117881 27455
rect 100628 27424 117881 27452
rect 100628 27412 100634 27424
rect 117869 27421 117881 27424
rect 117915 27421 117927 27455
rect 117869 27415 117927 27421
rect 118050 27316 118056 27328
rect 118011 27288 118056 27316
rect 118050 27276 118056 27288
rect 118108 27276 118114 27328
rect 1104 27226 118864 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 81014 27226
rect 81066 27174 81078 27226
rect 81130 27174 81142 27226
rect 81194 27174 81206 27226
rect 81258 27174 81270 27226
rect 81322 27174 111734 27226
rect 111786 27174 111798 27226
rect 111850 27174 111862 27226
rect 111914 27174 111926 27226
rect 111978 27174 111990 27226
rect 112042 27174 118864 27226
rect 1104 27152 118864 27174
rect 99834 26936 99840 26988
rect 99892 26976 99898 26988
rect 117869 26979 117927 26985
rect 117869 26976 117881 26979
rect 99892 26948 117881 26976
rect 99892 26936 99898 26948
rect 117869 26945 117881 26948
rect 117915 26945 117927 26979
rect 117869 26939 117927 26945
rect 118050 26772 118056 26784
rect 118011 26744 118056 26772
rect 118050 26732 118056 26744
rect 118108 26732 118114 26784
rect 1104 26682 118864 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 96374 26682
rect 96426 26630 96438 26682
rect 96490 26630 96502 26682
rect 96554 26630 96566 26682
rect 96618 26630 96630 26682
rect 96682 26630 118864 26682
rect 1104 26608 118864 26630
rect 1104 26138 118864 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 81014 26138
rect 81066 26086 81078 26138
rect 81130 26086 81142 26138
rect 81194 26086 81206 26138
rect 81258 26086 81270 26138
rect 81322 26086 111734 26138
rect 111786 26086 111798 26138
rect 111850 26086 111862 26138
rect 111914 26086 111926 26138
rect 111978 26086 111990 26138
rect 112042 26086 118864 26138
rect 1104 26064 118864 26086
rect 98086 25848 98092 25900
rect 98144 25888 98150 25900
rect 117501 25891 117559 25897
rect 117501 25888 117513 25891
rect 98144 25860 117513 25888
rect 98144 25848 98150 25860
rect 117501 25857 117513 25860
rect 117547 25888 117559 25891
rect 117869 25891 117927 25897
rect 117869 25888 117881 25891
rect 117547 25860 117881 25888
rect 117547 25857 117559 25860
rect 117501 25851 117559 25857
rect 117869 25857 117881 25860
rect 117915 25857 117927 25891
rect 117869 25851 117927 25857
rect 118050 25684 118056 25696
rect 118011 25656 118056 25684
rect 118050 25644 118056 25656
rect 118108 25644 118114 25696
rect 1104 25594 118864 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 96374 25594
rect 96426 25542 96438 25594
rect 96490 25542 96502 25594
rect 96554 25542 96566 25594
rect 96618 25542 96630 25594
rect 96682 25542 118864 25594
rect 1104 25520 118864 25542
rect 1104 25050 118864 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 81014 25050
rect 81066 24998 81078 25050
rect 81130 24998 81142 25050
rect 81194 24998 81206 25050
rect 81258 24998 81270 25050
rect 81322 24998 111734 25050
rect 111786 24998 111798 25050
rect 111850 24998 111862 25050
rect 111914 24998 111926 25050
rect 111978 24998 111990 25050
rect 112042 24998 118864 25050
rect 1104 24976 118864 24998
rect 96890 24760 96896 24812
rect 96948 24800 96954 24812
rect 117501 24803 117559 24809
rect 117501 24800 117513 24803
rect 96948 24772 117513 24800
rect 96948 24760 96954 24772
rect 117501 24769 117513 24772
rect 117547 24800 117559 24803
rect 117869 24803 117927 24809
rect 117869 24800 117881 24803
rect 117547 24772 117881 24800
rect 117547 24769 117559 24772
rect 117501 24763 117559 24769
rect 117869 24769 117881 24772
rect 117915 24769 117927 24803
rect 117869 24763 117927 24769
rect 118050 24596 118056 24608
rect 118011 24568 118056 24596
rect 118050 24556 118056 24568
rect 118108 24556 118114 24608
rect 1104 24506 118864 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 96374 24506
rect 96426 24454 96438 24506
rect 96490 24454 96502 24506
rect 96554 24454 96566 24506
rect 96618 24454 96630 24506
rect 96682 24454 118864 24506
rect 1104 24432 118864 24454
rect 1104 23962 118864 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 81014 23962
rect 81066 23910 81078 23962
rect 81130 23910 81142 23962
rect 81194 23910 81206 23962
rect 81258 23910 81270 23962
rect 81322 23910 111734 23962
rect 111786 23910 111798 23962
rect 111850 23910 111862 23962
rect 111914 23910 111926 23962
rect 111978 23910 111990 23962
rect 112042 23910 118864 23962
rect 1104 23888 118864 23910
rect 95970 23672 95976 23724
rect 96028 23712 96034 23724
rect 117501 23715 117559 23721
rect 117501 23712 117513 23715
rect 96028 23684 117513 23712
rect 96028 23672 96034 23684
rect 117501 23681 117513 23684
rect 117547 23712 117559 23715
rect 117869 23715 117927 23721
rect 117869 23712 117881 23715
rect 117547 23684 117881 23712
rect 117547 23681 117559 23684
rect 117501 23675 117559 23681
rect 117869 23681 117881 23684
rect 117915 23681 117927 23715
rect 117869 23675 117927 23681
rect 118050 23576 118056 23588
rect 118011 23548 118056 23576
rect 118050 23536 118056 23548
rect 118108 23536 118114 23588
rect 1104 23418 118864 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 96374 23418
rect 96426 23366 96438 23418
rect 96490 23366 96502 23418
rect 96554 23366 96566 23418
rect 96618 23366 96630 23418
rect 96682 23366 118864 23418
rect 1104 23344 118864 23366
rect 93118 23060 93124 23112
rect 93176 23100 93182 23112
rect 117501 23103 117559 23109
rect 117501 23100 117513 23103
rect 93176 23072 117513 23100
rect 93176 23060 93182 23072
rect 117501 23069 117513 23072
rect 117547 23100 117559 23103
rect 117869 23103 117927 23109
rect 117869 23100 117881 23103
rect 117547 23072 117881 23100
rect 117547 23069 117559 23072
rect 117501 23063 117559 23069
rect 117869 23069 117881 23072
rect 117915 23069 117927 23103
rect 117869 23063 117927 23069
rect 118050 22964 118056 22976
rect 118011 22936 118056 22964
rect 118050 22924 118056 22936
rect 118108 22924 118114 22976
rect 1104 22874 118864 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 81014 22874
rect 81066 22822 81078 22874
rect 81130 22822 81142 22874
rect 81194 22822 81206 22874
rect 81258 22822 81270 22874
rect 81322 22822 111734 22874
rect 111786 22822 111798 22874
rect 111850 22822 111862 22874
rect 111914 22822 111926 22874
rect 111978 22822 111990 22874
rect 112042 22822 118864 22874
rect 1104 22800 118864 22822
rect 1104 22330 118864 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 96374 22330
rect 96426 22278 96438 22330
rect 96490 22278 96502 22330
rect 96554 22278 96566 22330
rect 96618 22278 96630 22330
rect 96682 22278 118864 22330
rect 1104 22256 118864 22278
rect 117869 22015 117927 22021
rect 117869 22012 117881 22015
rect 117516 21984 117881 22012
rect 92382 21836 92388 21888
rect 92440 21876 92446 21888
rect 117516 21885 117544 21984
rect 117869 21981 117881 21984
rect 117915 21981 117927 22015
rect 117869 21975 117927 21981
rect 117501 21879 117559 21885
rect 117501 21876 117513 21879
rect 92440 21848 117513 21876
rect 92440 21836 92446 21848
rect 117501 21845 117513 21848
rect 117547 21845 117559 21879
rect 118050 21876 118056 21888
rect 118011 21848 118056 21876
rect 117501 21839 117559 21845
rect 118050 21836 118056 21848
rect 118108 21836 118114 21888
rect 1104 21786 118864 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 81014 21786
rect 81066 21734 81078 21786
rect 81130 21734 81142 21786
rect 81194 21734 81206 21786
rect 81258 21734 81270 21786
rect 81322 21734 111734 21786
rect 111786 21734 111798 21786
rect 111850 21734 111862 21786
rect 111914 21734 111926 21786
rect 111978 21734 111990 21786
rect 112042 21734 118864 21786
rect 1104 21712 118864 21734
rect 1104 21242 118864 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 96374 21242
rect 96426 21190 96438 21242
rect 96490 21190 96502 21242
rect 96554 21190 96566 21242
rect 96618 21190 96630 21242
rect 96682 21190 118864 21242
rect 1104 21168 118864 21190
rect 91002 20884 91008 20936
rect 91060 20924 91066 20936
rect 117501 20927 117559 20933
rect 117501 20924 117513 20927
rect 91060 20896 117513 20924
rect 91060 20884 91066 20896
rect 117501 20893 117513 20896
rect 117547 20924 117559 20927
rect 117869 20927 117927 20933
rect 117869 20924 117881 20927
rect 117547 20896 117881 20924
rect 117547 20893 117559 20896
rect 117501 20887 117559 20893
rect 117869 20893 117881 20896
rect 117915 20893 117927 20927
rect 117869 20887 117927 20893
rect 118050 20788 118056 20800
rect 118011 20760 118056 20788
rect 118050 20748 118056 20760
rect 118108 20748 118114 20800
rect 1104 20698 118864 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 81014 20698
rect 81066 20646 81078 20698
rect 81130 20646 81142 20698
rect 81194 20646 81206 20698
rect 81258 20646 81270 20698
rect 81322 20646 111734 20698
rect 111786 20646 111798 20698
rect 111850 20646 111862 20698
rect 111914 20646 111926 20698
rect 111978 20646 111990 20698
rect 112042 20646 118864 20698
rect 1104 20624 118864 20646
rect 89438 20408 89444 20460
rect 89496 20448 89502 20460
rect 117501 20451 117559 20457
rect 117501 20448 117513 20451
rect 89496 20420 117513 20448
rect 89496 20408 89502 20420
rect 117501 20417 117513 20420
rect 117547 20448 117559 20451
rect 117869 20451 117927 20457
rect 117869 20448 117881 20451
rect 117547 20420 117881 20448
rect 117547 20417 117559 20420
rect 117501 20411 117559 20417
rect 117869 20417 117881 20420
rect 117915 20417 117927 20451
rect 117869 20411 117927 20417
rect 118050 20244 118056 20256
rect 118011 20216 118056 20244
rect 118050 20204 118056 20216
rect 118108 20204 118114 20256
rect 1104 20154 118864 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 96374 20154
rect 96426 20102 96438 20154
rect 96490 20102 96502 20154
rect 96554 20102 96566 20154
rect 96618 20102 96630 20154
rect 96682 20102 118864 20154
rect 1104 20080 118864 20102
rect 1104 19610 118864 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 81014 19610
rect 81066 19558 81078 19610
rect 81130 19558 81142 19610
rect 81194 19558 81206 19610
rect 81258 19558 81270 19610
rect 81322 19558 111734 19610
rect 111786 19558 111798 19610
rect 111850 19558 111862 19610
rect 111914 19558 111926 19610
rect 111978 19558 111990 19610
rect 112042 19558 118864 19610
rect 1104 19536 118864 19558
rect 117869 19363 117927 19369
rect 117869 19360 117881 19363
rect 117516 19332 117881 19360
rect 117406 19116 117412 19168
rect 117464 19156 117470 19168
rect 117516 19165 117544 19332
rect 117869 19329 117881 19332
rect 117915 19329 117927 19363
rect 117869 19323 117927 19329
rect 117501 19159 117559 19165
rect 117501 19156 117513 19159
rect 117464 19128 117513 19156
rect 117464 19116 117470 19128
rect 117501 19125 117513 19128
rect 117547 19125 117559 19159
rect 118050 19156 118056 19168
rect 118011 19128 118056 19156
rect 117501 19119 117559 19125
rect 118050 19116 118056 19128
rect 118108 19116 118114 19168
rect 1104 19066 118864 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 96374 19066
rect 96426 19014 96438 19066
rect 96490 19014 96502 19066
rect 96554 19014 96566 19066
rect 96618 19014 96630 19066
rect 96682 19014 118864 19066
rect 1104 18992 118864 19014
rect 1104 18522 118864 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 81014 18522
rect 81066 18470 81078 18522
rect 81130 18470 81142 18522
rect 81194 18470 81206 18522
rect 81258 18470 81270 18522
rect 81322 18470 111734 18522
rect 111786 18470 111798 18522
rect 111850 18470 111862 18522
rect 111914 18470 111926 18522
rect 111978 18470 111990 18522
rect 112042 18470 118864 18522
rect 1104 18448 118864 18470
rect 117869 18275 117927 18281
rect 117869 18272 117881 18275
rect 117516 18244 117881 18272
rect 86678 18028 86684 18080
rect 86736 18068 86742 18080
rect 117516 18077 117544 18244
rect 117869 18241 117881 18244
rect 117915 18241 117927 18275
rect 117869 18235 117927 18241
rect 117501 18071 117559 18077
rect 117501 18068 117513 18071
rect 86736 18040 117513 18068
rect 86736 18028 86742 18040
rect 117501 18037 117513 18040
rect 117547 18037 117559 18071
rect 118050 18068 118056 18080
rect 118011 18040 118056 18068
rect 117501 18031 117559 18037
rect 118050 18028 118056 18040
rect 118108 18028 118114 18080
rect 1104 17978 118864 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 96374 17978
rect 96426 17926 96438 17978
rect 96490 17926 96502 17978
rect 96554 17926 96566 17978
rect 96618 17926 96630 17978
rect 96682 17926 118864 17978
rect 1104 17904 118864 17926
rect 85206 17620 85212 17672
rect 85264 17660 85270 17672
rect 117501 17663 117559 17669
rect 117501 17660 117513 17663
rect 85264 17632 117513 17660
rect 85264 17620 85270 17632
rect 117501 17629 117513 17632
rect 117547 17660 117559 17663
rect 117869 17663 117927 17669
rect 117869 17660 117881 17663
rect 117547 17632 117881 17660
rect 117547 17629 117559 17632
rect 117501 17623 117559 17629
rect 117869 17629 117881 17632
rect 117915 17629 117927 17663
rect 117869 17623 117927 17629
rect 118050 17524 118056 17536
rect 118011 17496 118056 17524
rect 118050 17484 118056 17496
rect 118108 17484 118114 17536
rect 1104 17434 118864 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 81014 17434
rect 81066 17382 81078 17434
rect 81130 17382 81142 17434
rect 81194 17382 81206 17434
rect 81258 17382 81270 17434
rect 81322 17382 111734 17434
rect 111786 17382 111798 17434
rect 111850 17382 111862 17434
rect 111914 17382 111926 17434
rect 111978 17382 111990 17434
rect 112042 17382 118864 17434
rect 1104 17360 118864 17382
rect 1104 16890 118864 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 96374 16890
rect 96426 16838 96438 16890
rect 96490 16838 96502 16890
rect 96554 16838 96566 16890
rect 96618 16838 96630 16890
rect 96682 16838 118864 16890
rect 1104 16816 118864 16838
rect 117869 16575 117927 16581
rect 117869 16572 117881 16575
rect 117516 16544 117881 16572
rect 117516 16448 117544 16544
rect 117869 16541 117881 16544
rect 117915 16541 117927 16575
rect 117869 16535 117927 16541
rect 117498 16436 117504 16448
rect 117459 16408 117504 16436
rect 117498 16396 117504 16408
rect 117556 16396 117562 16448
rect 118050 16436 118056 16448
rect 118011 16408 118056 16436
rect 118050 16396 118056 16408
rect 118108 16396 118114 16448
rect 1104 16346 118864 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 81014 16346
rect 81066 16294 81078 16346
rect 81130 16294 81142 16346
rect 81194 16294 81206 16346
rect 81258 16294 81270 16346
rect 81322 16294 111734 16346
rect 111786 16294 111798 16346
rect 111850 16294 111862 16346
rect 111914 16294 111926 16346
rect 111978 16294 111990 16346
rect 112042 16294 118864 16346
rect 1104 16272 118864 16294
rect 1104 15802 118864 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 96374 15802
rect 96426 15750 96438 15802
rect 96490 15750 96502 15802
rect 96554 15750 96566 15802
rect 96618 15750 96630 15802
rect 96682 15750 118864 15802
rect 1104 15728 118864 15750
rect 82814 15444 82820 15496
rect 82872 15484 82878 15496
rect 117501 15487 117559 15493
rect 117501 15484 117513 15487
rect 82872 15456 117513 15484
rect 82872 15444 82878 15456
rect 117501 15453 117513 15456
rect 117547 15484 117559 15487
rect 117869 15487 117927 15493
rect 117869 15484 117881 15487
rect 117547 15456 117881 15484
rect 117547 15453 117559 15456
rect 117501 15447 117559 15453
rect 117869 15453 117881 15456
rect 117915 15453 117927 15487
rect 117869 15447 117927 15453
rect 118050 15348 118056 15360
rect 118011 15320 118056 15348
rect 118050 15308 118056 15320
rect 118108 15308 118114 15360
rect 1104 15258 118864 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 81014 15258
rect 81066 15206 81078 15258
rect 81130 15206 81142 15258
rect 81194 15206 81206 15258
rect 81258 15206 81270 15258
rect 81322 15206 111734 15258
rect 111786 15206 111798 15258
rect 111850 15206 111862 15258
rect 111914 15206 111926 15258
rect 111978 15206 111990 15258
rect 112042 15206 118864 15258
rect 1104 15184 118864 15206
rect 1104 14714 118864 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 96374 14714
rect 96426 14662 96438 14714
rect 96490 14662 96502 14714
rect 96554 14662 96566 14714
rect 96618 14662 96630 14714
rect 96682 14662 118864 14714
rect 1104 14640 118864 14662
rect 81710 14356 81716 14408
rect 81768 14396 81774 14408
rect 117501 14399 117559 14405
rect 117501 14396 117513 14399
rect 81768 14368 117513 14396
rect 81768 14356 81774 14368
rect 117501 14365 117513 14368
rect 117547 14396 117559 14399
rect 117869 14399 117927 14405
rect 117869 14396 117881 14399
rect 117547 14368 117881 14396
rect 117547 14365 117559 14368
rect 117501 14359 117559 14365
rect 117869 14365 117881 14368
rect 117915 14365 117927 14399
rect 117869 14359 117927 14365
rect 118050 14260 118056 14272
rect 118011 14232 118056 14260
rect 118050 14220 118056 14232
rect 118108 14220 118114 14272
rect 1104 14170 118864 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 81014 14170
rect 81066 14118 81078 14170
rect 81130 14118 81142 14170
rect 81194 14118 81206 14170
rect 81258 14118 81270 14170
rect 81322 14118 111734 14170
rect 111786 14118 111798 14170
rect 111850 14118 111862 14170
rect 111914 14118 111926 14170
rect 111978 14118 111990 14170
rect 112042 14118 118864 14170
rect 1104 14096 118864 14118
rect 79594 13880 79600 13932
rect 79652 13920 79658 13932
rect 117501 13923 117559 13929
rect 117501 13920 117513 13923
rect 79652 13892 117513 13920
rect 79652 13880 79658 13892
rect 117501 13889 117513 13892
rect 117547 13920 117559 13923
rect 117869 13923 117927 13929
rect 117869 13920 117881 13923
rect 117547 13892 117881 13920
rect 117547 13889 117559 13892
rect 117501 13883 117559 13889
rect 117869 13889 117881 13892
rect 117915 13889 117927 13923
rect 117869 13883 117927 13889
rect 118050 13716 118056 13728
rect 118011 13688 118056 13716
rect 118050 13676 118056 13688
rect 118108 13676 118114 13728
rect 1104 13626 118864 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 96374 13626
rect 96426 13574 96438 13626
rect 96490 13574 96502 13626
rect 96554 13574 96566 13626
rect 96618 13574 96630 13626
rect 96682 13574 118864 13626
rect 1104 13552 118864 13574
rect 1104 13082 118864 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 81014 13082
rect 81066 13030 81078 13082
rect 81130 13030 81142 13082
rect 81194 13030 81206 13082
rect 81258 13030 81270 13082
rect 81322 13030 111734 13082
rect 111786 13030 111798 13082
rect 111850 13030 111862 13082
rect 111914 13030 111926 13082
rect 111978 13030 111990 13082
rect 112042 13030 118864 13082
rect 1104 13008 118864 13030
rect 89438 12968 89444 12980
rect 89399 12940 89444 12968
rect 89438 12928 89444 12940
rect 89496 12928 89502 12980
rect 78674 12792 78680 12844
rect 78732 12832 78738 12844
rect 78732 12804 84194 12832
rect 78732 12792 78738 12804
rect 84166 12764 84194 12804
rect 88794 12792 88800 12844
rect 88852 12832 88858 12844
rect 89257 12835 89315 12841
rect 89257 12832 89269 12835
rect 88852 12804 89269 12832
rect 88852 12792 88858 12804
rect 89257 12801 89269 12804
rect 89303 12801 89315 12835
rect 117501 12835 117559 12841
rect 117501 12832 117513 12835
rect 89257 12795 89315 12801
rect 93826 12804 117513 12832
rect 93826 12764 93854 12804
rect 117501 12801 117513 12804
rect 117547 12832 117559 12835
rect 117869 12835 117927 12841
rect 117869 12832 117881 12835
rect 117547 12804 117881 12832
rect 117547 12801 117559 12804
rect 117501 12795 117559 12801
rect 117869 12801 117881 12804
rect 117915 12801 117927 12835
rect 117869 12795 117927 12801
rect 84166 12736 93854 12764
rect 118050 12628 118056 12640
rect 118011 12600 118056 12628
rect 118050 12588 118056 12600
rect 118108 12588 118114 12640
rect 1104 12538 118864 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 96374 12538
rect 96426 12486 96438 12538
rect 96490 12486 96502 12538
rect 96554 12486 96566 12538
rect 96618 12486 96630 12538
rect 96682 12486 118864 12538
rect 1104 12464 118864 12486
rect 1104 11994 118864 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 81014 11994
rect 81066 11942 81078 11994
rect 81130 11942 81142 11994
rect 81194 11942 81206 11994
rect 81258 11942 81270 11994
rect 81322 11942 111734 11994
rect 111786 11942 111798 11994
rect 111850 11942 111862 11994
rect 111914 11942 111926 11994
rect 111978 11942 111990 11994
rect 112042 11942 118864 11994
rect 1104 11920 118864 11942
rect 117869 11747 117927 11753
rect 117869 11744 117881 11747
rect 117516 11716 117881 11744
rect 76650 11500 76656 11552
rect 76708 11540 76714 11552
rect 117516 11549 117544 11716
rect 117869 11713 117881 11716
rect 117915 11713 117927 11747
rect 117869 11707 117927 11713
rect 118050 11608 118056 11620
rect 118011 11580 118056 11608
rect 118050 11568 118056 11580
rect 118108 11568 118114 11620
rect 117501 11543 117559 11549
rect 117501 11540 117513 11543
rect 76708 11512 117513 11540
rect 76708 11500 76714 11512
rect 117501 11509 117513 11512
rect 117547 11509 117559 11543
rect 117501 11503 117559 11509
rect 1104 11450 118864 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 96374 11450
rect 96426 11398 96438 11450
rect 96490 11398 96502 11450
rect 96554 11398 96566 11450
rect 96618 11398 96630 11450
rect 96682 11398 118864 11450
rect 1104 11376 118864 11398
rect 118050 11268 118056 11280
rect 118011 11240 118056 11268
rect 118050 11228 118056 11240
rect 118108 11228 118114 11280
rect 76098 11092 76104 11144
rect 76156 11132 76162 11144
rect 117501 11135 117559 11141
rect 117501 11132 117513 11135
rect 76156 11104 117513 11132
rect 76156 11092 76162 11104
rect 117501 11101 117513 11104
rect 117547 11132 117559 11135
rect 117869 11135 117927 11141
rect 117869 11132 117881 11135
rect 117547 11104 117881 11132
rect 117547 11101 117559 11104
rect 117501 11095 117559 11101
rect 117869 11101 117881 11104
rect 117915 11101 117927 11135
rect 117869 11095 117927 11101
rect 1104 10906 118864 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 81014 10906
rect 81066 10854 81078 10906
rect 81130 10854 81142 10906
rect 81194 10854 81206 10906
rect 81258 10854 81270 10906
rect 81322 10854 111734 10906
rect 111786 10854 111798 10906
rect 111850 10854 111862 10906
rect 111914 10854 111926 10906
rect 111978 10854 111990 10906
rect 112042 10854 118864 10906
rect 1104 10832 118864 10854
rect 1104 10362 118864 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 96374 10362
rect 96426 10310 96438 10362
rect 96490 10310 96502 10362
rect 96554 10310 96566 10362
rect 96618 10310 96630 10362
rect 96682 10310 118864 10362
rect 1104 10288 118864 10310
rect 76098 10248 76104 10260
rect 76059 10220 76104 10248
rect 76098 10208 76104 10220
rect 76156 10208 76162 10260
rect 74626 10004 74632 10056
rect 74684 10044 74690 10056
rect 75917 10047 75975 10053
rect 75917 10044 75929 10047
rect 74684 10016 75929 10044
rect 74684 10004 74690 10016
rect 75917 10013 75929 10016
rect 75963 10013 75975 10047
rect 75917 10007 75975 10013
rect 117774 9976 117780 9988
rect 117735 9948 117780 9976
rect 117774 9936 117780 9948
rect 117832 9936 117838 9988
rect 107654 9868 107660 9920
rect 107712 9908 107718 9920
rect 117869 9911 117927 9917
rect 117869 9908 117881 9911
rect 107712 9880 117881 9908
rect 107712 9868 107718 9880
rect 117869 9877 117881 9880
rect 117915 9877 117927 9911
rect 117869 9871 117927 9877
rect 1104 9818 118864 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 81014 9818
rect 81066 9766 81078 9818
rect 81130 9766 81142 9818
rect 81194 9766 81206 9818
rect 81258 9766 81270 9818
rect 81322 9766 111734 9818
rect 111786 9766 111798 9818
rect 111850 9766 111862 9818
rect 111914 9766 111926 9818
rect 111978 9766 111990 9818
rect 112042 9766 118864 9818
rect 1104 9744 118864 9766
rect 1104 9274 118864 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 96374 9274
rect 96426 9222 96438 9274
rect 96490 9222 96502 9274
rect 96554 9222 96566 9274
rect 96618 9222 96630 9274
rect 96682 9222 118864 9274
rect 1104 9200 118864 9222
rect 117774 8888 117780 8900
rect 117735 8860 117780 8888
rect 117774 8848 117780 8860
rect 117832 8848 117838 8900
rect 73522 8780 73528 8832
rect 73580 8820 73586 8832
rect 117869 8823 117927 8829
rect 117869 8820 117881 8823
rect 73580 8792 117881 8820
rect 73580 8780 73586 8792
rect 117869 8789 117881 8792
rect 117915 8789 117927 8823
rect 117869 8783 117927 8789
rect 1104 8730 118864 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 81014 8730
rect 81066 8678 81078 8730
rect 81130 8678 81142 8730
rect 81194 8678 81206 8730
rect 81258 8678 81270 8730
rect 81322 8678 111734 8730
rect 111786 8678 111798 8730
rect 111850 8678 111862 8730
rect 111914 8678 111926 8730
rect 111978 8678 111990 8730
rect 112042 8678 118864 8730
rect 1104 8656 118864 8678
rect 1104 8186 118864 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 96374 8186
rect 96426 8134 96438 8186
rect 96490 8134 96502 8186
rect 96554 8134 96566 8186
rect 96618 8134 96630 8186
rect 96682 8134 118864 8186
rect 1104 8112 118864 8134
rect 117774 7800 117780 7812
rect 117735 7772 117780 7800
rect 117774 7760 117780 7772
rect 117832 7760 117838 7812
rect 71682 7692 71688 7744
rect 71740 7732 71746 7744
rect 117869 7735 117927 7741
rect 117869 7732 117881 7735
rect 71740 7704 117881 7732
rect 71740 7692 71746 7704
rect 117869 7701 117881 7704
rect 117915 7701 117927 7735
rect 117869 7695 117927 7701
rect 1104 7642 118864 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 81014 7642
rect 81066 7590 81078 7642
rect 81130 7590 81142 7642
rect 81194 7590 81206 7642
rect 81258 7590 81270 7642
rect 81322 7590 111734 7642
rect 111786 7590 111798 7642
rect 111850 7590 111862 7642
rect 111914 7590 111926 7642
rect 111978 7590 111990 7642
rect 112042 7590 118864 7642
rect 1104 7568 118864 7590
rect 117774 7392 117780 7404
rect 117735 7364 117780 7392
rect 117774 7352 117780 7364
rect 117832 7352 117838 7404
rect 116854 7148 116860 7200
rect 116912 7188 116918 7200
rect 117869 7191 117927 7197
rect 117869 7188 117881 7191
rect 116912 7160 117881 7188
rect 116912 7148 116918 7160
rect 117869 7157 117881 7160
rect 117915 7157 117927 7191
rect 117869 7151 117927 7157
rect 1104 7098 118864 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 96374 7098
rect 96426 7046 96438 7098
rect 96490 7046 96502 7098
rect 96554 7046 96566 7098
rect 96618 7046 96630 7098
rect 96682 7046 118864 7098
rect 1104 7024 118864 7046
rect 1104 6554 118864 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 81014 6554
rect 81066 6502 81078 6554
rect 81130 6502 81142 6554
rect 81194 6502 81206 6554
rect 81258 6502 81270 6554
rect 81322 6502 111734 6554
rect 111786 6502 111798 6554
rect 111850 6502 111862 6554
rect 111914 6502 111926 6554
rect 111978 6502 111990 6554
rect 112042 6502 118864 6554
rect 1104 6480 118864 6502
rect 91002 6440 91008 6452
rect 90963 6412 91008 6440
rect 91002 6400 91008 6412
rect 91060 6400 91066 6452
rect 88334 6264 88340 6316
rect 88392 6304 88398 6316
rect 88797 6307 88855 6313
rect 88797 6304 88809 6307
rect 88392 6276 88809 6304
rect 88392 6264 88398 6276
rect 88797 6273 88809 6276
rect 88843 6273 88855 6307
rect 90818 6304 90824 6316
rect 90779 6276 90824 6304
rect 88797 6267 88855 6273
rect 90818 6264 90824 6276
rect 90876 6264 90882 6316
rect 117406 6304 117412 6316
rect 99346 6276 117412 6304
rect 88981 6103 89039 6109
rect 88981 6069 88993 6103
rect 89027 6100 89039 6103
rect 99346 6100 99374 6276
rect 117406 6264 117412 6276
rect 117464 6264 117470 6316
rect 117774 6304 117780 6316
rect 117735 6276 117780 6304
rect 117774 6264 117780 6276
rect 117832 6264 117838 6316
rect 89027 6072 99374 6100
rect 89027 6069 89039 6072
rect 88981 6063 89039 6069
rect 117498 6060 117504 6112
rect 117556 6100 117562 6112
rect 117869 6103 117927 6109
rect 117869 6100 117881 6103
rect 117556 6072 117881 6100
rect 117556 6060 117562 6072
rect 117869 6069 117881 6072
rect 117915 6069 117927 6103
rect 117869 6063 117927 6069
rect 1104 6010 118864 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 96374 6010
rect 96426 5958 96438 6010
rect 96490 5958 96502 6010
rect 96554 5958 96566 6010
rect 96618 5958 96630 6010
rect 96682 5958 118864 6010
rect 1104 5936 118864 5958
rect 117682 5652 117688 5704
rect 117740 5692 117746 5704
rect 117961 5695 118019 5701
rect 117961 5692 117973 5695
rect 117740 5664 117973 5692
rect 117740 5652 117746 5664
rect 117961 5661 117973 5664
rect 118007 5661 118019 5695
rect 117961 5655 118019 5661
rect 116302 5516 116308 5568
rect 116360 5556 116366 5568
rect 117777 5559 117835 5565
rect 117777 5556 117789 5559
rect 116360 5528 117789 5556
rect 116360 5516 116366 5528
rect 117777 5525 117789 5528
rect 117823 5525 117835 5559
rect 117777 5519 117835 5525
rect 1104 5466 118864 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 81014 5466
rect 81066 5414 81078 5466
rect 81130 5414 81142 5466
rect 81194 5414 81206 5466
rect 81258 5414 81270 5466
rect 81322 5414 111734 5466
rect 111786 5414 111798 5466
rect 111850 5414 111862 5466
rect 111914 5414 111926 5466
rect 111978 5414 111990 5466
rect 112042 5414 118864 5466
rect 1104 5392 118864 5414
rect 117774 5216 117780 5228
rect 117735 5188 117780 5216
rect 117774 5176 117780 5188
rect 117832 5176 117838 5228
rect 117866 5012 117872 5024
rect 117827 4984 117872 5012
rect 117866 4972 117872 4984
rect 117924 4972 117930 5024
rect 1104 4922 118864 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 96374 4922
rect 96426 4870 96438 4922
rect 96490 4870 96502 4922
rect 96554 4870 96566 4922
rect 96618 4870 96630 4922
rect 96682 4870 118864 4922
rect 1104 4848 118864 4870
rect 116397 4811 116455 4817
rect 116397 4777 116409 4811
rect 116443 4808 116455 4811
rect 117590 4808 117596 4820
rect 116443 4780 117596 4808
rect 116443 4777 116455 4780
rect 116397 4771 116455 4777
rect 117590 4768 117596 4780
rect 117648 4768 117654 4820
rect 116210 4604 116216 4616
rect 116171 4576 116216 4604
rect 116210 4564 116216 4576
rect 116268 4564 116274 4616
rect 117774 4536 117780 4548
rect 117735 4508 117780 4536
rect 117774 4496 117780 4508
rect 117832 4496 117838 4548
rect 97534 4428 97540 4480
rect 97592 4468 97598 4480
rect 104158 4468 104164 4480
rect 97592 4440 104164 4468
rect 97592 4428 97598 4440
rect 104158 4428 104164 4440
rect 104216 4428 104222 4480
rect 115290 4428 115296 4480
rect 115348 4468 115354 4480
rect 117869 4471 117927 4477
rect 117869 4468 117881 4471
rect 115348 4440 117881 4468
rect 115348 4428 115354 4440
rect 117869 4437 117881 4440
rect 117915 4437 117927 4471
rect 117869 4431 117927 4437
rect 1104 4378 118864 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 81014 4378
rect 81066 4326 81078 4378
rect 81130 4326 81142 4378
rect 81194 4326 81206 4378
rect 81258 4326 81270 4378
rect 81322 4326 111734 4378
rect 111786 4326 111798 4378
rect 111850 4326 111862 4378
rect 111914 4326 111926 4378
rect 111978 4326 111990 4378
rect 112042 4326 118864 4378
rect 1104 4304 118864 4326
rect 58250 4224 58256 4276
rect 58308 4264 58314 4276
rect 97534 4264 97540 4276
rect 58308 4236 97540 4264
rect 58308 4224 58314 4236
rect 97534 4224 97540 4236
rect 97592 4224 97598 4276
rect 97813 4267 97871 4273
rect 97813 4233 97825 4267
rect 97859 4264 97871 4267
rect 97994 4264 98000 4276
rect 97859 4236 98000 4264
rect 97859 4233 97871 4236
rect 97813 4227 97871 4233
rect 97994 4224 98000 4236
rect 98052 4224 98058 4276
rect 100386 4224 100392 4276
rect 100444 4264 100450 4276
rect 100665 4267 100723 4273
rect 100665 4264 100677 4267
rect 100444 4236 100677 4264
rect 100444 4224 100450 4236
rect 100665 4233 100677 4236
rect 100711 4233 100723 4267
rect 100665 4227 100723 4233
rect 104158 4224 104164 4276
rect 104216 4264 104222 4276
rect 116118 4264 116124 4276
rect 104216 4236 116124 4264
rect 104216 4224 104222 4236
rect 116118 4224 116124 4236
rect 116176 4224 116182 4276
rect 117498 4264 117504 4276
rect 116228 4236 117504 4264
rect 25682 4156 25688 4208
rect 25740 4196 25746 4208
rect 85022 4196 85028 4208
rect 25740 4168 85028 4196
rect 25740 4156 25746 4168
rect 85022 4156 85028 4168
rect 85080 4156 85086 4208
rect 97828 4168 98132 4196
rect 97828 4152 97856 4168
rect 67358 4088 67364 4140
rect 67416 4128 67422 4140
rect 97644 4128 97856 4152
rect 67416 4124 97856 4128
rect 67416 4100 97672 4124
rect 67416 4088 67422 4100
rect 97902 4088 97908 4140
rect 97960 4128 97966 4140
rect 97997 4131 98055 4137
rect 97997 4128 98009 4131
rect 97960 4100 98009 4128
rect 97960 4088 97966 4100
rect 97997 4097 98009 4100
rect 98043 4097 98055 4131
rect 98104 4128 98132 4168
rect 100772 4168 101076 4196
rect 100772 4128 100800 4168
rect 98104 4100 100800 4128
rect 97997 4091 98055 4097
rect 100846 4088 100852 4140
rect 100904 4128 100910 4140
rect 101048 4128 101076 4168
rect 114738 4156 114744 4208
rect 114796 4196 114802 4208
rect 116228 4196 116256 4236
rect 117498 4224 117504 4236
rect 117556 4224 117562 4276
rect 114796 4168 116256 4196
rect 114796 4156 114802 4168
rect 117222 4156 117228 4208
rect 117280 4196 117286 4208
rect 117777 4199 117835 4205
rect 117777 4196 117789 4199
rect 117280 4168 117789 4196
rect 117280 4156 117286 4168
rect 117777 4165 117789 4168
rect 117823 4165 117835 4199
rect 117777 4159 117835 4165
rect 100904 4100 100949 4128
rect 101048 4100 113496 4128
rect 100904 4088 100910 4100
rect 63126 4020 63132 4072
rect 63184 4060 63190 4072
rect 113358 4060 113364 4072
rect 63184 4032 113364 4060
rect 63184 4020 63190 4032
rect 113358 4020 113364 4032
rect 113416 4020 113422 4072
rect 113468 4060 113496 4100
rect 114830 4088 114836 4140
rect 114888 4128 114894 4140
rect 115109 4131 115167 4137
rect 115109 4128 115121 4131
rect 114888 4100 115121 4128
rect 114888 4088 114894 4100
rect 115109 4097 115121 4100
rect 115155 4097 115167 4131
rect 115842 4128 115848 4140
rect 115803 4100 115848 4128
rect 115109 4091 115167 4097
rect 115842 4088 115848 4100
rect 115900 4088 115906 4140
rect 116578 4128 116584 4140
rect 116539 4100 116584 4128
rect 116578 4088 116584 4100
rect 116636 4088 116642 4140
rect 116670 4088 116676 4140
rect 116728 4128 116734 4140
rect 118142 4128 118148 4140
rect 116728 4100 118148 4128
rect 116728 4088 116734 4100
rect 118142 4088 118148 4100
rect 118200 4088 118206 4140
rect 117866 4060 117872 4072
rect 113468 4032 117872 4060
rect 117866 4020 117872 4032
rect 117924 4020 117930 4072
rect 68830 3952 68836 4004
rect 68888 3992 68894 4004
rect 68888 3964 111656 3992
rect 68888 3952 68894 3964
rect 64966 3884 64972 3936
rect 65024 3924 65030 3936
rect 111518 3924 111524 3936
rect 65024 3896 111524 3924
rect 65024 3884 65030 3896
rect 111518 3884 111524 3896
rect 111576 3884 111582 3936
rect 111628 3924 111656 3964
rect 111702 3952 111708 4004
rect 111760 3992 111766 4004
rect 117961 3995 118019 4001
rect 117961 3992 117973 3995
rect 111760 3964 117973 3992
rect 111760 3952 111766 3964
rect 117961 3961 117973 3964
rect 118007 3961 118019 3995
rect 117961 3955 118019 3961
rect 114738 3924 114744 3936
rect 111628 3896 114744 3924
rect 114738 3884 114744 3896
rect 114796 3884 114802 3936
rect 114925 3927 114983 3933
rect 114925 3893 114937 3927
rect 114971 3924 114983 3927
rect 115382 3924 115388 3936
rect 114971 3896 115388 3924
rect 114971 3893 114983 3896
rect 114925 3887 114983 3893
rect 115382 3884 115388 3896
rect 115440 3884 115446 3936
rect 116029 3927 116087 3933
rect 116029 3893 116041 3927
rect 116075 3924 116087 3927
rect 116670 3924 116676 3936
rect 116075 3896 116676 3924
rect 116075 3893 116087 3896
rect 116029 3887 116087 3893
rect 116670 3884 116676 3896
rect 116728 3884 116734 3936
rect 116765 3927 116823 3933
rect 116765 3893 116777 3927
rect 116811 3924 116823 3927
rect 118418 3924 118424 3936
rect 116811 3896 118424 3924
rect 116811 3893 116823 3896
rect 116765 3887 116823 3893
rect 118418 3884 118424 3896
rect 118476 3884 118482 3936
rect 1104 3834 118864 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 96374 3834
rect 96426 3782 96438 3834
rect 96490 3782 96502 3834
rect 96554 3782 96566 3834
rect 96618 3782 96630 3834
rect 96682 3782 118864 3834
rect 1104 3760 118864 3782
rect 61654 3680 61660 3732
rect 61712 3720 61718 3732
rect 113266 3720 113272 3732
rect 61712 3692 113272 3720
rect 61712 3680 61718 3692
rect 113266 3680 113272 3692
rect 113324 3680 113330 3732
rect 113358 3680 113364 3732
rect 113416 3720 113422 3732
rect 117869 3723 117927 3729
rect 117869 3720 117881 3723
rect 113416 3692 117881 3720
rect 113416 3680 113422 3692
rect 117869 3689 117881 3692
rect 117915 3689 117927 3723
rect 117869 3683 117927 3689
rect 57146 3612 57152 3664
rect 57204 3652 57210 3664
rect 98638 3652 98644 3664
rect 57204 3624 98644 3652
rect 57204 3612 57210 3624
rect 98638 3612 98644 3624
rect 98696 3612 98702 3664
rect 98914 3612 98920 3664
rect 98972 3652 98978 3664
rect 99009 3655 99067 3661
rect 99009 3652 99021 3655
rect 98972 3624 99021 3652
rect 98972 3612 98978 3624
rect 99009 3621 99021 3624
rect 99055 3621 99067 3655
rect 105998 3652 106004 3664
rect 99009 3615 99067 3621
rect 99116 3624 101444 3652
rect 105959 3624 106004 3652
rect 45186 3544 45192 3596
rect 45244 3584 45250 3596
rect 98730 3584 98736 3596
rect 45244 3556 98736 3584
rect 45244 3544 45250 3556
rect 98730 3544 98736 3556
rect 98788 3544 98794 3596
rect 63126 3516 63132 3528
rect 63087 3488 63132 3516
rect 63126 3476 63132 3488
rect 63184 3476 63190 3528
rect 68278 3476 68284 3528
rect 68336 3516 68342 3528
rect 68373 3519 68431 3525
rect 68373 3516 68385 3519
rect 68336 3488 68385 3516
rect 68336 3476 68342 3488
rect 68373 3485 68385 3488
rect 68419 3516 68431 3519
rect 68830 3516 68836 3528
rect 68419 3488 68836 3516
rect 68419 3485 68431 3488
rect 68373 3479 68431 3485
rect 68830 3476 68836 3488
rect 68888 3476 68894 3528
rect 76282 3476 76288 3528
rect 76340 3516 76346 3528
rect 76561 3519 76619 3525
rect 76561 3516 76573 3519
rect 76340 3488 76573 3516
rect 76340 3476 76346 3488
rect 76561 3485 76573 3488
rect 76607 3485 76619 3519
rect 76561 3479 76619 3485
rect 81986 3476 81992 3528
rect 82044 3516 82050 3528
rect 82265 3519 82323 3525
rect 82265 3516 82277 3519
rect 82044 3488 82277 3516
rect 82044 3476 82050 3488
rect 82265 3485 82277 3488
rect 82311 3485 82323 3519
rect 82265 3479 82323 3485
rect 83458 3476 83464 3528
rect 83516 3516 83522 3528
rect 83737 3519 83795 3525
rect 83737 3516 83749 3519
rect 83516 3488 83749 3516
rect 83516 3476 83522 3488
rect 83737 3485 83749 3488
rect 83783 3485 83795 3519
rect 83737 3479 83795 3485
rect 84838 3476 84844 3528
rect 84896 3516 84902 3528
rect 85117 3519 85175 3525
rect 85117 3516 85129 3519
rect 84896 3488 85129 3516
rect 84896 3476 84902 3488
rect 85117 3485 85129 3488
rect 85163 3485 85175 3519
rect 85117 3479 85175 3485
rect 86310 3476 86316 3528
rect 86368 3516 86374 3528
rect 86589 3519 86647 3525
rect 86589 3516 86601 3519
rect 86368 3488 86601 3516
rect 86368 3476 86374 3488
rect 86589 3485 86601 3488
rect 86635 3485 86647 3519
rect 86589 3479 86647 3485
rect 87690 3476 87696 3528
rect 87748 3516 87754 3528
rect 87969 3519 88027 3525
rect 87969 3516 87981 3519
rect 87748 3488 87981 3516
rect 87748 3476 87754 3488
rect 87969 3485 87981 3488
rect 88015 3485 88027 3519
rect 87969 3479 88027 3485
rect 91741 3519 91799 3525
rect 91741 3485 91753 3519
rect 91787 3516 91799 3519
rect 92014 3516 92020 3528
rect 91787 3488 92020 3516
rect 91787 3485 91799 3488
rect 91741 3479 91799 3485
rect 92014 3476 92020 3488
rect 92072 3476 92078 3528
rect 92198 3516 92204 3528
rect 92159 3488 92204 3516
rect 92198 3476 92204 3488
rect 92256 3476 92262 3528
rect 96154 3476 96160 3528
rect 96212 3516 96218 3528
rect 96709 3519 96767 3525
rect 96709 3516 96721 3519
rect 96212 3488 96721 3516
rect 96212 3476 96218 3488
rect 96709 3485 96721 3488
rect 96755 3485 96767 3519
rect 96709 3479 96767 3485
rect 97718 3476 97724 3528
rect 97776 3516 97782 3528
rect 97905 3519 97963 3525
rect 97905 3516 97917 3519
rect 97776 3488 97917 3516
rect 97776 3476 97782 3488
rect 97905 3485 97917 3488
rect 97951 3485 97963 3519
rect 97905 3479 97963 3485
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99116 3516 99144 3624
rect 101416 3584 101444 3624
rect 105998 3612 106004 3624
rect 106056 3612 106062 3664
rect 106090 3612 106096 3664
rect 106148 3652 106154 3664
rect 107654 3652 107660 3664
rect 106148 3624 107660 3652
rect 106148 3612 106154 3624
rect 107654 3612 107660 3624
rect 107712 3612 107718 3664
rect 114922 3612 114928 3664
rect 114980 3652 114986 3664
rect 115753 3655 115811 3661
rect 114980 3624 115025 3652
rect 114980 3612 114986 3624
rect 115753 3621 115765 3655
rect 115799 3621 115811 3655
rect 115753 3615 115811 3621
rect 114002 3584 114008 3596
rect 101416 3556 114008 3584
rect 114002 3544 114008 3556
rect 114060 3544 114066 3596
rect 114094 3544 114100 3596
rect 114152 3584 114158 3596
rect 114152 3556 115152 3584
rect 114152 3544 114158 3556
rect 98696 3488 99144 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3528
rect 99340 3516 99346 3528
rect 99653 3519 99711 3525
rect 99653 3516 99665 3519
rect 99340 3488 99665 3516
rect 99340 3476 99346 3488
rect 99653 3485 99665 3488
rect 99699 3485 99711 3519
rect 99653 3479 99711 3485
rect 100294 3476 100300 3528
rect 100352 3516 100358 3528
rect 100389 3519 100447 3525
rect 100389 3516 100401 3519
rect 100352 3488 100401 3516
rect 100352 3476 100358 3488
rect 100389 3485 100401 3488
rect 100435 3485 100447 3519
rect 105814 3516 105820 3528
rect 105775 3488 105820 3516
rect 100389 3479 100447 3485
rect 105814 3476 105820 3488
rect 105872 3476 105878 3528
rect 106274 3476 106280 3528
rect 106332 3516 106338 3528
rect 107013 3519 107071 3525
rect 107013 3516 107025 3519
rect 106332 3488 107025 3516
rect 106332 3476 106338 3488
rect 107013 3485 107025 3488
rect 107059 3485 107071 3519
rect 112254 3516 112260 3528
rect 112215 3488 112260 3516
rect 107013 3479 107071 3485
rect 112254 3476 112260 3488
rect 112312 3476 112318 3528
rect 115124 3525 115152 3556
rect 115198 3544 115204 3596
rect 115256 3584 115262 3596
rect 115768 3584 115796 3615
rect 116394 3584 116400 3596
rect 115256 3556 115796 3584
rect 116355 3556 116400 3584
rect 115256 3544 115262 3556
rect 116394 3544 116400 3556
rect 116452 3544 116458 3596
rect 114741 3519 114799 3525
rect 114741 3485 114753 3519
rect 114787 3485 114799 3519
rect 114741 3479 114799 3485
rect 115109 3519 115167 3525
rect 115109 3485 115121 3519
rect 115155 3485 115167 3519
rect 116118 3516 116124 3528
rect 115109 3479 115167 3485
rect 115216 3488 115888 3516
rect 116079 3488 116124 3516
rect 65518 3408 65524 3460
rect 65576 3448 65582 3460
rect 76190 3448 76196 3460
rect 65576 3420 76196 3448
rect 65576 3408 65582 3420
rect 76190 3408 76196 3420
rect 76248 3408 76254 3460
rect 88886 3408 88892 3460
rect 88944 3448 88950 3460
rect 97626 3448 97632 3460
rect 88944 3420 97632 3448
rect 88944 3408 88950 3420
rect 97626 3408 97632 3420
rect 97684 3408 97690 3460
rect 98825 3451 98883 3457
rect 98825 3417 98837 3451
rect 98871 3448 98883 3451
rect 99098 3448 99104 3460
rect 98871 3420 99104 3448
rect 98871 3417 98883 3420
rect 98825 3411 98883 3417
rect 99098 3408 99104 3420
rect 99156 3408 99162 3460
rect 99558 3408 99564 3460
rect 99616 3448 99622 3460
rect 114756 3448 114784 3479
rect 114922 3448 114928 3460
rect 99616 3420 112208 3448
rect 114756 3420 114928 3448
rect 99616 3408 99622 3420
rect 62945 3383 63003 3389
rect 62945 3349 62957 3383
rect 62991 3380 63003 3383
rect 63586 3380 63592 3392
rect 62991 3352 63592 3380
rect 62991 3349 63003 3352
rect 62945 3343 63003 3349
rect 63586 3340 63592 3352
rect 63644 3340 63650 3392
rect 68649 3383 68707 3389
rect 68649 3349 68661 3383
rect 68695 3380 68707 3383
rect 69106 3380 69112 3392
rect 68695 3352 69112 3380
rect 68695 3349 68707 3352
rect 68649 3343 68707 3349
rect 69106 3340 69112 3352
rect 69164 3340 69170 3392
rect 76377 3383 76435 3389
rect 76377 3349 76389 3383
rect 76423 3380 76435 3383
rect 76466 3380 76472 3392
rect 76423 3352 76472 3380
rect 76423 3349 76435 3352
rect 76377 3343 76435 3349
rect 76466 3340 76472 3352
rect 76524 3340 76530 3392
rect 82081 3383 82139 3389
rect 82081 3349 82093 3383
rect 82127 3380 82139 3383
rect 83090 3380 83096 3392
rect 82127 3352 83096 3380
rect 82127 3349 82139 3352
rect 82081 3343 82139 3349
rect 83090 3340 83096 3352
rect 83148 3340 83154 3392
rect 83550 3380 83556 3392
rect 83511 3352 83556 3380
rect 83550 3340 83556 3352
rect 83608 3340 83614 3392
rect 84930 3380 84936 3392
rect 84891 3352 84936 3380
rect 84930 3340 84936 3352
rect 84988 3340 84994 3392
rect 86402 3380 86408 3392
rect 86363 3352 86408 3380
rect 86402 3340 86408 3352
rect 86460 3340 86466 3392
rect 87782 3380 87788 3392
rect 87743 3352 87788 3380
rect 87782 3340 87788 3352
rect 87840 3340 87846 3392
rect 91554 3380 91560 3392
rect 91515 3352 91560 3380
rect 91554 3340 91560 3352
rect 91612 3340 91618 3392
rect 92382 3380 92388 3392
rect 92343 3352 92388 3380
rect 92382 3340 92388 3352
rect 92440 3340 92446 3392
rect 96525 3383 96583 3389
rect 96525 3349 96537 3383
rect 96571 3380 96583 3383
rect 96982 3380 96988 3392
rect 96571 3352 96988 3380
rect 96571 3349 96583 3352
rect 96525 3343 96583 3349
rect 96982 3340 96988 3352
rect 97040 3340 97046 3392
rect 98086 3380 98092 3392
rect 98047 3352 98092 3380
rect 98086 3340 98092 3352
rect 98144 3340 98150 3392
rect 99834 3340 99840 3392
rect 99892 3380 99898 3392
rect 99892 3352 99937 3380
rect 99892 3340 99898 3352
rect 100570 3340 100576 3392
rect 100628 3380 100634 3392
rect 100628 3352 100673 3380
rect 100628 3340 100634 3352
rect 100754 3340 100760 3392
rect 100812 3380 100818 3392
rect 105998 3380 106004 3392
rect 100812 3352 106004 3380
rect 100812 3340 100818 3352
rect 105998 3340 106004 3352
rect 106056 3340 106062 3392
rect 106090 3340 106096 3392
rect 106148 3380 106154 3392
rect 106829 3383 106887 3389
rect 106829 3380 106841 3383
rect 106148 3352 106841 3380
rect 106148 3340 106154 3352
rect 106829 3349 106841 3352
rect 106875 3349 106887 3383
rect 112070 3380 112076 3392
rect 112031 3352 112076 3380
rect 106829 3343 106887 3349
rect 112070 3340 112076 3352
rect 112128 3340 112134 3392
rect 112180 3380 112208 3420
rect 114922 3408 114928 3420
rect 114980 3408 114986 3460
rect 115216 3380 115244 3488
rect 115860 3448 115888 3488
rect 116118 3476 116124 3488
rect 116176 3476 116182 3528
rect 116213 3519 116271 3525
rect 116213 3485 116225 3519
rect 116259 3516 116271 3519
rect 116302 3516 116308 3528
rect 116259 3488 116308 3516
rect 116259 3485 116271 3488
rect 116213 3479 116271 3485
rect 116302 3476 116308 3488
rect 116360 3476 116366 3528
rect 116854 3448 116860 3460
rect 115860 3420 116860 3448
rect 116854 3408 116860 3420
rect 116912 3408 116918 3460
rect 117130 3408 117136 3460
rect 117188 3448 117194 3460
rect 117777 3451 117835 3457
rect 117777 3448 117789 3451
rect 117188 3420 117789 3448
rect 117188 3408 117194 3420
rect 117777 3417 117789 3420
rect 117823 3417 117835 3451
rect 117777 3411 117835 3417
rect 112180 3352 115244 3380
rect 115293 3383 115351 3389
rect 115293 3349 115305 3383
rect 115339 3380 115351 3383
rect 117958 3380 117964 3392
rect 115339 3352 117964 3380
rect 115339 3349 115351 3352
rect 115293 3343 115351 3349
rect 117958 3340 117964 3352
rect 118016 3340 118022 3392
rect 1104 3290 118864 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 81014 3290
rect 81066 3238 81078 3290
rect 81130 3238 81142 3290
rect 81194 3238 81206 3290
rect 81258 3238 81270 3290
rect 81322 3238 111734 3290
rect 111786 3238 111798 3290
rect 111850 3238 111862 3290
rect 111914 3238 111926 3290
rect 111978 3238 111990 3290
rect 112042 3238 118864 3290
rect 1104 3216 118864 3238
rect 17034 3136 17040 3188
rect 17092 3176 17098 3188
rect 65518 3176 65524 3188
rect 17092 3148 65524 3176
rect 17092 3136 17098 3148
rect 65518 3136 65524 3148
rect 65576 3136 65582 3188
rect 65797 3179 65855 3185
rect 65797 3145 65809 3179
rect 65843 3145 65855 3179
rect 76650 3176 76656 3188
rect 76611 3148 76656 3176
rect 65797 3139 65855 3145
rect 61378 3108 61384 3120
rect 60292 3080 61384 3108
rect 54846 3000 54852 3052
rect 54904 3040 54910 3052
rect 55401 3043 55459 3049
rect 55401 3040 55413 3043
rect 54904 3012 55413 3040
rect 54904 3000 54910 3012
rect 55401 3009 55413 3012
rect 55447 3009 55459 3043
rect 55401 3003 55459 3009
rect 59170 3000 59176 3052
rect 59228 3040 59234 3052
rect 59265 3043 59323 3049
rect 59265 3040 59277 3043
rect 59228 3012 59277 3040
rect 59228 3000 59234 3012
rect 59265 3009 59277 3012
rect 59311 3009 59323 3043
rect 59265 3003 59323 3009
rect 59538 3000 59544 3052
rect 59596 3040 59602 3052
rect 60292 3049 60320 3080
rect 61378 3068 61384 3080
rect 61436 3068 61442 3120
rect 65812 3108 65840 3139
rect 76650 3136 76656 3148
rect 76708 3136 76714 3188
rect 78674 3176 78680 3188
rect 78635 3148 78680 3176
rect 78674 3136 78680 3148
rect 78732 3136 78738 3188
rect 79594 3176 79600 3188
rect 79555 3148 79600 3176
rect 79594 3136 79600 3148
rect 79652 3136 79658 3188
rect 81710 3176 81716 3188
rect 81671 3148 81716 3176
rect 81710 3136 81716 3148
rect 81768 3136 81774 3188
rect 82814 3176 82820 3188
rect 82775 3148 82820 3176
rect 82814 3136 82820 3148
rect 82872 3136 82878 3188
rect 85206 3176 85212 3188
rect 85167 3148 85212 3176
rect 85206 3136 85212 3148
rect 85264 3136 85270 3188
rect 86678 3176 86684 3188
rect 86639 3148 86684 3176
rect 86678 3136 86684 3148
rect 86736 3136 86742 3188
rect 92566 3176 92572 3188
rect 87432 3148 92572 3176
rect 70118 3108 70124 3120
rect 65812 3080 66300 3108
rect 60277 3043 60335 3049
rect 60277 3040 60289 3043
rect 59596 3012 60289 3040
rect 59596 3000 59602 3012
rect 60277 3009 60289 3012
rect 60323 3009 60335 3043
rect 60277 3003 60335 3009
rect 60737 3043 60795 3049
rect 60737 3009 60749 3043
rect 60783 3009 60795 3043
rect 60737 3003 60795 3009
rect 60752 2972 60780 3003
rect 61010 3000 61016 3052
rect 61068 3040 61074 3052
rect 61654 3040 61660 3052
rect 61068 3012 61660 3040
rect 61068 3000 61074 3012
rect 61654 3000 61660 3012
rect 61712 3000 61718 3052
rect 63586 3040 63592 3052
rect 63547 3012 63592 3040
rect 63586 3000 63592 3012
rect 63644 3000 63650 3052
rect 64874 3040 64880 3052
rect 64835 3012 64880 3040
rect 64874 3000 64880 3012
rect 64932 3000 64938 3052
rect 66272 3049 66300 3080
rect 66364 3080 70124 3108
rect 65981 3043 66039 3049
rect 65981 3009 65993 3043
rect 66027 3009 66039 3043
rect 65981 3003 66039 3009
rect 66257 3043 66315 3049
rect 66257 3009 66269 3043
rect 66303 3009 66315 3043
rect 66257 3003 66315 3009
rect 60108 2944 60780 2972
rect 51902 2864 51908 2916
rect 51960 2904 51966 2916
rect 56686 2904 56692 2916
rect 51960 2876 56692 2904
rect 51960 2864 51966 2876
rect 56686 2864 56692 2876
rect 56744 2864 56750 2916
rect 60108 2913 60136 2944
rect 64414 2932 64420 2984
rect 64472 2972 64478 2984
rect 64966 2972 64972 2984
rect 64472 2944 64972 2972
rect 64472 2932 64478 2944
rect 64966 2932 64972 2944
rect 65024 2932 65030 2984
rect 65518 2972 65524 2984
rect 65431 2944 65524 2972
rect 65518 2932 65524 2944
rect 65576 2972 65582 2984
rect 65996 2972 66024 3003
rect 66364 2972 66392 3080
rect 70118 3068 70124 3080
rect 70176 3068 70182 3120
rect 87432 3108 87460 3148
rect 92566 3136 92572 3148
rect 92624 3136 92630 3188
rect 92661 3179 92719 3185
rect 92661 3145 92673 3179
rect 92707 3176 92719 3179
rect 93946 3176 93952 3188
rect 92707 3148 93952 3176
rect 92707 3145 92719 3148
rect 92661 3139 92719 3145
rect 93946 3136 93952 3148
rect 94004 3136 94010 3188
rect 95970 3176 95976 3188
rect 95931 3148 95976 3176
rect 95970 3136 95976 3148
rect 96028 3136 96034 3188
rect 96709 3179 96767 3185
rect 96709 3145 96721 3179
rect 96755 3176 96767 3179
rect 96890 3176 96896 3188
rect 96755 3148 96896 3176
rect 96755 3145 96767 3148
rect 96709 3139 96767 3145
rect 96890 3136 96896 3148
rect 96948 3136 96954 3188
rect 99101 3179 99159 3185
rect 99101 3145 99113 3179
rect 99147 3176 99159 3179
rect 99282 3176 99288 3188
rect 99147 3148 99288 3176
rect 99147 3145 99159 3148
rect 99101 3139 99159 3145
rect 99282 3136 99288 3148
rect 99340 3136 99346 3188
rect 99561 3179 99619 3185
rect 99561 3145 99573 3179
rect 99607 3176 99619 3179
rect 101033 3179 101091 3185
rect 101033 3176 101045 3179
rect 99607 3148 101045 3176
rect 99607 3145 99619 3148
rect 99561 3139 99619 3145
rect 101033 3145 101045 3148
rect 101079 3145 101091 3179
rect 102410 3176 102416 3188
rect 102371 3148 102416 3176
rect 101033 3139 101091 3145
rect 102410 3136 102416 3148
rect 102468 3136 102474 3188
rect 104434 3176 104440 3188
rect 104395 3148 104440 3176
rect 104434 3136 104440 3148
rect 104492 3136 104498 3188
rect 106090 3176 106096 3188
rect 106051 3148 106096 3176
rect 106090 3136 106096 3148
rect 106148 3136 106154 3188
rect 107013 3179 107071 3185
rect 107013 3145 107025 3179
rect 107059 3176 107071 3179
rect 107102 3176 107108 3188
rect 107059 3148 107108 3176
rect 107059 3145 107071 3148
rect 107013 3139 107071 3145
rect 107102 3136 107108 3148
rect 107160 3136 107166 3188
rect 108482 3176 108488 3188
rect 108443 3148 108488 3176
rect 108482 3136 108488 3148
rect 108540 3136 108546 3188
rect 110782 3176 110788 3188
rect 109006 3148 110552 3176
rect 110743 3148 110788 3176
rect 70366 3080 87460 3108
rect 87509 3111 87567 3117
rect 66714 3000 66720 3052
rect 66772 3040 66778 3052
rect 66901 3043 66959 3049
rect 66901 3040 66913 3043
rect 66772 3012 66913 3040
rect 66772 3000 66778 3012
rect 66901 3009 66913 3012
rect 66947 3040 66959 3043
rect 67358 3040 67364 3052
rect 66947 3012 67364 3040
rect 66947 3009 66959 3012
rect 66901 3003 66959 3009
rect 67358 3000 67364 3012
rect 67416 3000 67422 3052
rect 68189 3043 68247 3049
rect 68189 3009 68201 3043
rect 68235 3009 68247 3043
rect 69106 3040 69112 3052
rect 69067 3012 69112 3040
rect 68189 3003 68247 3009
rect 68204 2972 68232 3003
rect 69106 3000 69112 3012
rect 69164 3000 69170 3052
rect 70213 3043 70271 3049
rect 70213 3040 70225 3043
rect 69676 3012 70225 3040
rect 65576 2944 66392 2972
rect 67192 2944 68232 2972
rect 65576 2932 65582 2944
rect 60093 2907 60151 2913
rect 60093 2873 60105 2907
rect 60139 2873 60151 2907
rect 66162 2904 66168 2916
rect 60093 2867 60151 2873
rect 60200 2876 66168 2904
rect 55677 2839 55735 2845
rect 55677 2805 55689 2839
rect 55723 2836 55735 2839
rect 56502 2836 56508 2848
rect 55723 2808 56508 2836
rect 55723 2805 55735 2808
rect 55677 2799 55735 2805
rect 56502 2796 56508 2808
rect 56560 2796 56566 2848
rect 59449 2839 59507 2845
rect 59449 2805 59461 2839
rect 59495 2836 59507 2839
rect 60200 2836 60228 2876
rect 66162 2864 66168 2876
rect 66220 2864 66226 2916
rect 67192 2913 67220 2944
rect 67177 2907 67235 2913
rect 67177 2873 67189 2907
rect 67223 2873 67235 2907
rect 67177 2867 67235 2873
rect 59495 2808 60228 2836
rect 60921 2839 60979 2845
rect 59495 2805 59507 2808
rect 59449 2799 59507 2805
rect 60921 2805 60933 2839
rect 60967 2836 60979 2839
rect 61102 2836 61108 2848
rect 60967 2808 61108 2836
rect 60967 2805 60979 2808
rect 60921 2799 60979 2805
rect 61102 2796 61108 2808
rect 61160 2796 61166 2848
rect 61473 2839 61531 2845
rect 61473 2805 61485 2839
rect 61519 2836 61531 2839
rect 62114 2836 62120 2848
rect 61519 2808 62120 2836
rect 61519 2805 61531 2808
rect 61473 2799 61531 2805
rect 62114 2796 62120 2808
rect 62172 2796 62178 2848
rect 63494 2796 63500 2848
rect 63552 2836 63558 2848
rect 63773 2839 63831 2845
rect 63773 2836 63785 2839
rect 63552 2808 63785 2836
rect 63552 2796 63558 2808
rect 63773 2805 63785 2808
rect 63819 2805 63831 2839
rect 63773 2799 63831 2805
rect 64966 2796 64972 2848
rect 65024 2836 65030 2848
rect 65061 2839 65119 2845
rect 65061 2836 65073 2839
rect 65024 2808 65073 2836
rect 65024 2796 65030 2808
rect 65061 2805 65073 2808
rect 65107 2805 65119 2839
rect 65061 2799 65119 2805
rect 66346 2796 66352 2848
rect 66404 2836 66410 2848
rect 66441 2839 66499 2845
rect 66441 2836 66453 2839
rect 66404 2808 66453 2836
rect 66404 2796 66410 2808
rect 66441 2805 66453 2808
rect 66487 2805 66499 2839
rect 66441 2799 66499 2805
rect 67726 2796 67732 2848
rect 67784 2836 67790 2848
rect 68373 2839 68431 2845
rect 68373 2836 68385 2839
rect 67784 2808 68385 2836
rect 67784 2796 67790 2808
rect 68373 2805 68385 2808
rect 68419 2805 68431 2839
rect 68373 2799 68431 2805
rect 69198 2796 69204 2848
rect 69256 2836 69262 2848
rect 69293 2839 69351 2845
rect 69293 2836 69305 2839
rect 69256 2808 69305 2836
rect 69256 2796 69262 2808
rect 69293 2805 69305 2808
rect 69339 2805 69351 2839
rect 69293 2799 69351 2805
rect 69566 2796 69572 2848
rect 69624 2836 69630 2848
rect 69676 2845 69704 3012
rect 70213 3009 70225 3012
rect 70259 3040 70271 3043
rect 70366 3040 70394 3080
rect 87509 3077 87521 3111
rect 87555 3108 87567 3111
rect 88886 3108 88892 3120
rect 87555 3080 88892 3108
rect 87555 3077 87567 3080
rect 87509 3071 87567 3077
rect 88886 3068 88892 3080
rect 88944 3068 88950 3120
rect 99650 3108 99656 3120
rect 88996 3080 99656 3108
rect 70259 3012 70394 3040
rect 70673 3043 70731 3049
rect 70259 3009 70271 3012
rect 70213 3003 70271 3009
rect 70673 3009 70685 3043
rect 70719 3009 70731 3043
rect 71682 3040 71688 3052
rect 71643 3012 71688 3040
rect 70673 3003 70731 3009
rect 70688 2972 70716 3003
rect 71682 3000 71688 3012
rect 71740 3000 71746 3052
rect 72145 3043 72203 3049
rect 72145 3009 72157 3043
rect 72191 3009 72203 3043
rect 73522 3040 73528 3052
rect 73483 3012 73528 3040
rect 72145 3003 72203 3009
rect 72160 2972 72188 3003
rect 73522 3000 73528 3012
rect 73580 3000 73586 3052
rect 74902 3000 74908 3052
rect 74960 3040 74966 3052
rect 75181 3043 75239 3049
rect 75181 3040 75193 3043
rect 74960 3012 75193 3040
rect 74960 3000 74966 3012
rect 75181 3009 75193 3012
rect 75227 3009 75239 3043
rect 76558 3040 76564 3052
rect 76519 3012 76564 3040
rect 75181 3003 75239 3009
rect 76558 3000 76564 3012
rect 76616 3000 76622 3052
rect 77754 3000 77760 3052
rect 77812 3040 77818 3052
rect 77941 3043 77999 3049
rect 77941 3040 77953 3043
rect 77812 3012 77953 3040
rect 77812 3000 77818 3012
rect 77941 3009 77953 3012
rect 77987 3009 77999 3043
rect 78582 3040 78588 3052
rect 78543 3012 78588 3040
rect 77941 3003 77999 3009
rect 78582 3000 78588 3012
rect 78640 3000 78646 3052
rect 79502 3040 79508 3052
rect 79463 3012 79508 3040
rect 79502 3000 79508 3012
rect 79560 3000 79566 3052
rect 80606 3000 80612 3052
rect 80664 3040 80670 3052
rect 80885 3043 80943 3049
rect 80885 3040 80897 3043
rect 80664 3012 80897 3040
rect 80664 3000 80670 3012
rect 80885 3009 80897 3012
rect 80931 3009 80943 3043
rect 81618 3040 81624 3052
rect 81579 3012 81624 3040
rect 80885 3003 80943 3009
rect 81618 3000 81624 3012
rect 81676 3000 81682 3052
rect 82538 3040 82544 3052
rect 82499 3012 82544 3040
rect 82538 3000 82544 3012
rect 82596 3000 82602 3052
rect 83734 3040 83740 3052
rect 83695 3012 83740 3040
rect 83734 3000 83740 3012
rect 83792 3000 83798 3052
rect 85114 3040 85120 3052
rect 85075 3012 85120 3040
rect 85114 3000 85120 3012
rect 85172 3000 85178 3052
rect 86586 3040 86592 3052
rect 86547 3012 86592 3040
rect 86586 3000 86592 3012
rect 86644 3000 86650 3052
rect 70044 2944 70716 2972
rect 71516 2944 72188 2972
rect 84013 2975 84071 2981
rect 70044 2913 70072 2944
rect 70029 2907 70087 2913
rect 70029 2873 70041 2907
rect 70075 2873 70087 2907
rect 70029 2867 70087 2873
rect 70118 2864 70124 2916
rect 70176 2904 70182 2916
rect 71516 2913 71544 2944
rect 84013 2941 84025 2975
rect 84059 2972 84071 2975
rect 88996 2972 89024 3080
rect 99650 3068 99656 3080
rect 99708 3068 99714 3120
rect 100570 3068 100576 3120
rect 100628 3108 100634 3120
rect 109006 3108 109034 3148
rect 100628 3080 109034 3108
rect 109773 3111 109831 3117
rect 100628 3068 100634 3080
rect 109773 3077 109785 3111
rect 109819 3108 109831 3111
rect 110417 3111 110475 3117
rect 110417 3108 110429 3111
rect 109819 3080 110429 3108
rect 109819 3077 109831 3080
rect 109773 3071 109831 3077
rect 110417 3077 110429 3080
rect 110463 3077 110475 3111
rect 110524 3108 110552 3148
rect 110782 3136 110788 3148
rect 110840 3136 110846 3188
rect 111889 3179 111947 3185
rect 111889 3145 111901 3179
rect 111935 3176 111947 3179
rect 112162 3176 112168 3188
rect 111935 3148 112168 3176
rect 111935 3145 111947 3148
rect 111889 3139 111947 3145
rect 112162 3136 112168 3148
rect 112220 3136 112226 3188
rect 114002 3136 114008 3188
rect 114060 3176 114066 3188
rect 115109 3179 115167 3185
rect 115109 3176 115121 3179
rect 114060 3148 115121 3176
rect 114060 3136 114066 3148
rect 115109 3145 115121 3148
rect 115155 3176 115167 3179
rect 115477 3179 115535 3185
rect 115477 3176 115489 3179
rect 115155 3148 115489 3176
rect 115155 3145 115167 3148
rect 115109 3139 115167 3145
rect 115477 3145 115489 3148
rect 115523 3145 115535 3179
rect 115477 3139 115535 3145
rect 115845 3179 115903 3185
rect 115845 3145 115857 3179
rect 115891 3176 115903 3179
rect 116210 3176 116216 3188
rect 115891 3148 116216 3176
rect 115891 3145 115903 3148
rect 115845 3139 115903 3145
rect 110524 3080 115428 3108
rect 110417 3071 110475 3077
rect 89162 3000 89168 3052
rect 89220 3040 89226 3052
rect 89717 3043 89775 3049
rect 89717 3040 89729 3043
rect 89220 3012 89729 3040
rect 89220 3000 89226 3012
rect 89717 3009 89729 3012
rect 89763 3009 89775 3043
rect 89717 3003 89775 3009
rect 90634 3000 90640 3052
rect 90692 3040 90698 3052
rect 90913 3043 90971 3049
rect 90913 3040 90925 3043
rect 90692 3012 90925 3040
rect 90692 3000 90698 3012
rect 90913 3009 90925 3012
rect 90959 3009 90971 3043
rect 90913 3003 90971 3009
rect 91462 3000 91468 3052
rect 91520 3040 91526 3052
rect 92566 3040 92572 3052
rect 91520 3012 92572 3040
rect 91520 3000 91526 3012
rect 92566 3000 92572 3012
rect 92624 3000 92630 3052
rect 92658 3000 92664 3052
rect 92716 3040 92722 3052
rect 92716 3012 93854 3040
rect 92716 3000 92722 3012
rect 84059 2944 89024 2972
rect 89073 2975 89131 2981
rect 84059 2941 84071 2944
rect 84013 2935 84071 2941
rect 89073 2941 89085 2975
rect 89119 2972 89131 2975
rect 89438 2972 89444 2984
rect 89119 2944 89444 2972
rect 89119 2941 89131 2944
rect 89073 2935 89131 2941
rect 89438 2932 89444 2944
rect 89496 2932 89502 2984
rect 92290 2932 92296 2984
rect 92348 2972 92354 2984
rect 92753 2975 92811 2981
rect 92753 2972 92765 2975
rect 92348 2944 92765 2972
rect 92348 2932 92354 2944
rect 92753 2941 92765 2944
rect 92799 2941 92811 2975
rect 92753 2935 92811 2941
rect 92842 2932 92848 2984
rect 92900 2972 92906 2984
rect 93213 2975 93271 2981
rect 93213 2972 93225 2975
rect 92900 2944 93225 2972
rect 92900 2932 92906 2944
rect 93213 2941 93225 2944
rect 93259 2941 93271 2975
rect 93826 2972 93854 3012
rect 94866 3000 94872 3052
rect 94924 3040 94930 3052
rect 95145 3043 95203 3049
rect 95145 3040 95157 3043
rect 94924 3012 95157 3040
rect 94924 3000 94930 3012
rect 95145 3009 95157 3012
rect 95191 3009 95203 3043
rect 95786 3040 95792 3052
rect 95747 3012 95792 3040
rect 95145 3003 95203 3009
rect 95786 3000 95792 3012
rect 95844 3000 95850 3052
rect 96246 3000 96252 3052
rect 96304 3040 96310 3052
rect 96525 3043 96583 3049
rect 96525 3040 96537 3043
rect 96304 3012 96537 3040
rect 96304 3000 96310 3012
rect 96525 3009 96537 3012
rect 96571 3009 96583 3043
rect 97626 3040 97632 3052
rect 97587 3012 97632 3040
rect 96525 3003 96583 3009
rect 97626 3000 97632 3012
rect 97684 3000 97690 3052
rect 98273 3043 98331 3049
rect 98273 3009 98285 3043
rect 98319 3040 98331 3043
rect 98638 3040 98644 3052
rect 98319 3012 98644 3040
rect 98319 3009 98331 3012
rect 98273 3003 98331 3009
rect 98638 3000 98644 3012
rect 98696 3000 98702 3052
rect 99466 3000 99472 3052
rect 99524 3040 99530 3052
rect 100113 3043 100171 3049
rect 100113 3040 100125 3043
rect 99524 3012 100125 3040
rect 99524 3000 99530 3012
rect 100113 3009 100125 3012
rect 100159 3009 100171 3043
rect 100113 3003 100171 3009
rect 100389 3044 100447 3049
rect 100389 3043 100524 3044
rect 100389 3009 100401 3043
rect 100435 3016 100524 3043
rect 101214 3040 101220 3052
rect 100435 3009 100447 3016
rect 100389 3003 100447 3009
rect 99558 2972 99564 2984
rect 93826 2944 99564 2972
rect 93213 2935 93271 2941
rect 99558 2932 99564 2944
rect 99616 2932 99622 2984
rect 99742 2972 99748 2984
rect 99703 2944 99748 2972
rect 99742 2932 99748 2944
rect 99800 2932 99806 2984
rect 100496 2972 100524 3016
rect 101175 3012 101220 3040
rect 101214 3000 101220 3012
rect 101272 3000 101278 3052
rect 102134 3000 102140 3052
rect 102192 3040 102198 3052
rect 102229 3043 102287 3049
rect 102229 3040 102241 3043
rect 102192 3012 102241 3040
rect 102192 3000 102198 3012
rect 102229 3009 102241 3012
rect 102275 3009 102287 3043
rect 102229 3003 102287 3009
rect 103149 3043 103207 3049
rect 103149 3009 103161 3043
rect 103195 3009 103207 3043
rect 104250 3040 104256 3052
rect 104211 3012 104256 3040
rect 103149 3003 103207 3009
rect 100754 2972 100760 2984
rect 100496 2944 100760 2972
rect 100754 2932 100760 2944
rect 100812 2932 100818 2984
rect 102042 2932 102048 2984
rect 102100 2972 102106 2984
rect 103164 2972 103192 3003
rect 104250 3000 104256 3012
rect 104308 3000 104314 3052
rect 104894 3000 104900 3052
rect 104952 3040 104958 3052
rect 104989 3043 105047 3049
rect 104989 3040 105001 3043
rect 104952 3012 105001 3040
rect 104952 3000 104958 3012
rect 104989 3009 105001 3012
rect 105035 3009 105047 3043
rect 104989 3003 105047 3009
rect 105262 3000 105268 3052
rect 105320 3040 105326 3052
rect 105357 3043 105415 3049
rect 105357 3040 105369 3043
rect 105320 3012 105369 3040
rect 105320 3000 105326 3012
rect 105357 3009 105369 3012
rect 105403 3040 105415 3043
rect 106001 3043 106059 3049
rect 106001 3040 106013 3043
rect 105403 3012 106013 3040
rect 105403 3009 105415 3012
rect 105357 3003 105415 3009
rect 106001 3009 106013 3012
rect 106047 3009 106059 3043
rect 106001 3003 106059 3009
rect 106829 3043 106887 3049
rect 106829 3009 106841 3043
rect 106875 3009 106887 3043
rect 106829 3003 106887 3009
rect 102100 2944 103192 2972
rect 102100 2932 102106 2944
rect 106182 2932 106188 2984
rect 106240 2972 106246 2984
rect 106240 2944 106285 2972
rect 106240 2932 106246 2944
rect 71501 2907 71559 2913
rect 70176 2876 70992 2904
rect 70176 2864 70182 2876
rect 69661 2839 69719 2845
rect 69661 2836 69673 2839
rect 69624 2808 69673 2836
rect 69624 2796 69630 2808
rect 69661 2805 69673 2808
rect 69707 2805 69719 2839
rect 69661 2799 69719 2805
rect 70578 2796 70584 2848
rect 70636 2836 70642 2848
rect 70857 2839 70915 2845
rect 70857 2836 70869 2839
rect 70636 2808 70869 2836
rect 70636 2796 70642 2808
rect 70857 2805 70869 2808
rect 70903 2805 70915 2839
rect 70964 2836 70992 2876
rect 71501 2873 71513 2907
rect 71547 2873 71559 2907
rect 105633 2907 105691 2913
rect 71501 2867 71559 2873
rect 71608 2876 105308 2904
rect 71608 2836 71636 2876
rect 70964 2808 71636 2836
rect 70857 2799 70915 2805
rect 72050 2796 72056 2848
rect 72108 2836 72114 2848
rect 72329 2839 72387 2845
rect 72329 2836 72341 2839
rect 72108 2808 72341 2836
rect 72108 2796 72114 2808
rect 72329 2805 72341 2808
rect 72375 2805 72387 2839
rect 72329 2799 72387 2805
rect 73341 2839 73399 2845
rect 73341 2805 73353 2839
rect 73387 2836 73399 2839
rect 73522 2836 73528 2848
rect 73387 2808 73528 2836
rect 73387 2805 73399 2808
rect 73341 2799 73399 2805
rect 73522 2796 73528 2808
rect 73580 2796 73586 2848
rect 74994 2836 75000 2848
rect 74955 2808 75000 2836
rect 74994 2796 75000 2808
rect 75052 2796 75058 2848
rect 77662 2796 77668 2848
rect 77720 2836 77726 2848
rect 77757 2839 77815 2845
rect 77757 2836 77769 2839
rect 77720 2808 77769 2836
rect 77720 2796 77726 2808
rect 77757 2805 77769 2808
rect 77803 2805 77815 2839
rect 77757 2799 77815 2805
rect 80701 2839 80759 2845
rect 80701 2805 80713 2839
rect 80747 2836 80759 2839
rect 81526 2836 81532 2848
rect 80747 2808 81532 2836
rect 80747 2805 80759 2808
rect 80701 2799 80759 2805
rect 81526 2796 81532 2808
rect 81584 2796 81590 2848
rect 86862 2796 86868 2848
rect 86920 2836 86926 2848
rect 87601 2839 87659 2845
rect 87601 2836 87613 2839
rect 86920 2808 87613 2836
rect 86920 2796 86926 2808
rect 87601 2805 87613 2808
rect 87647 2805 87659 2839
rect 87601 2799 87659 2805
rect 89254 2796 89260 2848
rect 89312 2836 89318 2848
rect 89533 2839 89591 2845
rect 89533 2836 89545 2839
rect 89312 2808 89545 2836
rect 89312 2796 89318 2808
rect 89533 2805 89545 2808
rect 89579 2805 89591 2839
rect 89533 2799 89591 2805
rect 90542 2796 90548 2848
rect 90600 2836 90606 2848
rect 90729 2839 90787 2845
rect 90729 2836 90741 2839
rect 90600 2808 90741 2836
rect 90600 2796 90606 2808
rect 90729 2805 90741 2808
rect 90775 2805 90787 2839
rect 91462 2836 91468 2848
rect 91423 2808 91468 2836
rect 90729 2799 90787 2805
rect 91462 2796 91468 2808
rect 91520 2836 91526 2848
rect 91833 2839 91891 2845
rect 91833 2836 91845 2839
rect 91520 2808 91845 2836
rect 91520 2796 91526 2808
rect 91833 2805 91845 2808
rect 91879 2805 91891 2839
rect 91833 2799 91891 2805
rect 92201 2839 92259 2845
rect 92201 2805 92213 2839
rect 92247 2836 92259 2839
rect 92934 2836 92940 2848
rect 92247 2808 92940 2836
rect 92247 2805 92259 2808
rect 92201 2799 92259 2805
rect 92934 2796 92940 2808
rect 92992 2796 92998 2848
rect 94961 2839 95019 2845
rect 94961 2805 94973 2839
rect 95007 2836 95019 2839
rect 95510 2836 95516 2848
rect 95007 2808 95516 2836
rect 95007 2805 95019 2808
rect 94961 2799 95019 2805
rect 95510 2796 95516 2808
rect 95568 2796 95574 2848
rect 97721 2839 97779 2845
rect 97721 2805 97733 2839
rect 97767 2836 97779 2839
rect 97902 2836 97908 2848
rect 97767 2808 97908 2836
rect 97767 2805 97779 2808
rect 97721 2799 97779 2805
rect 97902 2796 97908 2808
rect 97960 2796 97966 2848
rect 98454 2836 98460 2848
rect 98415 2808 98460 2836
rect 98454 2796 98460 2808
rect 98512 2796 98518 2848
rect 98638 2796 98644 2848
rect 98696 2836 98702 2848
rect 100481 2839 100539 2845
rect 100481 2836 100493 2839
rect 98696 2808 100493 2836
rect 98696 2796 98702 2808
rect 100481 2805 100493 2808
rect 100527 2836 100539 2839
rect 102318 2836 102324 2848
rect 100527 2808 102324 2836
rect 100527 2805 100539 2808
rect 100481 2799 100539 2805
rect 102318 2796 102324 2808
rect 102376 2796 102382 2848
rect 102962 2836 102968 2848
rect 102923 2808 102968 2836
rect 102962 2796 102968 2808
rect 103020 2796 103026 2848
rect 104805 2839 104863 2845
rect 104805 2805 104817 2839
rect 104851 2836 104863 2839
rect 105170 2836 105176 2848
rect 104851 2808 105176 2836
rect 104851 2805 104863 2808
rect 104805 2799 104863 2805
rect 105170 2796 105176 2808
rect 105228 2796 105234 2848
rect 105280 2836 105308 2876
rect 105633 2873 105645 2907
rect 105679 2904 105691 2907
rect 106844 2904 106872 3003
rect 107746 3000 107752 3052
rect 107804 3040 107810 3052
rect 107841 3043 107899 3049
rect 107841 3040 107853 3043
rect 107804 3012 107853 3040
rect 107804 3000 107810 3012
rect 107841 3009 107853 3012
rect 107887 3009 107899 3043
rect 108298 3040 108304 3052
rect 108259 3012 108304 3040
rect 107841 3003 107899 3009
rect 108298 3000 108304 3012
rect 108356 3000 108362 3052
rect 109034 3000 109040 3052
rect 109092 3040 109098 3052
rect 109788 3040 109816 3071
rect 109092 3012 109816 3040
rect 109865 3043 109923 3049
rect 109092 3000 109098 3012
rect 109865 3009 109877 3043
rect 109911 3040 109923 3043
rect 110506 3040 110512 3052
rect 109911 3012 110512 3040
rect 109911 3009 109923 3012
rect 109865 3003 109923 3009
rect 110506 3000 110512 3012
rect 110564 3000 110570 3052
rect 110601 3043 110659 3049
rect 110601 3009 110613 3043
rect 110647 3040 110659 3043
rect 110690 3040 110696 3052
rect 110647 3012 110696 3040
rect 110647 3009 110659 3012
rect 110601 3003 110659 3009
rect 110690 3000 110696 3012
rect 110748 3000 110754 3052
rect 111705 3043 111763 3049
rect 111705 3009 111717 3043
rect 111751 3009 111763 3043
rect 112530 3040 112536 3052
rect 112491 3012 112536 3040
rect 111705 3003 111763 3009
rect 109954 2932 109960 2984
rect 110012 2972 110018 2984
rect 110012 2944 110057 2972
rect 110012 2932 110018 2944
rect 109405 2907 109463 2913
rect 105679 2876 106872 2904
rect 106936 2876 109034 2904
rect 105679 2873 105691 2876
rect 105633 2867 105691 2873
rect 106936 2836 106964 2876
rect 107654 2836 107660 2848
rect 105280 2808 106964 2836
rect 107615 2808 107660 2836
rect 107654 2796 107660 2808
rect 107712 2796 107718 2848
rect 109006 2836 109034 2876
rect 109405 2873 109417 2907
rect 109451 2904 109463 2907
rect 111720 2904 111748 3003
rect 112530 3000 112536 3012
rect 112588 3000 112594 3052
rect 113450 3000 113456 3052
rect 113508 3040 113514 3052
rect 113729 3043 113787 3049
rect 113729 3040 113741 3043
rect 113508 3012 113741 3040
rect 113508 3000 113514 3012
rect 113729 3009 113741 3012
rect 113775 3009 113787 3043
rect 113729 3003 113787 3009
rect 115290 2972 115296 2984
rect 109451 2876 111748 2904
rect 111812 2944 115296 2972
rect 109451 2873 109463 2876
rect 109405 2867 109463 2873
rect 111812 2836 111840 2944
rect 115290 2932 115296 2944
rect 115348 2932 115354 2984
rect 115400 2904 115428 3080
rect 115492 3040 115520 3139
rect 116210 3136 116216 3148
rect 116268 3136 116274 3188
rect 116305 3179 116363 3185
rect 116305 3145 116317 3179
rect 116351 3176 116363 3179
rect 117041 3179 117099 3185
rect 117041 3176 117053 3179
rect 116351 3148 117053 3176
rect 116351 3145 116363 3148
rect 116305 3139 116363 3145
rect 117041 3145 117053 3148
rect 117087 3145 117099 3179
rect 117041 3139 117099 3145
rect 116857 3111 116915 3117
rect 116857 3108 116869 3111
rect 116228 3080 116869 3108
rect 116228 3049 116256 3080
rect 116857 3077 116869 3080
rect 116903 3077 116915 3111
rect 116857 3071 116915 3077
rect 116213 3043 116271 3049
rect 116213 3040 116225 3043
rect 115492 3012 116225 3040
rect 116213 3009 116225 3012
rect 116259 3009 116271 3043
rect 116213 3003 116271 3009
rect 116302 3000 116308 3052
rect 116360 3040 116366 3052
rect 117225 3043 117283 3049
rect 117225 3040 117237 3043
rect 116360 3012 117237 3040
rect 116360 3000 116366 3012
rect 117225 3009 117237 3012
rect 117271 3009 117283 3043
rect 117774 3040 117780 3052
rect 117735 3012 117780 3040
rect 117225 3003 117283 3009
rect 117774 3000 117780 3012
rect 117832 3000 117838 3052
rect 115474 2932 115480 2984
rect 115532 2972 115538 2984
rect 116394 2972 116400 2984
rect 115532 2944 116400 2972
rect 115532 2932 115538 2944
rect 116394 2932 116400 2944
rect 116452 2932 116458 2984
rect 117406 2904 117412 2916
rect 115400 2876 117412 2904
rect 117406 2864 117412 2876
rect 117464 2864 117470 2916
rect 112622 2836 112628 2848
rect 109006 2808 111840 2836
rect 112583 2808 112628 2836
rect 112622 2796 112628 2808
rect 112680 2796 112686 2848
rect 113542 2836 113548 2848
rect 113503 2808 113548 2836
rect 113542 2796 113548 2808
rect 113600 2796 113606 2848
rect 113634 2796 113640 2848
rect 113692 2836 113698 2848
rect 117869 2839 117927 2845
rect 117869 2836 117881 2839
rect 113692 2808 117881 2836
rect 113692 2796 113698 2808
rect 117869 2805 117881 2808
rect 117915 2805 117927 2839
rect 117869 2799 117927 2805
rect 1104 2746 118864 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 96374 2746
rect 96426 2694 96438 2746
rect 96490 2694 96502 2746
rect 96554 2694 96566 2746
rect 96618 2694 96630 2746
rect 96682 2694 118864 2746
rect 1104 2672 118864 2694
rect 5000 2604 55996 2632
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2397 1455 2431
rect 2130 2428 2136 2440
rect 2091 2400 2136 2428
rect 1397 2391 1455 2397
rect 1412 2360 1440 2391
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 5000 2437 5028 2604
rect 17034 2564 17040 2576
rect 16995 2536 17040 2564
rect 17034 2524 17040 2536
rect 17092 2524 17098 2576
rect 22557 2567 22615 2573
rect 21376 2536 22048 2564
rect 21376 2496 21404 2536
rect 5092 2468 21404 2496
rect 22020 2496 22048 2536
rect 22557 2533 22569 2567
rect 22603 2564 22615 2567
rect 55858 2564 55864 2576
rect 22603 2536 55864 2564
rect 22603 2533 22615 2536
rect 22557 2527 22615 2533
rect 55858 2524 55864 2536
rect 55916 2524 55922 2576
rect 35894 2496 35900 2508
rect 22020 2468 35900 2496
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 5092 2360 5120 2468
rect 35894 2456 35900 2468
rect 35952 2456 35958 2508
rect 35986 2456 35992 2508
rect 36044 2496 36050 2508
rect 45370 2496 45376 2508
rect 36044 2468 45376 2496
rect 36044 2456 36050 2468
rect 45370 2456 45376 2468
rect 45428 2456 45434 2508
rect 45462 2456 45468 2508
rect 45520 2496 45526 2508
rect 55766 2496 55772 2508
rect 45520 2468 55772 2496
rect 45520 2456 45526 2468
rect 55766 2456 55772 2468
rect 55824 2456 55830 2508
rect 55968 2496 55996 2604
rect 56134 2592 56140 2644
rect 56192 2632 56198 2644
rect 56781 2635 56839 2641
rect 56781 2632 56793 2635
rect 56192 2604 56793 2632
rect 56192 2592 56198 2604
rect 56781 2601 56793 2604
rect 56827 2632 56839 2635
rect 57146 2632 57152 2644
rect 56827 2604 57152 2632
rect 56827 2601 56839 2604
rect 56781 2595 56839 2601
rect 57146 2592 57152 2604
rect 57204 2592 57210 2644
rect 58250 2632 58256 2644
rect 58211 2604 58256 2632
rect 58250 2592 58256 2604
rect 58308 2592 58314 2644
rect 58434 2592 58440 2644
rect 58492 2632 58498 2644
rect 59633 2635 59691 2641
rect 59633 2632 59645 2635
rect 58492 2604 59645 2632
rect 58492 2592 58498 2604
rect 59633 2601 59645 2604
rect 59679 2601 59691 2635
rect 64138 2632 64144 2644
rect 59633 2595 59691 2601
rect 60292 2604 60504 2632
rect 64099 2604 64144 2632
rect 56042 2524 56048 2576
rect 56100 2564 56106 2576
rect 60292 2564 60320 2604
rect 56100 2536 60320 2564
rect 60476 2564 60504 2604
rect 64138 2592 64144 2604
rect 64196 2592 64202 2644
rect 64693 2635 64751 2641
rect 64693 2601 64705 2635
rect 64739 2632 64751 2635
rect 64874 2632 64880 2644
rect 64739 2604 64880 2632
rect 64739 2601 64751 2604
rect 64693 2595 64751 2601
rect 64874 2592 64880 2604
rect 64932 2592 64938 2644
rect 65150 2632 65156 2644
rect 65111 2604 65156 2632
rect 65150 2592 65156 2604
rect 65208 2592 65214 2644
rect 65242 2592 65248 2644
rect 65300 2632 65306 2644
rect 74626 2632 74632 2644
rect 65300 2604 74534 2632
rect 74587 2604 74632 2632
rect 65300 2592 65306 2604
rect 74506 2564 74534 2604
rect 74626 2592 74632 2604
rect 74684 2592 74690 2644
rect 75917 2635 75975 2641
rect 75917 2601 75929 2635
rect 75963 2632 75975 2635
rect 76558 2632 76564 2644
rect 75963 2604 76564 2632
rect 75963 2601 75975 2604
rect 75917 2595 75975 2601
rect 76558 2592 76564 2604
rect 76616 2592 76622 2644
rect 77205 2635 77263 2641
rect 77205 2601 77217 2635
rect 77251 2632 77263 2635
rect 78582 2632 78588 2644
rect 77251 2604 78588 2632
rect 77251 2601 77263 2604
rect 77205 2595 77263 2601
rect 78582 2592 78588 2604
rect 78640 2592 78646 2644
rect 78677 2635 78735 2641
rect 78677 2601 78689 2635
rect 78723 2632 78735 2635
rect 79502 2632 79508 2644
rect 78723 2604 79508 2632
rect 78723 2601 78735 2604
rect 78677 2595 78735 2601
rect 79502 2592 79508 2604
rect 79560 2592 79566 2644
rect 79594 2592 79600 2644
rect 79652 2632 79658 2644
rect 80882 2632 80888 2644
rect 79652 2604 80888 2632
rect 79652 2592 79658 2604
rect 80882 2592 80888 2604
rect 80940 2592 80946 2644
rect 81069 2635 81127 2641
rect 81069 2601 81081 2635
rect 81115 2632 81127 2635
rect 81618 2632 81624 2644
rect 81115 2604 81624 2632
rect 81115 2601 81127 2604
rect 81069 2595 81127 2601
rect 81618 2592 81624 2604
rect 81676 2592 81682 2644
rect 82538 2592 82544 2644
rect 82596 2632 82602 2644
rect 82633 2635 82691 2641
rect 82633 2632 82645 2635
rect 82596 2604 82645 2632
rect 82596 2592 82602 2604
rect 82633 2601 82645 2604
rect 82679 2601 82691 2635
rect 82633 2595 82691 2601
rect 83645 2635 83703 2641
rect 83645 2601 83657 2635
rect 83691 2632 83703 2635
rect 83734 2632 83740 2644
rect 83691 2604 83740 2632
rect 83691 2601 83703 2604
rect 83645 2595 83703 2601
rect 83734 2592 83740 2604
rect 83792 2592 83798 2644
rect 84841 2635 84899 2641
rect 84841 2601 84853 2635
rect 84887 2632 84899 2635
rect 85114 2632 85120 2644
rect 84887 2604 85120 2632
rect 84887 2601 84899 2604
rect 84841 2595 84899 2601
rect 85114 2592 85120 2604
rect 85172 2592 85178 2644
rect 86221 2635 86279 2641
rect 86221 2601 86233 2635
rect 86267 2632 86279 2635
rect 86586 2632 86592 2644
rect 86267 2604 86592 2632
rect 86267 2601 86279 2604
rect 86221 2595 86279 2601
rect 86586 2592 86592 2604
rect 86644 2592 86650 2644
rect 87509 2635 87567 2641
rect 87509 2601 87521 2635
rect 87555 2632 87567 2635
rect 88334 2632 88340 2644
rect 87555 2604 88340 2632
rect 87555 2601 87567 2604
rect 87509 2595 87567 2601
rect 88334 2592 88340 2604
rect 88392 2592 88398 2644
rect 88794 2632 88800 2644
rect 88755 2604 88800 2632
rect 88794 2592 88800 2604
rect 88852 2592 88858 2644
rect 90085 2635 90143 2641
rect 90085 2601 90097 2635
rect 90131 2632 90143 2635
rect 90818 2632 90824 2644
rect 90131 2604 90824 2632
rect 90131 2601 90143 2604
rect 90085 2595 90143 2601
rect 90818 2592 90824 2604
rect 90876 2592 90882 2644
rect 91557 2635 91615 2641
rect 91557 2601 91569 2635
rect 91603 2632 91615 2635
rect 92198 2632 92204 2644
rect 91603 2604 92204 2632
rect 91603 2601 91615 2604
rect 91557 2595 91615 2601
rect 92198 2592 92204 2604
rect 92256 2592 92262 2644
rect 93118 2632 93124 2644
rect 93079 2604 93124 2632
rect 93118 2592 93124 2604
rect 93176 2592 93182 2644
rect 93946 2592 93952 2644
rect 94004 2632 94010 2644
rect 95053 2635 95111 2641
rect 94004 2604 94049 2632
rect 94004 2592 94010 2604
rect 95053 2601 95065 2635
rect 95099 2632 95111 2635
rect 95786 2632 95792 2644
rect 95099 2604 95792 2632
rect 95099 2601 95111 2604
rect 95053 2595 95111 2601
rect 95786 2592 95792 2604
rect 95844 2592 95850 2644
rect 96246 2592 96252 2644
rect 96304 2632 96310 2644
rect 96525 2635 96583 2641
rect 96525 2632 96537 2635
rect 96304 2604 96537 2632
rect 96304 2592 96310 2604
rect 96525 2601 96537 2604
rect 96571 2601 96583 2635
rect 96525 2595 96583 2601
rect 97902 2592 97908 2644
rect 97960 2632 97966 2644
rect 100294 2632 100300 2644
rect 97960 2604 99788 2632
rect 100255 2604 100300 2632
rect 97960 2592 97966 2604
rect 97534 2564 97540 2576
rect 60476 2536 73752 2564
rect 74506 2536 97540 2564
rect 56100 2524 56106 2536
rect 60274 2496 60280 2508
rect 55968 2468 60280 2496
rect 60274 2456 60280 2468
rect 60332 2456 60338 2508
rect 60642 2456 60648 2508
rect 60700 2496 60706 2508
rect 60826 2496 60832 2508
rect 60700 2468 60832 2496
rect 60700 2456 60706 2468
rect 60826 2456 60832 2468
rect 60884 2456 60890 2508
rect 61286 2456 61292 2508
rect 61344 2496 61350 2508
rect 73724 2496 73752 2536
rect 97534 2524 97540 2536
rect 97592 2524 97598 2576
rect 97718 2564 97724 2576
rect 97679 2536 97724 2564
rect 97718 2524 97724 2536
rect 97776 2524 97782 2576
rect 74810 2496 74816 2508
rect 61344 2468 73660 2496
rect 73724 2468 74816 2496
rect 61344 2456 61350 2468
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 7561 2431 7619 2437
rect 6503 2400 6914 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 1412 2332 5120 2360
rect 658 2252 664 2304
rect 716 2292 722 2304
rect 1581 2295 1639 2301
rect 1581 2292 1593 2295
rect 716 2264 1593 2292
rect 716 2252 722 2264
rect 1581 2261 1593 2264
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 2038 2252 2044 2304
rect 2096 2292 2102 2304
rect 2317 2295 2375 2301
rect 2317 2292 2329 2295
rect 2096 2264 2329 2292
rect 2096 2252 2102 2264
rect 2317 2261 2329 2264
rect 2363 2261 2375 2295
rect 2317 2255 2375 2261
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3568 2264 3985 2292
rect 3568 2252 3574 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 4890 2252 4896 2304
rect 4948 2292 4954 2304
rect 5169 2295 5227 2301
rect 5169 2292 5181 2295
rect 4948 2264 5181 2292
rect 4948 2252 4954 2264
rect 5169 2261 5181 2264
rect 5215 2261 5227 2295
rect 5169 2255 5227 2261
rect 6362 2252 6368 2304
rect 6420 2292 6426 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6420 2264 6653 2292
rect 6420 2252 6426 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6886 2292 6914 2400
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 7834 2428 7840 2440
rect 7607 2400 7840 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10686 2428 10692 2440
rect 10459 2400 10692 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 9324 2360 9352 2391
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 12158 2428 12164 2440
rect 12119 2400 12164 2428
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22281 2431 22339 2437
rect 22281 2428 22293 2431
rect 22060 2400 22293 2428
rect 22060 2388 22066 2400
rect 22281 2397 22293 2400
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 22388 2400 25544 2428
rect 9953 2363 10011 2369
rect 9953 2360 9965 2363
rect 9324 2332 9965 2360
rect 9953 2329 9965 2332
rect 9999 2360 10011 2363
rect 9999 2332 14412 2360
rect 9999 2329 10011 2332
rect 9953 2323 10011 2329
rect 7098 2292 7104 2304
rect 6886 2264 7104 2292
rect 6641 2255 6699 2261
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7800 2264 8033 2292
rect 7800 2252 7806 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 9493 2295 9551 2301
rect 9493 2292 9505 2295
rect 9272 2264 9505 2292
rect 9272 2252 9278 2264
rect 9493 2261 9505 2264
rect 9539 2261 9551 2295
rect 9493 2255 9551 2261
rect 10594 2252 10600 2304
rect 10652 2292 10658 2304
rect 10873 2295 10931 2301
rect 10873 2292 10885 2295
rect 10652 2264 10885 2292
rect 10652 2252 10658 2264
rect 10873 2261 10885 2264
rect 10919 2261 10931 2295
rect 10873 2255 10931 2261
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12345 2295 12403 2301
rect 12345 2292 12357 2295
rect 12124 2264 12357 2292
rect 12124 2252 12130 2264
rect 12345 2261 12357 2264
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 13446 2252 13452 2304
rect 13504 2292 13510 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13504 2264 14289 2292
rect 13504 2252 13510 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14384 2292 14412 2332
rect 14918 2320 14924 2372
rect 14976 2360 14982 2372
rect 15105 2363 15163 2369
rect 15105 2360 15117 2363
rect 14976 2332 15117 2360
rect 14976 2320 14982 2332
rect 15105 2329 15117 2332
rect 15151 2329 15163 2363
rect 15470 2360 15476 2372
rect 15431 2332 15476 2360
rect 15105 2323 15163 2329
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 16298 2320 16304 2372
rect 16356 2360 16362 2372
rect 16761 2363 16819 2369
rect 16761 2360 16773 2363
rect 16356 2332 16773 2360
rect 16356 2320 16362 2332
rect 16761 2329 16773 2332
rect 16807 2329 16819 2363
rect 16761 2323 16819 2329
rect 17770 2320 17776 2372
rect 17828 2360 17834 2372
rect 17957 2363 18015 2369
rect 17957 2360 17969 2363
rect 17828 2332 17969 2360
rect 17828 2320 17834 2332
rect 17957 2329 17969 2332
rect 18003 2329 18015 2363
rect 18322 2360 18328 2372
rect 18283 2332 18328 2360
rect 17957 2323 18015 2329
rect 18322 2320 18328 2332
rect 18380 2320 18386 2372
rect 19150 2320 19156 2372
rect 19208 2360 19214 2372
rect 19337 2363 19395 2369
rect 19337 2360 19349 2363
rect 19208 2332 19349 2360
rect 19208 2320 19214 2332
rect 19337 2329 19349 2332
rect 19383 2329 19395 2363
rect 19337 2323 19395 2329
rect 20622 2320 20628 2372
rect 20680 2360 20686 2372
rect 20809 2363 20867 2369
rect 20809 2360 20821 2363
rect 20680 2332 20821 2360
rect 20680 2320 20686 2332
rect 20809 2329 20821 2332
rect 20855 2329 20867 2363
rect 20809 2323 20867 2329
rect 22097 2363 22155 2369
rect 22097 2329 22109 2363
rect 22143 2360 22155 2363
rect 22388 2360 22416 2400
rect 22143 2332 22416 2360
rect 22143 2329 22155 2332
rect 22097 2323 22155 2329
rect 19426 2292 19432 2304
rect 14384 2264 19432 2292
rect 14277 2255 14335 2261
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 19613 2295 19671 2301
rect 19613 2261 19625 2295
rect 19659 2292 19671 2295
rect 19978 2292 19984 2304
rect 19659 2264 19984 2292
rect 19659 2261 19671 2264
rect 19613 2255 19671 2261
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 20073 2295 20131 2301
rect 20073 2261 20085 2295
rect 20119 2292 20131 2295
rect 20441 2295 20499 2301
rect 20441 2292 20453 2295
rect 20119 2264 20453 2292
rect 20119 2261 20131 2264
rect 20073 2255 20131 2261
rect 20441 2261 20453 2264
rect 20487 2292 20499 2295
rect 21085 2295 21143 2301
rect 21085 2292 21097 2295
rect 20487 2264 21097 2292
rect 20487 2261 20499 2264
rect 20441 2255 20499 2261
rect 21085 2261 21097 2264
rect 21131 2292 21143 2295
rect 22112 2292 22140 2323
rect 23474 2320 23480 2372
rect 23532 2360 23538 2372
rect 24489 2363 24547 2369
rect 24489 2360 24501 2363
rect 23532 2332 24501 2360
rect 23532 2320 23538 2332
rect 24489 2329 24501 2332
rect 24535 2329 24547 2363
rect 24489 2323 24547 2329
rect 24946 2320 24952 2372
rect 25004 2360 25010 2372
rect 25409 2363 25467 2369
rect 25409 2360 25421 2363
rect 25004 2332 25421 2360
rect 25004 2320 25010 2332
rect 25409 2329 25421 2332
rect 25455 2329 25467 2363
rect 25516 2360 25544 2400
rect 25774 2388 25780 2440
rect 25832 2428 25838 2440
rect 35710 2428 35716 2440
rect 25832 2400 35716 2428
rect 25832 2388 25838 2400
rect 35710 2388 35716 2400
rect 35768 2388 35774 2440
rect 35802 2388 35808 2440
rect 35860 2428 35866 2440
rect 35860 2400 59676 2428
rect 35860 2388 35866 2400
rect 26234 2360 26240 2372
rect 25516 2332 26240 2360
rect 25409 2323 25467 2329
rect 26234 2320 26240 2332
rect 26292 2320 26298 2372
rect 26326 2320 26332 2372
rect 26384 2360 26390 2372
rect 27065 2363 27123 2369
rect 27065 2360 27077 2363
rect 26384 2332 27077 2360
rect 26384 2320 26390 2332
rect 27065 2329 27077 2332
rect 27111 2329 27123 2363
rect 27065 2323 27123 2329
rect 27706 2320 27712 2372
rect 27764 2360 27770 2372
rect 27985 2363 28043 2369
rect 27985 2360 27997 2363
rect 27764 2332 27997 2360
rect 27764 2320 27770 2332
rect 27985 2329 27997 2332
rect 28031 2329 28043 2363
rect 27985 2323 28043 2329
rect 29178 2320 29184 2372
rect 29236 2360 29242 2372
rect 29641 2363 29699 2369
rect 29641 2360 29653 2363
rect 29236 2332 29653 2360
rect 29236 2320 29242 2332
rect 29641 2329 29653 2332
rect 29687 2329 29699 2363
rect 30006 2360 30012 2372
rect 29967 2332 30012 2360
rect 29641 2323 29699 2329
rect 30006 2320 30012 2332
rect 30064 2320 30070 2372
rect 30834 2320 30840 2372
rect 30892 2360 30898 2372
rect 30892 2332 30937 2360
rect 31036 2332 31984 2360
rect 30892 2320 30898 2332
rect 24762 2292 24768 2304
rect 21131 2264 22140 2292
rect 24723 2264 24768 2292
rect 21131 2261 21143 2264
rect 21085 2255 21143 2261
rect 24762 2252 24768 2264
rect 24820 2252 24826 2304
rect 25682 2252 25688 2304
rect 25740 2292 25746 2304
rect 27338 2292 27344 2304
rect 25740 2264 25785 2292
rect 27299 2264 27344 2292
rect 25740 2252 25746 2264
rect 27338 2252 27344 2264
rect 27396 2252 27402 2304
rect 28261 2295 28319 2301
rect 28261 2261 28273 2295
rect 28307 2292 28319 2295
rect 31036 2292 31064 2332
rect 28307 2264 31064 2292
rect 31113 2295 31171 2301
rect 28307 2261 28319 2264
rect 28261 2255 28319 2261
rect 31113 2261 31125 2295
rect 31159 2292 31171 2295
rect 31662 2292 31668 2304
rect 31159 2264 31668 2292
rect 31159 2261 31171 2264
rect 31113 2255 31171 2261
rect 31662 2252 31668 2264
rect 31720 2252 31726 2304
rect 31956 2292 31984 2332
rect 32030 2320 32036 2372
rect 32088 2360 32094 2372
rect 32217 2363 32275 2369
rect 32217 2360 32229 2363
rect 32088 2332 32229 2360
rect 32088 2320 32094 2332
rect 32217 2329 32229 2332
rect 32263 2329 32275 2363
rect 32582 2360 32588 2372
rect 32543 2332 32588 2360
rect 32217 2323 32275 2329
rect 32582 2320 32588 2332
rect 32640 2320 32646 2372
rect 33410 2360 33416 2372
rect 32876 2332 33416 2360
rect 32876 2292 32904 2332
rect 33410 2320 33416 2332
rect 33468 2320 33474 2372
rect 33502 2320 33508 2372
rect 33560 2360 33566 2372
rect 33689 2363 33747 2369
rect 33689 2360 33701 2363
rect 33560 2332 33701 2360
rect 33560 2320 33566 2332
rect 33689 2329 33701 2332
rect 33735 2329 33747 2363
rect 33689 2323 33747 2329
rect 35158 2320 35164 2372
rect 35216 2360 35222 2372
rect 37274 2360 37280 2372
rect 35216 2332 35261 2360
rect 35360 2332 37280 2360
rect 35216 2320 35222 2332
rect 31956 2264 32904 2292
rect 32953 2295 33011 2301
rect 32953 2261 32965 2295
rect 32999 2292 33011 2295
rect 33321 2295 33379 2301
rect 33321 2292 33333 2295
rect 32999 2264 33333 2292
rect 32999 2261 33011 2264
rect 32953 2255 33011 2261
rect 33321 2261 33333 2264
rect 33367 2292 33379 2295
rect 33965 2295 34023 2301
rect 33965 2292 33977 2295
rect 33367 2264 33977 2292
rect 33367 2261 33379 2264
rect 33321 2255 33379 2261
rect 33965 2261 33977 2264
rect 34011 2292 34023 2295
rect 34977 2295 35035 2301
rect 34977 2292 34989 2295
rect 34011 2264 34989 2292
rect 34011 2261 34023 2264
rect 33965 2255 34023 2261
rect 34977 2261 34989 2264
rect 35023 2292 35035 2295
rect 35360 2292 35388 2332
rect 37274 2320 37280 2332
rect 37332 2320 37338 2372
rect 37369 2363 37427 2369
rect 37369 2329 37381 2363
rect 37415 2329 37427 2363
rect 37369 2323 37427 2329
rect 35023 2264 35388 2292
rect 35437 2295 35495 2301
rect 35023 2261 35035 2264
rect 34977 2255 35035 2261
rect 35437 2261 35449 2295
rect 35483 2292 35495 2295
rect 35526 2292 35532 2304
rect 35483 2264 35532 2292
rect 35483 2261 35495 2264
rect 35437 2255 35495 2261
rect 35526 2252 35532 2264
rect 35584 2252 35590 2304
rect 36354 2252 36360 2304
rect 36412 2292 36418 2304
rect 37384 2292 37412 2323
rect 37734 2320 37740 2372
rect 37792 2360 37798 2372
rect 38289 2363 38347 2369
rect 38289 2360 38301 2363
rect 37792 2332 38301 2360
rect 37792 2320 37798 2332
rect 38289 2329 38301 2332
rect 38335 2329 38347 2363
rect 38289 2323 38347 2329
rect 39206 2320 39212 2372
rect 39264 2360 39270 2372
rect 39945 2363 40003 2369
rect 39945 2360 39957 2363
rect 39264 2332 39957 2360
rect 39264 2320 39270 2332
rect 39945 2329 39957 2332
rect 39991 2329 40003 2363
rect 39945 2323 40003 2329
rect 40586 2320 40592 2372
rect 40644 2360 40650 2372
rect 40865 2363 40923 2369
rect 40865 2360 40877 2363
rect 40644 2332 40877 2360
rect 40644 2320 40650 2332
rect 40865 2329 40877 2332
rect 40911 2329 40923 2363
rect 40865 2323 40923 2329
rect 42058 2320 42064 2372
rect 42116 2360 42122 2372
rect 42521 2363 42579 2369
rect 42521 2360 42533 2363
rect 42116 2332 42533 2360
rect 42116 2320 42122 2332
rect 42521 2329 42533 2332
rect 42567 2329 42579 2363
rect 42521 2323 42579 2329
rect 43438 2320 43444 2372
rect 43496 2360 43502 2372
rect 43625 2363 43683 2369
rect 43625 2360 43637 2363
rect 43496 2332 43637 2360
rect 43496 2320 43502 2332
rect 43625 2329 43637 2332
rect 43671 2329 43683 2363
rect 43625 2323 43683 2329
rect 44910 2320 44916 2372
rect 44968 2360 44974 2372
rect 45097 2363 45155 2369
rect 45097 2360 45109 2363
rect 44968 2332 45109 2360
rect 44968 2320 44974 2332
rect 45097 2329 45109 2332
rect 45143 2329 45155 2363
rect 45097 2323 45155 2329
rect 46290 2320 46296 2372
rect 46348 2360 46354 2372
rect 46477 2363 46535 2369
rect 46477 2360 46489 2363
rect 46348 2332 46489 2360
rect 46348 2320 46354 2332
rect 46477 2329 46489 2332
rect 46523 2329 46535 2363
rect 46477 2323 46535 2329
rect 46845 2363 46903 2369
rect 46845 2329 46857 2363
rect 46891 2360 46903 2363
rect 47670 2360 47676 2372
rect 46891 2332 47676 2360
rect 46891 2329 46903 2332
rect 46845 2323 46903 2329
rect 47670 2320 47676 2332
rect 47728 2320 47734 2372
rect 47762 2320 47768 2372
rect 47820 2360 47826 2372
rect 47949 2363 48007 2369
rect 47949 2360 47961 2363
rect 47820 2332 47961 2360
rect 47820 2320 47826 2332
rect 47949 2329 47961 2332
rect 47995 2329 48007 2363
rect 49050 2360 49056 2372
rect 47949 2323 48007 2329
rect 48148 2332 49056 2360
rect 37642 2292 37648 2304
rect 36412 2264 37412 2292
rect 37603 2264 37648 2292
rect 36412 2252 36418 2264
rect 37642 2252 37648 2264
rect 37700 2252 37706 2304
rect 38562 2292 38568 2304
rect 38523 2264 38568 2292
rect 38562 2252 38568 2264
rect 38620 2252 38626 2304
rect 40221 2295 40279 2301
rect 40221 2261 40233 2295
rect 40267 2292 40279 2295
rect 40494 2292 40500 2304
rect 40267 2264 40500 2292
rect 40267 2261 40279 2264
rect 40221 2255 40279 2261
rect 40494 2252 40500 2264
rect 40552 2252 40558 2304
rect 41138 2292 41144 2304
rect 41099 2264 41144 2292
rect 41138 2252 41144 2264
rect 41196 2252 41202 2304
rect 42794 2292 42800 2304
rect 42755 2264 42800 2292
rect 42794 2252 42800 2264
rect 42852 2252 42858 2304
rect 43898 2292 43904 2304
rect 43859 2264 43904 2292
rect 43898 2252 43904 2264
rect 43956 2252 43962 2304
rect 45186 2252 45192 2304
rect 45244 2292 45250 2304
rect 45244 2264 45289 2292
rect 45244 2252 45250 2264
rect 45370 2252 45376 2304
rect 45428 2292 45434 2304
rect 48148 2292 48176 2332
rect 49050 2320 49056 2332
rect 49108 2320 49114 2372
rect 49142 2320 49148 2372
rect 49200 2360 49206 2372
rect 49237 2363 49295 2369
rect 49237 2360 49249 2363
rect 49200 2332 49249 2360
rect 49200 2320 49206 2332
rect 49237 2329 49249 2332
rect 49283 2329 49295 2363
rect 49237 2323 49295 2329
rect 49436 2332 50568 2360
rect 45428 2264 48176 2292
rect 48225 2295 48283 2301
rect 45428 2252 45434 2264
rect 48225 2261 48237 2295
rect 48271 2292 48283 2295
rect 49436 2292 49464 2332
rect 48271 2264 49464 2292
rect 49513 2295 49571 2301
rect 48271 2261 48283 2264
rect 48225 2255 48283 2261
rect 49513 2261 49525 2295
rect 49559 2292 49571 2295
rect 49602 2292 49608 2304
rect 49559 2264 49608 2292
rect 49559 2261 49571 2264
rect 49513 2255 49571 2261
rect 49602 2252 49608 2264
rect 49660 2252 49666 2304
rect 50540 2292 50568 2332
rect 50614 2320 50620 2372
rect 50672 2360 50678 2372
rect 50801 2363 50859 2369
rect 50801 2360 50813 2363
rect 50672 2332 50813 2360
rect 50672 2320 50678 2332
rect 50801 2329 50813 2332
rect 50847 2329 50859 2363
rect 50801 2323 50859 2329
rect 51169 2363 51227 2369
rect 51169 2329 51181 2363
rect 51215 2360 51227 2363
rect 51902 2360 51908 2372
rect 51215 2332 51908 2360
rect 51215 2329 51227 2332
rect 51169 2323 51227 2329
rect 51902 2320 51908 2332
rect 51960 2320 51966 2372
rect 51994 2320 52000 2372
rect 52052 2360 52058 2372
rect 52825 2363 52883 2369
rect 52825 2360 52837 2363
rect 52052 2332 52837 2360
rect 52052 2320 52058 2332
rect 52825 2329 52837 2332
rect 52871 2329 52883 2363
rect 53374 2360 53380 2372
rect 52825 2323 52883 2329
rect 53024 2332 53380 2360
rect 53024 2292 53052 2332
rect 53374 2320 53380 2332
rect 53432 2320 53438 2372
rect 53466 2320 53472 2372
rect 53524 2360 53530 2372
rect 53745 2363 53803 2369
rect 53745 2360 53757 2363
rect 53524 2332 53757 2360
rect 53524 2320 53530 2332
rect 53745 2329 53757 2332
rect 53791 2329 53803 2363
rect 53745 2323 53803 2329
rect 54113 2363 54171 2369
rect 54113 2329 54125 2363
rect 54159 2360 54171 2363
rect 56505 2363 56563 2369
rect 54159 2332 56364 2360
rect 54159 2329 54171 2332
rect 54113 2323 54171 2329
rect 50540 2264 53052 2292
rect 53101 2295 53159 2301
rect 53101 2261 53113 2295
rect 53147 2292 53159 2295
rect 55674 2292 55680 2304
rect 53147 2264 55680 2292
rect 53147 2261 53159 2264
rect 53101 2255 53159 2261
rect 55674 2252 55680 2264
rect 55732 2252 55738 2304
rect 55769 2295 55827 2301
rect 55769 2261 55781 2295
rect 55815 2292 55827 2295
rect 56134 2292 56140 2304
rect 55815 2264 56140 2292
rect 55815 2261 55827 2264
rect 55769 2255 55827 2261
rect 56134 2252 56140 2264
rect 56192 2252 56198 2304
rect 56336 2292 56364 2332
rect 56505 2329 56517 2363
rect 56551 2360 56563 2363
rect 56686 2360 56692 2372
rect 56551 2332 56692 2360
rect 56551 2329 56563 2332
rect 56505 2323 56563 2329
rect 56686 2320 56692 2332
rect 56744 2320 56750 2372
rect 57698 2320 57704 2372
rect 57756 2360 57762 2372
rect 57977 2363 58035 2369
rect 57977 2360 57989 2363
rect 57756 2332 57989 2360
rect 57756 2320 57762 2332
rect 57977 2329 57989 2332
rect 58023 2329 58035 2363
rect 59538 2360 59544 2372
rect 59499 2332 59544 2360
rect 57977 2323 58035 2329
rect 59538 2320 59544 2332
rect 59596 2320 59602 2372
rect 59648 2360 59676 2400
rect 59906 2388 59912 2440
rect 59964 2428 59970 2440
rect 61381 2431 61439 2437
rect 61381 2428 61393 2431
rect 59964 2424 60412 2428
rect 60476 2424 61393 2428
rect 59964 2400 61393 2424
rect 59964 2388 59970 2400
rect 60384 2396 60504 2400
rect 61381 2397 61393 2400
rect 61427 2397 61439 2431
rect 61381 2391 61439 2397
rect 62114 2388 62120 2440
rect 62172 2428 62178 2440
rect 62172 2400 62217 2428
rect 62172 2388 62178 2400
rect 63402 2388 63408 2440
rect 63460 2428 63466 2440
rect 63497 2431 63555 2437
rect 63497 2428 63509 2431
rect 63460 2400 63509 2428
rect 63460 2388 63466 2400
rect 63497 2397 63509 2400
rect 63543 2397 63555 2431
rect 63497 2391 63555 2397
rect 64049 2431 64107 2437
rect 64049 2397 64061 2431
rect 64095 2428 64107 2431
rect 64414 2428 64420 2440
rect 64095 2400 64420 2428
rect 64095 2397 64107 2400
rect 64049 2391 64107 2397
rect 64414 2388 64420 2400
rect 64472 2428 64478 2440
rect 64877 2431 64935 2437
rect 64877 2428 64889 2431
rect 64472 2400 64889 2428
rect 64472 2388 64478 2400
rect 64877 2397 64889 2400
rect 64923 2397 64935 2431
rect 64877 2391 64935 2397
rect 65518 2388 65524 2440
rect 65576 2428 65582 2440
rect 65705 2431 65763 2437
rect 65705 2428 65717 2431
rect 65576 2400 65717 2428
rect 65576 2388 65582 2400
rect 65705 2397 65717 2400
rect 65751 2397 65763 2431
rect 66714 2428 66720 2440
rect 66675 2400 66720 2428
rect 65705 2391 65763 2397
rect 66714 2388 66720 2400
rect 66772 2388 66778 2440
rect 68278 2428 68284 2440
rect 68239 2400 68284 2428
rect 68278 2388 68284 2400
rect 68336 2388 68342 2440
rect 69566 2428 69572 2440
rect 69527 2400 69572 2428
rect 69566 2388 69572 2400
rect 69624 2388 69630 2440
rect 69658 2388 69664 2440
rect 69716 2428 69722 2440
rect 72786 2428 72792 2440
rect 69716 2400 72556 2428
rect 72747 2400 72792 2428
rect 69716 2388 69722 2400
rect 60182 2360 60188 2372
rect 59648 2332 60188 2360
rect 60182 2320 60188 2332
rect 60240 2320 60246 2372
rect 61010 2320 61016 2372
rect 61068 2360 61074 2372
rect 61068 2332 61113 2360
rect 61068 2320 61074 2332
rect 63126 2320 63132 2372
rect 63184 2360 63190 2372
rect 63184 2332 63229 2360
rect 63184 2320 63190 2332
rect 63310 2320 63316 2372
rect 63368 2360 63374 2372
rect 63368 2332 69704 2360
rect 63368 2320 63374 2332
rect 59630 2292 59636 2304
rect 56336 2264 59636 2292
rect 59630 2252 59636 2264
rect 59688 2252 59694 2304
rect 59722 2252 59728 2304
rect 59780 2292 59786 2304
rect 61930 2292 61936 2304
rect 59780 2264 61936 2292
rect 59780 2252 59786 2264
rect 61930 2252 61936 2264
rect 61988 2252 61994 2304
rect 62022 2252 62028 2304
rect 62080 2292 62086 2304
rect 62301 2295 62359 2301
rect 62301 2292 62313 2295
rect 62080 2264 62313 2292
rect 62080 2252 62086 2264
rect 62301 2261 62313 2264
rect 62347 2261 62359 2295
rect 62301 2255 62359 2261
rect 65150 2252 65156 2304
rect 65208 2292 65214 2304
rect 65797 2295 65855 2301
rect 65797 2292 65809 2295
rect 65208 2264 65809 2292
rect 65208 2252 65214 2264
rect 65797 2261 65809 2264
rect 65843 2261 65855 2295
rect 66806 2292 66812 2304
rect 66767 2264 66812 2292
rect 65797 2255 65855 2261
rect 66806 2252 66812 2264
rect 66864 2292 66870 2304
rect 67361 2295 67419 2301
rect 67361 2292 67373 2295
rect 66864 2264 67373 2292
rect 66864 2252 66870 2264
rect 67361 2261 67373 2264
rect 67407 2261 67419 2295
rect 67361 2255 67419 2261
rect 67450 2252 67456 2304
rect 67508 2292 67514 2304
rect 69676 2301 69704 2332
rect 69750 2320 69756 2372
rect 69808 2360 69814 2372
rect 71041 2363 71099 2369
rect 69808 2332 70394 2360
rect 69808 2320 69814 2332
rect 68373 2295 68431 2301
rect 68373 2292 68385 2295
rect 67508 2264 68385 2292
rect 67508 2252 67514 2264
rect 68373 2261 68385 2264
rect 68419 2292 68431 2295
rect 68925 2295 68983 2301
rect 68925 2292 68937 2295
rect 68419 2264 68937 2292
rect 68419 2261 68431 2264
rect 68373 2255 68431 2261
rect 68925 2261 68937 2264
rect 68971 2261 68983 2295
rect 68925 2255 68983 2261
rect 69661 2295 69719 2301
rect 69661 2261 69673 2295
rect 69707 2292 69719 2295
rect 70213 2295 70271 2301
rect 70213 2292 70225 2295
rect 69707 2264 70225 2292
rect 69707 2261 69719 2264
rect 69661 2255 69719 2261
rect 70213 2261 70225 2264
rect 70259 2261 70271 2295
rect 70366 2292 70394 2332
rect 71041 2329 71053 2363
rect 71087 2360 71099 2363
rect 71682 2360 71688 2372
rect 71087 2332 71688 2360
rect 71087 2329 71099 2332
rect 71041 2323 71099 2329
rect 71682 2320 71688 2332
rect 71740 2320 71746 2372
rect 72421 2363 72479 2369
rect 72421 2329 72433 2363
rect 72467 2329 72479 2363
rect 72528 2360 72556 2400
rect 72786 2388 72792 2400
rect 72844 2388 72850 2440
rect 73522 2428 73528 2440
rect 73483 2400 73528 2428
rect 73522 2388 73528 2400
rect 73580 2388 73586 2440
rect 73632 2428 73660 2468
rect 74810 2456 74816 2468
rect 74868 2456 74874 2508
rect 74994 2456 75000 2508
rect 75052 2496 75058 2508
rect 75089 2499 75147 2505
rect 75089 2496 75101 2499
rect 75052 2468 75101 2496
rect 75052 2456 75058 2468
rect 75089 2465 75101 2468
rect 75135 2465 75147 2499
rect 75089 2459 75147 2465
rect 75273 2499 75331 2505
rect 75273 2465 75285 2499
rect 75319 2496 75331 2499
rect 76561 2499 76619 2505
rect 76561 2496 76573 2499
rect 75319 2468 76573 2496
rect 75319 2465 75331 2468
rect 75273 2459 75331 2465
rect 76561 2465 76573 2468
rect 76607 2496 76619 2499
rect 77849 2499 77907 2505
rect 77849 2496 77861 2499
rect 76607 2468 77861 2496
rect 76607 2465 76619 2468
rect 76561 2459 76619 2465
rect 77849 2465 77861 2468
rect 77895 2496 77907 2499
rect 79226 2496 79232 2508
rect 77895 2468 79232 2496
rect 77895 2465 77907 2468
rect 77849 2459 77907 2465
rect 79226 2456 79232 2468
rect 79284 2456 79290 2508
rect 81526 2496 81532 2508
rect 79336 2468 81388 2496
rect 81487 2468 81532 2496
rect 79336 2428 79364 2468
rect 73632 2400 79364 2428
rect 79410 2388 79416 2440
rect 79468 2428 79474 2440
rect 80057 2431 80115 2437
rect 80057 2428 80069 2431
rect 79468 2400 80069 2428
rect 79468 2388 79474 2400
rect 80057 2397 80069 2400
rect 80103 2397 80115 2431
rect 80057 2391 80115 2397
rect 72528 2332 73844 2360
rect 72421 2323 72479 2329
rect 71133 2295 71191 2301
rect 71133 2292 71145 2295
rect 70366 2264 71145 2292
rect 70213 2255 70271 2261
rect 71133 2261 71145 2264
rect 71179 2261 71191 2295
rect 72436 2292 72464 2323
rect 73338 2292 73344 2304
rect 72436 2264 73344 2292
rect 71133 2255 71191 2261
rect 73338 2252 73344 2264
rect 73396 2252 73402 2304
rect 73430 2252 73436 2304
rect 73488 2292 73494 2304
rect 73709 2295 73767 2301
rect 73709 2292 73721 2295
rect 73488 2264 73721 2292
rect 73488 2252 73494 2264
rect 73709 2261 73721 2264
rect 73755 2261 73767 2295
rect 73816 2292 73844 2332
rect 73890 2320 73896 2372
rect 73948 2360 73954 2372
rect 76098 2360 76104 2372
rect 73948 2332 76104 2360
rect 73948 2320 73954 2332
rect 76098 2320 76104 2332
rect 76156 2320 76162 2372
rect 76190 2320 76196 2372
rect 76248 2360 76254 2372
rect 76285 2363 76343 2369
rect 76285 2360 76297 2363
rect 76248 2332 76297 2360
rect 76248 2320 76254 2332
rect 76285 2329 76297 2332
rect 76331 2329 76343 2363
rect 76285 2323 76343 2329
rect 79137 2363 79195 2369
rect 79137 2329 79149 2363
rect 79183 2360 79195 2363
rect 81360 2360 81388 2468
rect 81526 2456 81532 2468
rect 81584 2456 81590 2508
rect 81713 2499 81771 2505
rect 81713 2465 81725 2499
rect 81759 2496 81771 2499
rect 83185 2499 83243 2505
rect 83185 2496 83197 2499
rect 81759 2468 83197 2496
rect 81759 2465 81771 2468
rect 81713 2459 81771 2465
rect 83185 2465 83197 2468
rect 83231 2465 83243 2499
rect 83185 2459 83243 2465
rect 81434 2388 81440 2440
rect 81492 2428 81498 2440
rect 83001 2431 83059 2437
rect 83001 2428 83013 2431
rect 81492 2400 83013 2428
rect 81492 2388 81498 2400
rect 83001 2397 83013 2400
rect 83047 2397 83059 2431
rect 83200 2428 83228 2459
rect 83550 2456 83556 2508
rect 83608 2496 83614 2508
rect 84105 2499 84163 2505
rect 84105 2496 84117 2499
rect 83608 2468 84117 2496
rect 83608 2456 83614 2468
rect 84105 2465 84117 2468
rect 84151 2465 84163 2499
rect 84105 2459 84163 2465
rect 84197 2499 84255 2505
rect 84197 2465 84209 2499
rect 84243 2465 84255 2499
rect 84197 2459 84255 2465
rect 84212 2428 84240 2459
rect 84930 2456 84936 2508
rect 84988 2496 84994 2508
rect 85301 2499 85359 2505
rect 85301 2496 85313 2499
rect 84988 2468 85313 2496
rect 84988 2456 84994 2468
rect 85301 2465 85313 2468
rect 85347 2465 85359 2499
rect 85301 2459 85359 2465
rect 85485 2499 85543 2505
rect 85485 2465 85497 2499
rect 85531 2496 85543 2499
rect 85574 2496 85580 2508
rect 85531 2468 85580 2496
rect 85531 2465 85543 2468
rect 85485 2459 85543 2465
rect 85574 2456 85580 2468
rect 85632 2456 85638 2508
rect 86402 2456 86408 2508
rect 86460 2496 86466 2508
rect 86681 2499 86739 2505
rect 86681 2496 86693 2499
rect 86460 2468 86693 2496
rect 86460 2456 86466 2468
rect 86681 2465 86693 2468
rect 86727 2465 86739 2499
rect 86681 2459 86739 2465
rect 86773 2499 86831 2505
rect 86773 2465 86785 2499
rect 86819 2496 86831 2499
rect 86862 2496 86868 2508
rect 86819 2468 86868 2496
rect 86819 2465 86831 2468
rect 86773 2459 86831 2465
rect 83200 2400 84240 2428
rect 83001 2391 83059 2397
rect 84102 2360 84108 2372
rect 79183 2332 79916 2360
rect 81360 2332 84108 2360
rect 79183 2329 79195 2332
rect 79137 2323 79195 2329
rect 74442 2292 74448 2304
rect 73816 2264 74448 2292
rect 73709 2255 73767 2261
rect 74442 2252 74448 2264
rect 74500 2252 74506 2304
rect 74994 2292 75000 2304
rect 74955 2264 75000 2292
rect 74994 2252 75000 2264
rect 75052 2252 75058 2304
rect 76377 2295 76435 2301
rect 76377 2261 76389 2295
rect 76423 2292 76435 2295
rect 76466 2292 76472 2304
rect 76423 2264 76472 2292
rect 76423 2261 76435 2264
rect 76377 2255 76435 2261
rect 76466 2252 76472 2264
rect 76524 2252 76530 2304
rect 77570 2292 77576 2304
rect 77531 2264 77576 2292
rect 77570 2252 77576 2264
rect 77628 2252 77634 2304
rect 77662 2252 77668 2304
rect 77720 2292 77726 2304
rect 79042 2292 79048 2304
rect 77720 2264 77765 2292
rect 79003 2264 79048 2292
rect 77720 2252 77726 2264
rect 79042 2252 79048 2264
rect 79100 2292 79106 2304
rect 79888 2301 79916 2332
rect 84102 2320 84108 2332
rect 84160 2320 84166 2372
rect 79689 2295 79747 2301
rect 79689 2292 79701 2295
rect 79100 2264 79701 2292
rect 79100 2252 79106 2264
rect 79689 2261 79701 2264
rect 79735 2261 79747 2295
rect 79689 2255 79747 2261
rect 79873 2295 79931 2301
rect 79873 2261 79885 2295
rect 79919 2261 79931 2295
rect 79873 2255 79931 2261
rect 80514 2252 80520 2304
rect 80572 2292 80578 2304
rect 80609 2295 80667 2301
rect 80609 2292 80621 2295
rect 80572 2264 80621 2292
rect 80572 2252 80578 2264
rect 80609 2261 80621 2264
rect 80655 2292 80667 2295
rect 81437 2295 81495 2301
rect 81437 2292 81449 2295
rect 80655 2264 81449 2292
rect 80655 2261 80667 2264
rect 80609 2255 80667 2261
rect 81437 2261 81449 2264
rect 81483 2292 81495 2295
rect 82081 2295 82139 2301
rect 82081 2292 82093 2295
rect 81483 2264 82093 2292
rect 81483 2261 81495 2264
rect 81437 2255 81495 2261
rect 82081 2261 82093 2264
rect 82127 2292 82139 2295
rect 82449 2295 82507 2301
rect 82449 2292 82461 2295
rect 82127 2264 82461 2292
rect 82127 2261 82139 2264
rect 82081 2255 82139 2261
rect 82449 2261 82461 2264
rect 82495 2261 82507 2295
rect 83090 2292 83096 2304
rect 83051 2264 83096 2292
rect 82449 2255 82507 2261
rect 83090 2252 83096 2264
rect 83148 2252 83154 2304
rect 84010 2292 84016 2304
rect 83971 2264 84016 2292
rect 84010 2252 84016 2264
rect 84068 2252 84074 2304
rect 84212 2292 84240 2400
rect 85022 2388 85028 2440
rect 85080 2428 85086 2440
rect 85209 2431 85267 2437
rect 85209 2428 85221 2431
rect 85080 2400 85221 2428
rect 85080 2388 85086 2400
rect 85209 2397 85221 2400
rect 85255 2397 85267 2431
rect 85592 2428 85620 2456
rect 86788 2428 86816 2459
rect 86862 2456 86868 2468
rect 86920 2456 86926 2508
rect 87782 2456 87788 2508
rect 87840 2496 87846 2508
rect 87969 2499 88027 2505
rect 87969 2496 87981 2499
rect 87840 2468 87981 2496
rect 87840 2456 87846 2468
rect 87969 2465 87981 2468
rect 88015 2465 88027 2499
rect 87969 2459 88027 2465
rect 88153 2499 88211 2505
rect 88153 2465 88165 2499
rect 88199 2465 88211 2499
rect 89254 2496 89260 2508
rect 89215 2468 89260 2496
rect 88153 2459 88211 2465
rect 85592 2400 86816 2428
rect 88168 2428 88196 2459
rect 89254 2456 89260 2468
rect 89312 2456 89318 2508
rect 89349 2499 89407 2505
rect 89349 2465 89361 2499
rect 89395 2465 89407 2499
rect 90542 2496 90548 2508
rect 90503 2468 90548 2496
rect 89349 2459 89407 2465
rect 89364 2428 89392 2459
rect 90542 2456 90548 2468
rect 90600 2456 90606 2508
rect 90729 2499 90787 2505
rect 90729 2465 90741 2499
rect 90775 2465 90787 2499
rect 90729 2459 90787 2465
rect 89438 2428 89444 2440
rect 88168 2400 89444 2428
rect 85209 2391 85267 2397
rect 89438 2388 89444 2400
rect 89496 2428 89502 2440
rect 90744 2428 90772 2459
rect 91554 2456 91560 2508
rect 91612 2496 91618 2508
rect 92017 2499 92075 2505
rect 92017 2496 92029 2499
rect 91612 2468 92029 2496
rect 91612 2456 91618 2468
rect 92017 2465 92029 2468
rect 92063 2465 92075 2499
rect 92017 2459 92075 2465
rect 92201 2499 92259 2505
rect 92201 2465 92213 2499
rect 92247 2496 92259 2499
rect 92290 2496 92296 2508
rect 92247 2468 92296 2496
rect 92247 2465 92259 2468
rect 92201 2459 92259 2465
rect 92216 2428 92244 2459
rect 92290 2456 92296 2468
rect 92348 2456 92354 2508
rect 95510 2496 95516 2508
rect 95471 2468 95516 2496
rect 95510 2456 95516 2468
rect 95568 2456 95574 2508
rect 95697 2499 95755 2505
rect 95697 2465 95709 2499
rect 95743 2465 95755 2499
rect 96982 2496 96988 2508
rect 96943 2468 96988 2496
rect 95697 2459 95755 2465
rect 92934 2428 92940 2440
rect 89496 2400 92244 2428
rect 92895 2400 92940 2428
rect 89496 2388 89502 2400
rect 92934 2388 92940 2400
rect 92992 2388 92998 2440
rect 93486 2388 93492 2440
rect 93544 2428 93550 2440
rect 94133 2431 94191 2437
rect 94133 2428 94145 2431
rect 93544 2400 94145 2428
rect 93544 2388 93550 2400
rect 94133 2397 94145 2400
rect 94179 2397 94191 2431
rect 95712 2428 95740 2459
rect 96982 2456 96988 2468
rect 97040 2456 97046 2508
rect 97169 2499 97227 2505
rect 97169 2465 97181 2499
rect 97215 2496 97227 2499
rect 97920 2496 97948 2592
rect 97215 2468 97948 2496
rect 97215 2465 97227 2468
rect 97169 2459 97227 2465
rect 97184 2428 97212 2459
rect 97994 2456 98000 2508
rect 98052 2496 98058 2508
rect 98181 2499 98239 2505
rect 98181 2496 98193 2499
rect 98052 2468 98193 2496
rect 98052 2456 98058 2468
rect 98181 2465 98193 2468
rect 98227 2465 98239 2499
rect 98181 2459 98239 2465
rect 98365 2499 98423 2505
rect 98365 2465 98377 2499
rect 98411 2496 98423 2499
rect 98472 2496 98500 2604
rect 99760 2576 99788 2604
rect 100294 2592 100300 2604
rect 100352 2592 100358 2644
rect 101677 2635 101735 2641
rect 101677 2601 101689 2635
rect 101723 2632 101735 2635
rect 102134 2632 102140 2644
rect 101723 2604 102140 2632
rect 101723 2601 101735 2604
rect 101677 2595 101735 2601
rect 102134 2592 102140 2604
rect 102192 2592 102198 2644
rect 102873 2635 102931 2641
rect 102873 2601 102885 2635
rect 102919 2632 102931 2635
rect 104250 2632 104256 2644
rect 102919 2604 104256 2632
rect 102919 2601 102931 2604
rect 102873 2595 102931 2601
rect 104250 2592 104256 2604
rect 104308 2592 104314 2644
rect 105081 2635 105139 2641
rect 105081 2601 105093 2635
rect 105127 2632 105139 2635
rect 105814 2632 105820 2644
rect 105127 2604 105820 2632
rect 105127 2601 105139 2604
rect 105081 2595 105139 2601
rect 105814 2592 105820 2604
rect 105872 2592 105878 2644
rect 107289 2635 107347 2641
rect 107289 2601 107301 2635
rect 107335 2632 107347 2635
rect 108298 2632 108304 2644
rect 107335 2604 108304 2632
rect 107335 2601 107347 2604
rect 107289 2595 107347 2601
rect 108298 2592 108304 2604
rect 108356 2592 108362 2644
rect 110506 2592 110512 2644
rect 110564 2632 110570 2644
rect 111061 2635 111119 2641
rect 111061 2632 111073 2635
rect 110564 2604 111073 2632
rect 110564 2592 110570 2604
rect 111061 2601 111073 2604
rect 111107 2601 111119 2635
rect 111061 2595 111119 2601
rect 111981 2635 112039 2641
rect 111981 2601 111993 2635
rect 112027 2632 112039 2635
rect 114094 2632 114100 2644
rect 112027 2604 114100 2632
rect 112027 2601 112039 2604
rect 111981 2595 112039 2601
rect 114094 2592 114100 2604
rect 114152 2592 114158 2644
rect 114925 2635 114983 2641
rect 114925 2601 114937 2635
rect 114971 2632 114983 2635
rect 116578 2632 116584 2644
rect 114971 2604 116584 2632
rect 114971 2601 114983 2604
rect 114925 2595 114983 2601
rect 116578 2592 116584 2604
rect 116636 2592 116642 2644
rect 99098 2564 99104 2576
rect 99059 2536 99104 2564
rect 99098 2524 99104 2536
rect 99156 2524 99162 2576
rect 99558 2524 99564 2576
rect 99616 2564 99622 2576
rect 99616 2536 99696 2564
rect 99616 2524 99622 2536
rect 99668 2505 99696 2536
rect 99742 2524 99748 2576
rect 99800 2564 99806 2576
rect 99800 2536 100892 2564
rect 99800 2524 99806 2536
rect 98411 2468 98500 2496
rect 99653 2499 99711 2505
rect 98411 2465 98423 2468
rect 98365 2459 98423 2465
rect 99653 2465 99665 2499
rect 99699 2465 99711 2499
rect 100294 2496 100300 2508
rect 99653 2459 99711 2465
rect 99760 2468 100300 2496
rect 95712 2400 97212 2428
rect 99561 2431 99619 2437
rect 94133 2391 94191 2397
rect 99561 2397 99573 2431
rect 99607 2428 99619 2431
rect 99760 2428 99788 2468
rect 100294 2456 100300 2468
rect 100352 2456 100358 2508
rect 100386 2456 100392 2508
rect 100444 2496 100450 2508
rect 100864 2505 100892 2536
rect 106182 2524 106188 2576
rect 106240 2564 106246 2576
rect 109405 2567 109463 2573
rect 106240 2536 107884 2564
rect 106240 2524 106246 2536
rect 100757 2499 100815 2505
rect 100757 2496 100769 2499
rect 100444 2468 100769 2496
rect 100444 2456 100450 2468
rect 100757 2465 100769 2468
rect 100803 2465 100815 2499
rect 100757 2459 100815 2465
rect 100849 2499 100907 2505
rect 100849 2465 100861 2499
rect 100895 2465 100907 2499
rect 102318 2496 102324 2508
rect 102231 2468 102324 2496
rect 100849 2459 100907 2465
rect 102318 2456 102324 2468
rect 102376 2496 102382 2508
rect 103514 2496 103520 2508
rect 102376 2468 103520 2496
rect 102376 2456 102382 2468
rect 103514 2456 103520 2468
rect 103572 2456 103578 2508
rect 104360 2468 105124 2496
rect 99607 2400 99788 2428
rect 102137 2431 102195 2437
rect 99607 2397 99619 2400
rect 99561 2391 99619 2397
rect 102137 2397 102149 2431
rect 102183 2428 102195 2431
rect 102962 2428 102968 2440
rect 102183 2400 102968 2428
rect 102183 2397 102195 2400
rect 102137 2391 102195 2397
rect 102962 2388 102968 2400
rect 103020 2388 103026 2440
rect 104360 2428 104388 2468
rect 103348 2400 104388 2428
rect 104437 2431 104495 2437
rect 84286 2320 84292 2372
rect 84344 2360 84350 2372
rect 84344 2332 99374 2360
rect 84344 2320 84350 2332
rect 85574 2292 85580 2304
rect 84212 2264 85580 2292
rect 85574 2252 85580 2264
rect 85632 2252 85638 2304
rect 86586 2292 86592 2304
rect 86547 2264 86592 2292
rect 86586 2252 86592 2264
rect 86644 2252 86650 2304
rect 87874 2292 87880 2304
rect 87835 2264 87880 2292
rect 87874 2252 87880 2264
rect 87932 2252 87938 2304
rect 88334 2252 88340 2304
rect 88392 2292 88398 2304
rect 89165 2295 89223 2301
rect 89165 2292 89177 2295
rect 88392 2264 89177 2292
rect 88392 2252 88398 2264
rect 89165 2261 89177 2264
rect 89211 2261 89223 2295
rect 90450 2292 90456 2304
rect 90411 2264 90456 2292
rect 89165 2255 89223 2261
rect 90450 2252 90456 2264
rect 90508 2252 90514 2304
rect 91922 2292 91928 2304
rect 91883 2264 91928 2292
rect 91922 2252 91928 2264
rect 91980 2252 91986 2304
rect 95418 2292 95424 2304
rect 95379 2264 95424 2292
rect 95418 2252 95424 2264
rect 95476 2252 95482 2304
rect 96890 2292 96896 2304
rect 96851 2264 96896 2292
rect 96890 2252 96896 2264
rect 96948 2252 96954 2304
rect 98086 2292 98092 2304
rect 98047 2264 98092 2292
rect 98086 2252 98092 2264
rect 98144 2252 98150 2304
rect 99346 2292 99374 2332
rect 99466 2320 99472 2372
rect 99524 2360 99530 2372
rect 100113 2363 100171 2369
rect 100113 2360 100125 2363
rect 99524 2332 100125 2360
rect 99524 2320 99530 2332
rect 100113 2329 100125 2332
rect 100159 2329 100171 2363
rect 103348 2360 103376 2400
rect 104437 2397 104449 2431
rect 104483 2397 104495 2431
rect 104437 2391 104495 2397
rect 100113 2323 100171 2329
rect 100496 2332 103376 2360
rect 100496 2292 100524 2332
rect 103422 2320 103428 2372
rect 103480 2360 103486 2372
rect 104452 2360 104480 2391
rect 103480 2332 104480 2360
rect 103480 2320 103486 2332
rect 100662 2292 100668 2304
rect 99346 2264 100524 2292
rect 100623 2264 100668 2292
rect 100662 2252 100668 2264
rect 100720 2252 100726 2304
rect 100754 2252 100760 2304
rect 100812 2292 100818 2304
rect 102045 2295 102103 2301
rect 102045 2292 102057 2295
rect 100812 2264 102057 2292
rect 100812 2252 100818 2264
rect 102045 2261 102057 2264
rect 102091 2261 102103 2295
rect 103238 2292 103244 2304
rect 103199 2264 103244 2292
rect 102045 2255 102103 2261
rect 103238 2252 103244 2264
rect 103296 2252 103302 2304
rect 103333 2295 103391 2301
rect 103333 2261 103345 2295
rect 103379 2292 103391 2295
rect 104253 2295 104311 2301
rect 104253 2292 104265 2295
rect 103379 2264 104265 2292
rect 103379 2261 103391 2264
rect 103333 2255 103391 2261
rect 104253 2261 104265 2264
rect 104299 2261 104311 2295
rect 105096 2292 105124 2468
rect 105170 2456 105176 2508
rect 105228 2496 105234 2508
rect 105541 2499 105599 2505
rect 105541 2496 105553 2499
rect 105228 2468 105553 2496
rect 105228 2456 105234 2468
rect 105541 2465 105553 2468
rect 105587 2465 105599 2499
rect 105541 2459 105599 2465
rect 105633 2499 105691 2505
rect 105633 2465 105645 2499
rect 105679 2465 105691 2499
rect 105633 2459 105691 2465
rect 105446 2428 105452 2440
rect 105407 2400 105452 2428
rect 105446 2388 105452 2400
rect 105504 2388 105510 2440
rect 105648 2360 105676 2459
rect 107654 2456 107660 2508
rect 107712 2496 107718 2508
rect 107856 2505 107884 2536
rect 109405 2533 109417 2567
rect 109451 2564 109463 2567
rect 110690 2564 110696 2576
rect 109451 2536 110696 2564
rect 109451 2533 109463 2536
rect 109405 2527 109463 2533
rect 110690 2524 110696 2536
rect 110748 2524 110754 2576
rect 113269 2567 113327 2573
rect 113269 2533 113281 2567
rect 113315 2564 113327 2567
rect 115842 2564 115848 2576
rect 113315 2536 115848 2564
rect 113315 2533 113327 2536
rect 113269 2527 113327 2533
rect 115842 2524 115848 2536
rect 115900 2524 115906 2576
rect 107749 2499 107807 2505
rect 107749 2496 107761 2499
rect 107712 2468 107761 2496
rect 107712 2456 107718 2468
rect 107749 2465 107761 2468
rect 107795 2465 107807 2499
rect 107749 2459 107807 2465
rect 107841 2499 107899 2505
rect 107841 2465 107853 2499
rect 107887 2496 107899 2499
rect 108853 2499 108911 2505
rect 108853 2496 108865 2499
rect 107887 2468 108865 2496
rect 107887 2465 107899 2468
rect 107841 2459 107899 2465
rect 108853 2465 108865 2468
rect 108899 2496 108911 2499
rect 109954 2496 109960 2508
rect 108899 2468 109960 2496
rect 108899 2465 108911 2468
rect 108853 2459 108911 2465
rect 109954 2456 109960 2468
rect 110012 2456 110018 2508
rect 110598 2456 110604 2508
rect 110656 2496 110662 2508
rect 110656 2468 111288 2496
rect 110656 2456 110662 2468
rect 105722 2388 105728 2440
rect 105780 2428 105786 2440
rect 109034 2428 109040 2440
rect 105780 2400 109040 2428
rect 105780 2388 105786 2400
rect 109034 2388 109040 2400
rect 109092 2388 109098 2440
rect 109126 2388 109132 2440
rect 109184 2428 109190 2440
rect 111260 2437 111288 2468
rect 112070 2456 112076 2508
rect 112128 2496 112134 2508
rect 112441 2499 112499 2505
rect 112441 2496 112453 2499
rect 112128 2468 112453 2496
rect 112128 2456 112134 2468
rect 112441 2465 112453 2468
rect 112487 2465 112499 2499
rect 112622 2496 112628 2508
rect 112583 2468 112628 2496
rect 112441 2459 112499 2465
rect 112622 2456 112628 2468
rect 112680 2496 112686 2508
rect 112680 2468 113174 2496
rect 112680 2456 112686 2468
rect 110785 2431 110843 2437
rect 110785 2428 110797 2431
rect 109184 2400 110797 2428
rect 109184 2388 109190 2400
rect 110785 2397 110797 2400
rect 110831 2397 110843 2431
rect 110785 2391 110843 2397
rect 111245 2431 111303 2437
rect 111245 2397 111257 2431
rect 111291 2397 111303 2431
rect 113146 2428 113174 2468
rect 113542 2456 113548 2508
rect 113600 2496 113606 2508
rect 113729 2499 113787 2505
rect 113729 2496 113741 2499
rect 113600 2468 113741 2496
rect 113600 2456 113606 2468
rect 113729 2465 113741 2468
rect 113775 2465 113787 2499
rect 113729 2459 113787 2465
rect 113821 2499 113879 2505
rect 113821 2465 113833 2499
rect 113867 2465 113879 2499
rect 115382 2496 115388 2508
rect 115343 2468 115388 2496
rect 113821 2459 113879 2465
rect 113836 2428 113864 2459
rect 115382 2456 115388 2468
rect 115440 2456 115446 2508
rect 115474 2456 115480 2508
rect 115532 2496 115538 2508
rect 117317 2499 117375 2505
rect 115532 2468 115625 2496
rect 115532 2456 115538 2468
rect 117317 2465 117329 2499
rect 117363 2496 117375 2499
rect 119154 2496 119160 2508
rect 117363 2468 119160 2496
rect 117363 2465 117375 2468
rect 117317 2459 117375 2465
rect 119154 2456 119160 2468
rect 119212 2456 119218 2508
rect 115492 2428 115520 2456
rect 116486 2428 116492 2440
rect 113146 2400 115520 2428
rect 116447 2400 116492 2428
rect 111245 2391 111303 2397
rect 116486 2388 116492 2400
rect 116544 2388 116550 2440
rect 117590 2428 117596 2440
rect 117551 2400 117596 2428
rect 117590 2388 117596 2400
rect 117648 2388 117654 2440
rect 106182 2360 106188 2372
rect 105648 2332 106188 2360
rect 106182 2320 106188 2332
rect 106240 2320 106246 2372
rect 108666 2360 108672 2372
rect 108627 2332 108672 2360
rect 108666 2320 108672 2332
rect 108724 2360 108730 2372
rect 112530 2360 112536 2372
rect 108724 2332 112536 2360
rect 108724 2320 108730 2332
rect 112530 2320 112536 2332
rect 112588 2320 112594 2372
rect 113634 2360 113640 2372
rect 113547 2332 113640 2360
rect 113634 2320 113640 2332
rect 113692 2360 113698 2372
rect 115937 2363 115995 2369
rect 115937 2360 115949 2363
rect 113692 2332 115949 2360
rect 113692 2320 113698 2332
rect 115937 2329 115949 2332
rect 115983 2329 115995 2363
rect 116762 2360 116768 2372
rect 116723 2332 116768 2360
rect 115937 2323 115995 2329
rect 116762 2320 116768 2332
rect 116820 2320 116826 2372
rect 107657 2295 107715 2301
rect 107657 2292 107669 2295
rect 105096 2264 107669 2292
rect 104253 2255 104311 2261
rect 107657 2261 107669 2264
rect 107703 2292 107715 2295
rect 108301 2295 108359 2301
rect 108301 2292 108313 2295
rect 107703 2264 108313 2292
rect 107703 2261 107715 2264
rect 107657 2255 107715 2261
rect 108301 2261 108313 2264
rect 108347 2261 108359 2295
rect 109770 2292 109776 2304
rect 109731 2264 109776 2292
rect 108301 2255 108359 2261
rect 109770 2252 109776 2264
rect 109828 2252 109834 2304
rect 109865 2295 109923 2301
rect 109865 2261 109877 2295
rect 109911 2292 109923 2295
rect 110601 2295 110659 2301
rect 110601 2292 110613 2295
rect 109911 2264 110613 2292
rect 109911 2261 109923 2264
rect 109865 2255 109923 2261
rect 110601 2261 110613 2264
rect 110647 2261 110659 2295
rect 111518 2292 111524 2304
rect 111479 2264 111524 2292
rect 110601 2255 110659 2261
rect 111518 2252 111524 2264
rect 111576 2292 111582 2304
rect 112349 2295 112407 2301
rect 112349 2292 112361 2295
rect 111576 2264 112361 2292
rect 111576 2252 111582 2264
rect 112349 2261 112361 2264
rect 112395 2261 112407 2295
rect 115290 2292 115296 2304
rect 115251 2264 115296 2292
rect 112349 2255 112407 2261
rect 115290 2252 115296 2264
rect 115348 2292 115354 2304
rect 116305 2295 116363 2301
rect 116305 2292 116317 2295
rect 115348 2264 116317 2292
rect 115348 2252 115354 2264
rect 116305 2261 116317 2264
rect 116351 2261 116363 2295
rect 116305 2255 116363 2261
rect 1104 2202 118864 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 81014 2202
rect 81066 2150 81078 2202
rect 81130 2150 81142 2202
rect 81194 2150 81206 2202
rect 81258 2150 81270 2202
rect 81322 2150 111734 2202
rect 111786 2150 111798 2202
rect 111850 2150 111862 2202
rect 111914 2150 111926 2202
rect 111978 2150 111990 2202
rect 112042 2150 118864 2202
rect 1104 2128 118864 2150
rect 2130 2048 2136 2100
rect 2188 2088 2194 2100
rect 51074 2088 51080 2100
rect 2188 2060 51080 2088
rect 2188 2048 2194 2060
rect 51074 2048 51080 2060
rect 51132 2048 51138 2100
rect 60182 2088 60188 2100
rect 51276 2060 60188 2088
rect 3786 1980 3792 2032
rect 3844 2020 3850 2032
rect 51276 2020 51304 2060
rect 60182 2048 60188 2060
rect 60240 2048 60246 2100
rect 60366 2048 60372 2100
rect 60424 2088 60430 2100
rect 66806 2088 66812 2100
rect 60424 2060 66812 2088
rect 60424 2048 60430 2060
rect 66806 2048 66812 2060
rect 66864 2048 66870 2100
rect 66898 2048 66904 2100
rect 66956 2088 66962 2100
rect 113634 2088 113640 2100
rect 66956 2060 113640 2088
rect 66956 2048 66962 2060
rect 113634 2048 113640 2060
rect 113692 2048 113698 2100
rect 3844 1992 51304 2020
rect 3844 1980 3850 1992
rect 51350 1980 51356 2032
rect 51408 2020 51414 2032
rect 59814 2020 59820 2032
rect 51408 1992 59820 2020
rect 51408 1980 51414 1992
rect 59814 1980 59820 1992
rect 59872 1980 59878 2032
rect 60706 1992 60964 2020
rect 24762 1912 24768 1964
rect 24820 1952 24826 1964
rect 60706 1952 60734 1992
rect 24820 1924 60734 1952
rect 60936 1952 60964 1992
rect 61930 1980 61936 2032
rect 61988 2020 61994 2032
rect 111518 2020 111524 2032
rect 61988 1992 111524 2020
rect 61988 1980 61994 1992
rect 111518 1980 111524 1992
rect 111576 1980 111582 2032
rect 76006 1952 76012 1964
rect 60936 1924 76012 1952
rect 24820 1912 24826 1924
rect 76006 1912 76012 1924
rect 76064 1912 76070 1964
rect 76098 1912 76104 1964
rect 76156 1952 76162 1964
rect 80514 1952 80520 1964
rect 76156 1924 80520 1952
rect 76156 1912 76162 1924
rect 80514 1912 80520 1924
rect 80572 1912 80578 1964
rect 80882 1912 80888 1964
rect 80940 1952 80946 1964
rect 84746 1952 84752 1964
rect 80940 1924 84752 1952
rect 80940 1912 80946 1924
rect 84746 1912 84752 1924
rect 84804 1912 84810 1964
rect 103514 1912 103520 1964
rect 103572 1952 103578 1964
rect 108666 1952 108672 1964
rect 103572 1924 108672 1952
rect 103572 1912 103578 1924
rect 108666 1912 108672 1924
rect 108724 1912 108730 1964
rect 19426 1844 19432 1896
rect 19484 1884 19490 1896
rect 25774 1884 25780 1896
rect 19484 1856 25780 1884
rect 19484 1844 19490 1856
rect 25774 1844 25780 1856
rect 25832 1844 25838 1896
rect 26234 1844 26240 1896
rect 26292 1884 26298 1896
rect 35618 1884 35624 1896
rect 26292 1856 35624 1884
rect 26292 1844 26298 1856
rect 35618 1844 35624 1856
rect 35676 1844 35682 1896
rect 60734 1884 60740 1896
rect 35728 1856 60740 1884
rect 27338 1776 27344 1828
rect 27396 1816 27402 1828
rect 35728 1816 35756 1856
rect 60734 1844 60740 1856
rect 60792 1844 60798 1896
rect 60918 1844 60924 1896
rect 60976 1884 60982 1896
rect 60976 1856 79272 1884
rect 60976 1844 60982 1856
rect 27396 1788 35756 1816
rect 27396 1776 27402 1788
rect 35802 1776 35808 1828
rect 35860 1816 35866 1828
rect 79134 1816 79140 1828
rect 35860 1788 79140 1816
rect 35860 1776 35866 1788
rect 79134 1776 79140 1788
rect 79192 1776 79198 1828
rect 19978 1708 19984 1760
rect 20036 1748 20042 1760
rect 79042 1748 79048 1760
rect 20036 1720 79048 1748
rect 20036 1708 20042 1720
rect 79042 1708 79048 1720
rect 79100 1708 79106 1760
rect 79244 1748 79272 1856
rect 79318 1844 79324 1896
rect 79376 1884 79382 1896
rect 79376 1856 79456 1884
rect 79376 1844 79382 1856
rect 79428 1816 79456 1856
rect 79502 1844 79508 1896
rect 79560 1884 79566 1896
rect 91462 1884 91468 1896
rect 79560 1856 91468 1884
rect 79560 1844 79566 1856
rect 91462 1844 91468 1856
rect 91520 1844 91526 1896
rect 100294 1844 100300 1896
rect 100352 1884 100358 1896
rect 117590 1884 117596 1896
rect 100352 1856 117596 1884
rect 100352 1844 100358 1856
rect 117590 1844 117596 1856
rect 117648 1844 117654 1896
rect 87874 1816 87880 1828
rect 79428 1788 87880 1816
rect 87874 1776 87880 1788
rect 87932 1776 87938 1828
rect 86586 1748 86592 1760
rect 79244 1720 86592 1748
rect 86586 1708 86592 1720
rect 86644 1708 86650 1760
rect 10686 1640 10692 1692
rect 10744 1680 10750 1692
rect 63310 1680 63316 1692
rect 10744 1652 63316 1680
rect 10744 1640 10750 1652
rect 63310 1640 63316 1652
rect 63368 1640 63374 1692
rect 66162 1640 66168 1692
rect 66220 1680 66226 1692
rect 70210 1680 70216 1692
rect 66220 1652 70216 1680
rect 66220 1640 66226 1652
rect 70210 1640 70216 1652
rect 70268 1640 70274 1692
rect 70302 1640 70308 1692
rect 70360 1680 70366 1692
rect 73890 1680 73896 1692
rect 70360 1652 73896 1680
rect 70360 1640 70366 1652
rect 73890 1640 73896 1652
rect 73948 1640 73954 1692
rect 73982 1640 73988 1692
rect 74040 1680 74046 1692
rect 99466 1680 99472 1692
rect 74040 1652 99472 1680
rect 74040 1640 74046 1652
rect 99466 1640 99472 1652
rect 99524 1640 99530 1692
rect 12158 1572 12164 1624
rect 12216 1612 12222 1624
rect 45554 1612 45560 1624
rect 12216 1584 45560 1612
rect 12216 1572 12222 1584
rect 45554 1572 45560 1584
rect 45612 1572 45618 1624
rect 45646 1572 45652 1624
rect 45704 1612 45710 1624
rect 99374 1612 99380 1624
rect 45704 1584 60780 1612
rect 45704 1572 45710 1584
rect 7834 1504 7840 1556
rect 7892 1544 7898 1556
rect 51074 1544 51080 1556
rect 7892 1516 51080 1544
rect 7892 1504 7898 1516
rect 51074 1504 51080 1516
rect 51132 1504 51138 1556
rect 51258 1504 51264 1556
rect 51316 1544 51322 1556
rect 60550 1544 60556 1556
rect 51316 1516 60556 1544
rect 51316 1504 51322 1516
rect 60550 1504 60556 1516
rect 60608 1504 60614 1556
rect 60752 1544 60780 1584
rect 60936 1584 99380 1612
rect 60936 1544 60964 1584
rect 99374 1572 99380 1584
rect 99432 1572 99438 1624
rect 60752 1516 60964 1544
rect 61746 1504 61752 1556
rect 61804 1544 61810 1556
rect 115290 1544 115296 1556
rect 61804 1516 115296 1544
rect 61804 1504 61810 1516
rect 115290 1504 115296 1516
rect 115348 1504 115354 1556
rect 14090 1436 14096 1488
rect 14148 1476 14154 1488
rect 45646 1476 45652 1488
rect 14148 1448 45652 1476
rect 14148 1436 14154 1448
rect 45646 1436 45652 1448
rect 45704 1436 45710 1488
rect 45738 1436 45744 1488
rect 45796 1476 45802 1488
rect 51166 1476 51172 1488
rect 45796 1448 51172 1476
rect 45796 1436 45802 1448
rect 51166 1436 51172 1448
rect 51224 1436 51230 1488
rect 51626 1436 51632 1488
rect 51684 1476 51690 1488
rect 60458 1476 60464 1488
rect 51684 1448 60464 1476
rect 51684 1436 51690 1448
rect 60458 1436 60464 1448
rect 60516 1436 60522 1488
rect 61010 1436 61016 1488
rect 61068 1476 61074 1488
rect 105262 1476 105268 1488
rect 61068 1448 105268 1476
rect 61068 1436 61074 1448
rect 105262 1436 105268 1448
rect 105320 1436 105326 1488
rect 7098 1368 7104 1420
rect 7156 1408 7162 1420
rect 51258 1408 51264 1420
rect 7156 1380 51264 1408
rect 7156 1368 7162 1380
rect 51258 1368 51264 1380
rect 51316 1368 51322 1420
rect 60734 1408 60740 1420
rect 51552 1380 60740 1408
rect 45554 1300 45560 1352
rect 45612 1340 45618 1352
rect 51552 1340 51580 1380
rect 60734 1368 60740 1380
rect 60792 1368 60798 1420
rect 61194 1368 61200 1420
rect 61252 1408 61258 1420
rect 72786 1408 72792 1420
rect 61252 1380 72792 1408
rect 61252 1368 61258 1380
rect 72786 1368 72792 1380
rect 72844 1368 72850 1420
rect 72878 1368 72884 1420
rect 72936 1408 72942 1420
rect 77570 1408 77576 1420
rect 72936 1380 77576 1408
rect 72936 1368 72942 1380
rect 77570 1368 77576 1380
rect 77628 1368 77634 1420
rect 77662 1368 77668 1420
rect 77720 1408 77726 1420
rect 84010 1408 84016 1420
rect 77720 1380 84016 1408
rect 77720 1368 77726 1380
rect 84010 1368 84016 1380
rect 84068 1368 84074 1420
rect 84746 1368 84752 1420
rect 84804 1408 84810 1420
rect 98454 1408 98460 1420
rect 84804 1380 98460 1408
rect 84804 1368 84810 1380
rect 98454 1368 98460 1380
rect 98512 1368 98518 1420
rect 99190 1368 99196 1420
rect 99248 1408 99254 1420
rect 101214 1408 101220 1420
rect 99248 1380 101220 1408
rect 99248 1368 99254 1380
rect 101214 1368 101220 1380
rect 101272 1368 101278 1420
rect 45612 1312 51580 1340
rect 45612 1300 45618 1312
rect 56318 1300 56324 1352
rect 56376 1340 56382 1352
rect 61746 1340 61752 1352
rect 56376 1312 61752 1340
rect 56376 1300 56382 1312
rect 61746 1300 61752 1312
rect 61804 1300 61810 1352
rect 65518 1300 65524 1352
rect 65576 1340 65582 1352
rect 109770 1340 109776 1352
rect 65576 1312 109776 1340
rect 65576 1300 65582 1312
rect 109770 1300 109776 1312
rect 109828 1300 109834 1352
rect 35526 1232 35532 1284
rect 35584 1272 35590 1284
rect 95418 1272 95424 1284
rect 35584 1244 95424 1272
rect 35584 1232 35590 1244
rect 95418 1232 95424 1244
rect 95476 1232 95482 1284
rect 45646 1164 45652 1216
rect 45704 1204 45710 1216
rect 51626 1204 51632 1216
rect 45704 1176 51632 1204
rect 45704 1164 45710 1176
rect 51626 1164 51632 1176
rect 51684 1164 51690 1216
rect 61378 1164 61384 1216
rect 61436 1204 61442 1216
rect 116762 1204 116768 1216
rect 61436 1176 116768 1204
rect 61436 1164 61442 1176
rect 116762 1164 116768 1176
rect 116820 1164 116826 1216
rect 38562 1096 38568 1148
rect 38620 1136 38626 1148
rect 98086 1136 98092 1148
rect 38620 1108 98092 1136
rect 38620 1096 38626 1108
rect 98086 1096 98092 1108
rect 98144 1096 98150 1148
rect 41138 1028 41144 1080
rect 41196 1068 41202 1080
rect 100662 1068 100668 1080
rect 41196 1040 100668 1068
rect 41196 1028 41202 1040
rect 100662 1028 100668 1040
rect 100720 1028 100726 1080
rect 32582 960 32588 1012
rect 32640 1000 32646 1012
rect 91922 1000 91928 1012
rect 32640 972 91928 1000
rect 32640 960 32646 972
rect 91922 960 91928 972
rect 91980 960 91986 1012
rect 31662 892 31668 944
rect 31720 932 31726 944
rect 90450 932 90456 944
rect 31720 904 90456 932
rect 31720 892 31726 904
rect 90450 892 90456 904
rect 90508 892 90514 944
rect 43898 824 43904 876
rect 43956 864 43962 876
rect 103238 864 103244 876
rect 43956 836 103244 864
rect 43956 824 43962 836
rect 103238 824 103244 836
rect 103296 824 103302 876
rect 30006 756 30012 808
rect 30064 796 30070 808
rect 88334 796 88340 808
rect 30064 768 88340 796
rect 30064 756 30070 768
rect 88334 756 88340 768
rect 88392 756 88398 808
rect 37642 688 37648 740
rect 37700 728 37706 740
rect 96890 728 96896 740
rect 37700 700 96896 728
rect 37700 688 37706 700
rect 96890 688 96896 700
rect 96948 688 96954 740
rect 42794 620 42800 672
rect 42852 660 42858 672
rect 100754 660 100760 672
rect 42852 632 100760 660
rect 42852 620 42858 632
rect 100754 620 100760 632
rect 100812 620 100818 672
rect 18322 552 18328 604
rect 18380 592 18386 604
rect 72878 592 72884 604
rect 18380 564 72884 592
rect 18380 552 18386 564
rect 72878 552 72884 564
rect 72936 552 72942 604
rect 15470 484 15476 536
rect 15528 524 15534 536
rect 74994 524 75000 536
rect 15528 496 75000 524
rect 15528 484 15534 496
rect 74994 484 75000 496
rect 75052 484 75058 536
rect 49602 348 49608 400
rect 49660 388 49666 400
rect 65518 388 65524 400
rect 49660 360 65524 388
rect 49660 348 49666 360
rect 65518 348 65524 360
rect 65576 348 65582 400
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 96374 37510 96426 37562
rect 96438 37510 96490 37562
rect 96502 37510 96554 37562
rect 96566 37510 96618 37562
rect 96630 37510 96682 37562
rect 117228 37408 117280 37460
rect 118056 37451 118108 37460
rect 118056 37417 118065 37451
rect 118065 37417 118099 37451
rect 118099 37417 118108 37451
rect 118056 37408 118108 37417
rect 114928 37204 114980 37256
rect 117596 37204 117648 37256
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 81014 36966 81066 37018
rect 81078 36966 81130 37018
rect 81142 36966 81194 37018
rect 81206 36966 81258 37018
rect 81270 36966 81322 37018
rect 111734 36966 111786 37018
rect 111798 36966 111850 37018
rect 111862 36966 111914 37018
rect 111926 36966 111978 37018
rect 111990 36966 112042 37018
rect 117136 36864 117188 36916
rect 98920 36728 98972 36780
rect 118424 36728 118476 36780
rect 118056 36635 118108 36644
rect 118056 36601 118065 36635
rect 118065 36601 118099 36635
rect 118099 36601 118108 36635
rect 118056 36592 118108 36601
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 96374 36422 96426 36474
rect 96438 36422 96490 36474
rect 96502 36422 96554 36474
rect 96566 36422 96618 36474
rect 96630 36422 96682 36474
rect 118148 36116 118200 36168
rect 118056 36023 118108 36032
rect 118056 35989 118065 36023
rect 118065 35989 118099 36023
rect 118099 35989 118108 36023
rect 118056 35980 118108 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 81014 35878 81066 35930
rect 81078 35878 81130 35930
rect 81142 35878 81194 35930
rect 81206 35878 81258 35930
rect 81270 35878 81322 35930
rect 111734 35878 111786 35930
rect 111798 35878 111850 35930
rect 111862 35878 111914 35930
rect 111926 35878 111978 35930
rect 111990 35878 112042 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 96374 35334 96426 35386
rect 96438 35334 96490 35386
rect 96502 35334 96554 35386
rect 96566 35334 96618 35386
rect 96630 35334 96682 35386
rect 117688 35028 117740 35080
rect 118056 34935 118108 34944
rect 118056 34901 118065 34935
rect 118065 34901 118099 34935
rect 118099 34901 118108 34935
rect 118056 34892 118108 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 81014 34790 81066 34842
rect 81078 34790 81130 34842
rect 81142 34790 81194 34842
rect 81206 34790 81258 34842
rect 81270 34790 81322 34842
rect 111734 34790 111786 34842
rect 111798 34790 111850 34842
rect 111862 34790 111914 34842
rect 111926 34790 111978 34842
rect 111990 34790 112042 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 96374 34246 96426 34298
rect 96438 34246 96490 34298
rect 96502 34246 96554 34298
rect 96566 34246 96618 34298
rect 96630 34246 96682 34298
rect 112168 33940 112220 33992
rect 118056 33847 118108 33856
rect 118056 33813 118065 33847
rect 118065 33813 118099 33847
rect 118099 33813 118108 33847
rect 118056 33804 118108 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 81014 33702 81066 33754
rect 81078 33702 81130 33754
rect 81142 33702 81194 33754
rect 81206 33702 81258 33754
rect 81270 33702 81322 33754
rect 111734 33702 111786 33754
rect 111798 33702 111850 33754
rect 111862 33702 111914 33754
rect 111926 33702 111978 33754
rect 111990 33702 112042 33754
rect 110788 33464 110840 33516
rect 118056 33303 118108 33312
rect 118056 33269 118065 33303
rect 118065 33269 118099 33303
rect 118099 33269 118108 33303
rect 118056 33260 118108 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 96374 33158 96426 33210
rect 96438 33158 96490 33210
rect 96502 33158 96554 33210
rect 96566 33158 96618 33210
rect 96630 33158 96682 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 81014 32614 81066 32666
rect 81078 32614 81130 32666
rect 81142 32614 81194 32666
rect 81206 32614 81258 32666
rect 81270 32614 81322 32666
rect 111734 32614 111786 32666
rect 111798 32614 111850 32666
rect 111862 32614 111914 32666
rect 111926 32614 111978 32666
rect 111990 32614 112042 32666
rect 108488 32376 108540 32428
rect 118056 32215 118108 32224
rect 118056 32181 118065 32215
rect 118065 32181 118099 32215
rect 118099 32181 118108 32215
rect 118056 32172 118108 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 96374 32070 96426 32122
rect 96438 32070 96490 32122
rect 96502 32070 96554 32122
rect 96566 32070 96618 32122
rect 96630 32070 96682 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 81014 31526 81066 31578
rect 81078 31526 81130 31578
rect 81142 31526 81194 31578
rect 81206 31526 81258 31578
rect 81270 31526 81322 31578
rect 111734 31526 111786 31578
rect 111798 31526 111850 31578
rect 111862 31526 111914 31578
rect 111926 31526 111978 31578
rect 111990 31526 112042 31578
rect 107108 31288 107160 31340
rect 118056 31127 118108 31136
rect 118056 31093 118065 31127
rect 118065 31093 118099 31127
rect 118099 31093 118108 31127
rect 118056 31084 118108 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 96374 30982 96426 31034
rect 96438 30982 96490 31034
rect 96502 30982 96554 31034
rect 96566 30982 96618 31034
rect 96630 30982 96682 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 81014 30438 81066 30490
rect 81078 30438 81130 30490
rect 81142 30438 81194 30490
rect 81206 30438 81258 30490
rect 81270 30438 81322 30490
rect 111734 30438 111786 30490
rect 111798 30438 111850 30490
rect 111862 30438 111914 30490
rect 111926 30438 111978 30490
rect 111990 30438 112042 30490
rect 106004 30200 106056 30252
rect 118056 30107 118108 30116
rect 118056 30073 118065 30107
rect 118065 30073 118099 30107
rect 118099 30073 118108 30107
rect 118056 30064 118108 30073
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 96374 29894 96426 29946
rect 96438 29894 96490 29946
rect 96502 29894 96554 29946
rect 96566 29894 96618 29946
rect 96630 29894 96682 29946
rect 104440 29588 104492 29640
rect 118056 29495 118108 29504
rect 118056 29461 118065 29495
rect 118065 29461 118099 29495
rect 118099 29461 118108 29495
rect 118056 29452 118108 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 81014 29350 81066 29402
rect 81078 29350 81130 29402
rect 81142 29350 81194 29402
rect 81206 29350 81258 29402
rect 81270 29350 81322 29402
rect 111734 29350 111786 29402
rect 111798 29350 111850 29402
rect 111862 29350 111914 29402
rect 111926 29350 111978 29402
rect 111990 29350 112042 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 96374 28806 96426 28858
rect 96438 28806 96490 28858
rect 96502 28806 96554 28858
rect 96566 28806 96618 28858
rect 96630 28806 96682 28858
rect 102416 28500 102468 28552
rect 118056 28407 118108 28416
rect 118056 28373 118065 28407
rect 118065 28373 118099 28407
rect 118099 28373 118108 28407
rect 118056 28364 118108 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 81014 28262 81066 28314
rect 81078 28262 81130 28314
rect 81142 28262 81194 28314
rect 81206 28262 81258 28314
rect 81270 28262 81322 28314
rect 111734 28262 111786 28314
rect 111798 28262 111850 28314
rect 111862 28262 111914 28314
rect 111926 28262 111978 28314
rect 111990 28262 112042 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 96374 27718 96426 27770
rect 96438 27718 96490 27770
rect 96502 27718 96554 27770
rect 96566 27718 96618 27770
rect 96630 27718 96682 27770
rect 100576 27412 100628 27464
rect 118056 27319 118108 27328
rect 118056 27285 118065 27319
rect 118065 27285 118099 27319
rect 118099 27285 118108 27319
rect 118056 27276 118108 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 81014 27174 81066 27226
rect 81078 27174 81130 27226
rect 81142 27174 81194 27226
rect 81206 27174 81258 27226
rect 81270 27174 81322 27226
rect 111734 27174 111786 27226
rect 111798 27174 111850 27226
rect 111862 27174 111914 27226
rect 111926 27174 111978 27226
rect 111990 27174 112042 27226
rect 99840 26936 99892 26988
rect 118056 26775 118108 26784
rect 118056 26741 118065 26775
rect 118065 26741 118099 26775
rect 118099 26741 118108 26775
rect 118056 26732 118108 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 96374 26630 96426 26682
rect 96438 26630 96490 26682
rect 96502 26630 96554 26682
rect 96566 26630 96618 26682
rect 96630 26630 96682 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 81014 26086 81066 26138
rect 81078 26086 81130 26138
rect 81142 26086 81194 26138
rect 81206 26086 81258 26138
rect 81270 26086 81322 26138
rect 111734 26086 111786 26138
rect 111798 26086 111850 26138
rect 111862 26086 111914 26138
rect 111926 26086 111978 26138
rect 111990 26086 112042 26138
rect 98092 25848 98144 25900
rect 118056 25687 118108 25696
rect 118056 25653 118065 25687
rect 118065 25653 118099 25687
rect 118099 25653 118108 25687
rect 118056 25644 118108 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 96374 25542 96426 25594
rect 96438 25542 96490 25594
rect 96502 25542 96554 25594
rect 96566 25542 96618 25594
rect 96630 25542 96682 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 81014 24998 81066 25050
rect 81078 24998 81130 25050
rect 81142 24998 81194 25050
rect 81206 24998 81258 25050
rect 81270 24998 81322 25050
rect 111734 24998 111786 25050
rect 111798 24998 111850 25050
rect 111862 24998 111914 25050
rect 111926 24998 111978 25050
rect 111990 24998 112042 25050
rect 96896 24760 96948 24812
rect 118056 24599 118108 24608
rect 118056 24565 118065 24599
rect 118065 24565 118099 24599
rect 118099 24565 118108 24599
rect 118056 24556 118108 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 96374 24454 96426 24506
rect 96438 24454 96490 24506
rect 96502 24454 96554 24506
rect 96566 24454 96618 24506
rect 96630 24454 96682 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 81014 23910 81066 23962
rect 81078 23910 81130 23962
rect 81142 23910 81194 23962
rect 81206 23910 81258 23962
rect 81270 23910 81322 23962
rect 111734 23910 111786 23962
rect 111798 23910 111850 23962
rect 111862 23910 111914 23962
rect 111926 23910 111978 23962
rect 111990 23910 112042 23962
rect 95976 23672 96028 23724
rect 118056 23579 118108 23588
rect 118056 23545 118065 23579
rect 118065 23545 118099 23579
rect 118099 23545 118108 23579
rect 118056 23536 118108 23545
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 96374 23366 96426 23418
rect 96438 23366 96490 23418
rect 96502 23366 96554 23418
rect 96566 23366 96618 23418
rect 96630 23366 96682 23418
rect 93124 23060 93176 23112
rect 118056 22967 118108 22976
rect 118056 22933 118065 22967
rect 118065 22933 118099 22967
rect 118099 22933 118108 22967
rect 118056 22924 118108 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 81014 22822 81066 22874
rect 81078 22822 81130 22874
rect 81142 22822 81194 22874
rect 81206 22822 81258 22874
rect 81270 22822 81322 22874
rect 111734 22822 111786 22874
rect 111798 22822 111850 22874
rect 111862 22822 111914 22874
rect 111926 22822 111978 22874
rect 111990 22822 112042 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 96374 22278 96426 22330
rect 96438 22278 96490 22330
rect 96502 22278 96554 22330
rect 96566 22278 96618 22330
rect 96630 22278 96682 22330
rect 92388 21836 92440 21888
rect 118056 21879 118108 21888
rect 118056 21845 118065 21879
rect 118065 21845 118099 21879
rect 118099 21845 118108 21879
rect 118056 21836 118108 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 81014 21734 81066 21786
rect 81078 21734 81130 21786
rect 81142 21734 81194 21786
rect 81206 21734 81258 21786
rect 81270 21734 81322 21786
rect 111734 21734 111786 21786
rect 111798 21734 111850 21786
rect 111862 21734 111914 21786
rect 111926 21734 111978 21786
rect 111990 21734 112042 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 96374 21190 96426 21242
rect 96438 21190 96490 21242
rect 96502 21190 96554 21242
rect 96566 21190 96618 21242
rect 96630 21190 96682 21242
rect 91008 20884 91060 20936
rect 118056 20791 118108 20800
rect 118056 20757 118065 20791
rect 118065 20757 118099 20791
rect 118099 20757 118108 20791
rect 118056 20748 118108 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 81014 20646 81066 20698
rect 81078 20646 81130 20698
rect 81142 20646 81194 20698
rect 81206 20646 81258 20698
rect 81270 20646 81322 20698
rect 111734 20646 111786 20698
rect 111798 20646 111850 20698
rect 111862 20646 111914 20698
rect 111926 20646 111978 20698
rect 111990 20646 112042 20698
rect 89444 20408 89496 20460
rect 118056 20247 118108 20256
rect 118056 20213 118065 20247
rect 118065 20213 118099 20247
rect 118099 20213 118108 20247
rect 118056 20204 118108 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 96374 20102 96426 20154
rect 96438 20102 96490 20154
rect 96502 20102 96554 20154
rect 96566 20102 96618 20154
rect 96630 20102 96682 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 81014 19558 81066 19610
rect 81078 19558 81130 19610
rect 81142 19558 81194 19610
rect 81206 19558 81258 19610
rect 81270 19558 81322 19610
rect 111734 19558 111786 19610
rect 111798 19558 111850 19610
rect 111862 19558 111914 19610
rect 111926 19558 111978 19610
rect 111990 19558 112042 19610
rect 117412 19116 117464 19168
rect 118056 19159 118108 19168
rect 118056 19125 118065 19159
rect 118065 19125 118099 19159
rect 118099 19125 118108 19159
rect 118056 19116 118108 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 96374 19014 96426 19066
rect 96438 19014 96490 19066
rect 96502 19014 96554 19066
rect 96566 19014 96618 19066
rect 96630 19014 96682 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 81014 18470 81066 18522
rect 81078 18470 81130 18522
rect 81142 18470 81194 18522
rect 81206 18470 81258 18522
rect 81270 18470 81322 18522
rect 111734 18470 111786 18522
rect 111798 18470 111850 18522
rect 111862 18470 111914 18522
rect 111926 18470 111978 18522
rect 111990 18470 112042 18522
rect 86684 18028 86736 18080
rect 118056 18071 118108 18080
rect 118056 18037 118065 18071
rect 118065 18037 118099 18071
rect 118099 18037 118108 18071
rect 118056 18028 118108 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 96374 17926 96426 17978
rect 96438 17926 96490 17978
rect 96502 17926 96554 17978
rect 96566 17926 96618 17978
rect 96630 17926 96682 17978
rect 85212 17620 85264 17672
rect 118056 17527 118108 17536
rect 118056 17493 118065 17527
rect 118065 17493 118099 17527
rect 118099 17493 118108 17527
rect 118056 17484 118108 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 81014 17382 81066 17434
rect 81078 17382 81130 17434
rect 81142 17382 81194 17434
rect 81206 17382 81258 17434
rect 81270 17382 81322 17434
rect 111734 17382 111786 17434
rect 111798 17382 111850 17434
rect 111862 17382 111914 17434
rect 111926 17382 111978 17434
rect 111990 17382 112042 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 96374 16838 96426 16890
rect 96438 16838 96490 16890
rect 96502 16838 96554 16890
rect 96566 16838 96618 16890
rect 96630 16838 96682 16890
rect 117504 16439 117556 16448
rect 117504 16405 117513 16439
rect 117513 16405 117547 16439
rect 117547 16405 117556 16439
rect 117504 16396 117556 16405
rect 118056 16439 118108 16448
rect 118056 16405 118065 16439
rect 118065 16405 118099 16439
rect 118099 16405 118108 16439
rect 118056 16396 118108 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 81014 16294 81066 16346
rect 81078 16294 81130 16346
rect 81142 16294 81194 16346
rect 81206 16294 81258 16346
rect 81270 16294 81322 16346
rect 111734 16294 111786 16346
rect 111798 16294 111850 16346
rect 111862 16294 111914 16346
rect 111926 16294 111978 16346
rect 111990 16294 112042 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 96374 15750 96426 15802
rect 96438 15750 96490 15802
rect 96502 15750 96554 15802
rect 96566 15750 96618 15802
rect 96630 15750 96682 15802
rect 82820 15444 82872 15496
rect 118056 15351 118108 15360
rect 118056 15317 118065 15351
rect 118065 15317 118099 15351
rect 118099 15317 118108 15351
rect 118056 15308 118108 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 81014 15206 81066 15258
rect 81078 15206 81130 15258
rect 81142 15206 81194 15258
rect 81206 15206 81258 15258
rect 81270 15206 81322 15258
rect 111734 15206 111786 15258
rect 111798 15206 111850 15258
rect 111862 15206 111914 15258
rect 111926 15206 111978 15258
rect 111990 15206 112042 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 96374 14662 96426 14714
rect 96438 14662 96490 14714
rect 96502 14662 96554 14714
rect 96566 14662 96618 14714
rect 96630 14662 96682 14714
rect 81716 14356 81768 14408
rect 118056 14263 118108 14272
rect 118056 14229 118065 14263
rect 118065 14229 118099 14263
rect 118099 14229 118108 14263
rect 118056 14220 118108 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 81014 14118 81066 14170
rect 81078 14118 81130 14170
rect 81142 14118 81194 14170
rect 81206 14118 81258 14170
rect 81270 14118 81322 14170
rect 111734 14118 111786 14170
rect 111798 14118 111850 14170
rect 111862 14118 111914 14170
rect 111926 14118 111978 14170
rect 111990 14118 112042 14170
rect 79600 13880 79652 13932
rect 118056 13719 118108 13728
rect 118056 13685 118065 13719
rect 118065 13685 118099 13719
rect 118099 13685 118108 13719
rect 118056 13676 118108 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 96374 13574 96426 13626
rect 96438 13574 96490 13626
rect 96502 13574 96554 13626
rect 96566 13574 96618 13626
rect 96630 13574 96682 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 81014 13030 81066 13082
rect 81078 13030 81130 13082
rect 81142 13030 81194 13082
rect 81206 13030 81258 13082
rect 81270 13030 81322 13082
rect 111734 13030 111786 13082
rect 111798 13030 111850 13082
rect 111862 13030 111914 13082
rect 111926 13030 111978 13082
rect 111990 13030 112042 13082
rect 89444 12971 89496 12980
rect 89444 12937 89453 12971
rect 89453 12937 89487 12971
rect 89487 12937 89496 12971
rect 89444 12928 89496 12937
rect 78680 12792 78732 12844
rect 88800 12792 88852 12844
rect 118056 12631 118108 12640
rect 118056 12597 118065 12631
rect 118065 12597 118099 12631
rect 118099 12597 118108 12631
rect 118056 12588 118108 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 96374 12486 96426 12538
rect 96438 12486 96490 12538
rect 96502 12486 96554 12538
rect 96566 12486 96618 12538
rect 96630 12486 96682 12538
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 81014 11942 81066 11994
rect 81078 11942 81130 11994
rect 81142 11942 81194 11994
rect 81206 11942 81258 11994
rect 81270 11942 81322 11994
rect 111734 11942 111786 11994
rect 111798 11942 111850 11994
rect 111862 11942 111914 11994
rect 111926 11942 111978 11994
rect 111990 11942 112042 11994
rect 76656 11500 76708 11552
rect 118056 11611 118108 11620
rect 118056 11577 118065 11611
rect 118065 11577 118099 11611
rect 118099 11577 118108 11611
rect 118056 11568 118108 11577
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 96374 11398 96426 11450
rect 96438 11398 96490 11450
rect 96502 11398 96554 11450
rect 96566 11398 96618 11450
rect 96630 11398 96682 11450
rect 118056 11271 118108 11280
rect 118056 11237 118065 11271
rect 118065 11237 118099 11271
rect 118099 11237 118108 11271
rect 118056 11228 118108 11237
rect 76104 11092 76156 11144
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 81014 10854 81066 10906
rect 81078 10854 81130 10906
rect 81142 10854 81194 10906
rect 81206 10854 81258 10906
rect 81270 10854 81322 10906
rect 111734 10854 111786 10906
rect 111798 10854 111850 10906
rect 111862 10854 111914 10906
rect 111926 10854 111978 10906
rect 111990 10854 112042 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 96374 10310 96426 10362
rect 96438 10310 96490 10362
rect 96502 10310 96554 10362
rect 96566 10310 96618 10362
rect 96630 10310 96682 10362
rect 76104 10251 76156 10260
rect 76104 10217 76113 10251
rect 76113 10217 76147 10251
rect 76147 10217 76156 10251
rect 76104 10208 76156 10217
rect 74632 10004 74684 10056
rect 117780 9979 117832 9988
rect 117780 9945 117789 9979
rect 117789 9945 117823 9979
rect 117823 9945 117832 9979
rect 117780 9936 117832 9945
rect 107660 9868 107712 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 81014 9766 81066 9818
rect 81078 9766 81130 9818
rect 81142 9766 81194 9818
rect 81206 9766 81258 9818
rect 81270 9766 81322 9818
rect 111734 9766 111786 9818
rect 111798 9766 111850 9818
rect 111862 9766 111914 9818
rect 111926 9766 111978 9818
rect 111990 9766 112042 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 96374 9222 96426 9274
rect 96438 9222 96490 9274
rect 96502 9222 96554 9274
rect 96566 9222 96618 9274
rect 96630 9222 96682 9274
rect 117780 8891 117832 8900
rect 117780 8857 117789 8891
rect 117789 8857 117823 8891
rect 117823 8857 117832 8891
rect 117780 8848 117832 8857
rect 73528 8780 73580 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 81014 8678 81066 8730
rect 81078 8678 81130 8730
rect 81142 8678 81194 8730
rect 81206 8678 81258 8730
rect 81270 8678 81322 8730
rect 111734 8678 111786 8730
rect 111798 8678 111850 8730
rect 111862 8678 111914 8730
rect 111926 8678 111978 8730
rect 111990 8678 112042 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 96374 8134 96426 8186
rect 96438 8134 96490 8186
rect 96502 8134 96554 8186
rect 96566 8134 96618 8186
rect 96630 8134 96682 8186
rect 117780 7803 117832 7812
rect 117780 7769 117789 7803
rect 117789 7769 117823 7803
rect 117823 7769 117832 7803
rect 117780 7760 117832 7769
rect 71688 7692 71740 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 81014 7590 81066 7642
rect 81078 7590 81130 7642
rect 81142 7590 81194 7642
rect 81206 7590 81258 7642
rect 81270 7590 81322 7642
rect 111734 7590 111786 7642
rect 111798 7590 111850 7642
rect 111862 7590 111914 7642
rect 111926 7590 111978 7642
rect 111990 7590 112042 7642
rect 117780 7395 117832 7404
rect 117780 7361 117789 7395
rect 117789 7361 117823 7395
rect 117823 7361 117832 7395
rect 117780 7352 117832 7361
rect 116860 7148 116912 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 96374 7046 96426 7098
rect 96438 7046 96490 7098
rect 96502 7046 96554 7098
rect 96566 7046 96618 7098
rect 96630 7046 96682 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 81014 6502 81066 6554
rect 81078 6502 81130 6554
rect 81142 6502 81194 6554
rect 81206 6502 81258 6554
rect 81270 6502 81322 6554
rect 111734 6502 111786 6554
rect 111798 6502 111850 6554
rect 111862 6502 111914 6554
rect 111926 6502 111978 6554
rect 111990 6502 112042 6554
rect 91008 6443 91060 6452
rect 91008 6409 91017 6443
rect 91017 6409 91051 6443
rect 91051 6409 91060 6443
rect 91008 6400 91060 6409
rect 88340 6264 88392 6316
rect 90824 6307 90876 6316
rect 90824 6273 90833 6307
rect 90833 6273 90867 6307
rect 90867 6273 90876 6307
rect 90824 6264 90876 6273
rect 117412 6264 117464 6316
rect 117780 6307 117832 6316
rect 117780 6273 117789 6307
rect 117789 6273 117823 6307
rect 117823 6273 117832 6307
rect 117780 6264 117832 6273
rect 117504 6060 117556 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 96374 5958 96426 6010
rect 96438 5958 96490 6010
rect 96502 5958 96554 6010
rect 96566 5958 96618 6010
rect 96630 5958 96682 6010
rect 117688 5652 117740 5704
rect 116308 5516 116360 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 81014 5414 81066 5466
rect 81078 5414 81130 5466
rect 81142 5414 81194 5466
rect 81206 5414 81258 5466
rect 81270 5414 81322 5466
rect 111734 5414 111786 5466
rect 111798 5414 111850 5466
rect 111862 5414 111914 5466
rect 111926 5414 111978 5466
rect 111990 5414 112042 5466
rect 117780 5219 117832 5228
rect 117780 5185 117789 5219
rect 117789 5185 117823 5219
rect 117823 5185 117832 5219
rect 117780 5176 117832 5185
rect 117872 5015 117924 5024
rect 117872 4981 117881 5015
rect 117881 4981 117915 5015
rect 117915 4981 117924 5015
rect 117872 4972 117924 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 96374 4870 96426 4922
rect 96438 4870 96490 4922
rect 96502 4870 96554 4922
rect 96566 4870 96618 4922
rect 96630 4870 96682 4922
rect 117596 4768 117648 4820
rect 116216 4607 116268 4616
rect 116216 4573 116225 4607
rect 116225 4573 116259 4607
rect 116259 4573 116268 4607
rect 116216 4564 116268 4573
rect 117780 4539 117832 4548
rect 117780 4505 117789 4539
rect 117789 4505 117823 4539
rect 117823 4505 117832 4539
rect 117780 4496 117832 4505
rect 97540 4428 97592 4480
rect 104164 4428 104216 4480
rect 115296 4428 115348 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 81014 4326 81066 4378
rect 81078 4326 81130 4378
rect 81142 4326 81194 4378
rect 81206 4326 81258 4378
rect 81270 4326 81322 4378
rect 111734 4326 111786 4378
rect 111798 4326 111850 4378
rect 111862 4326 111914 4378
rect 111926 4326 111978 4378
rect 111990 4326 112042 4378
rect 58256 4224 58308 4276
rect 97540 4224 97592 4276
rect 98000 4224 98052 4276
rect 100392 4224 100444 4276
rect 104164 4224 104216 4276
rect 116124 4224 116176 4276
rect 25688 4156 25740 4208
rect 85028 4156 85080 4208
rect 67364 4088 67416 4140
rect 97908 4088 97960 4140
rect 100852 4131 100904 4140
rect 100852 4097 100861 4131
rect 100861 4097 100895 4131
rect 100895 4097 100904 4131
rect 114744 4156 114796 4208
rect 117504 4224 117556 4276
rect 117228 4156 117280 4208
rect 100852 4088 100904 4097
rect 63132 4020 63184 4072
rect 113364 4020 113416 4072
rect 114836 4088 114888 4140
rect 115848 4131 115900 4140
rect 115848 4097 115857 4131
rect 115857 4097 115891 4131
rect 115891 4097 115900 4131
rect 115848 4088 115900 4097
rect 116584 4131 116636 4140
rect 116584 4097 116593 4131
rect 116593 4097 116627 4131
rect 116627 4097 116636 4131
rect 116584 4088 116636 4097
rect 116676 4088 116728 4140
rect 118148 4088 118200 4140
rect 117872 4020 117924 4072
rect 68836 3952 68888 4004
rect 64972 3884 65024 3936
rect 111524 3884 111576 3936
rect 111708 3952 111760 4004
rect 114744 3884 114796 3936
rect 115388 3884 115440 3936
rect 116676 3884 116728 3936
rect 118424 3884 118476 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 96374 3782 96426 3834
rect 96438 3782 96490 3834
rect 96502 3782 96554 3834
rect 96566 3782 96618 3834
rect 96630 3782 96682 3834
rect 61660 3680 61712 3732
rect 113272 3680 113324 3732
rect 113364 3680 113416 3732
rect 57152 3612 57204 3664
rect 98644 3612 98696 3664
rect 98920 3612 98972 3664
rect 106004 3655 106056 3664
rect 45192 3544 45244 3596
rect 98736 3544 98788 3596
rect 63132 3519 63184 3528
rect 63132 3485 63141 3519
rect 63141 3485 63175 3519
rect 63175 3485 63184 3519
rect 63132 3476 63184 3485
rect 68284 3476 68336 3528
rect 68836 3519 68888 3528
rect 68836 3485 68845 3519
rect 68845 3485 68879 3519
rect 68879 3485 68888 3519
rect 68836 3476 68888 3485
rect 76288 3476 76340 3528
rect 81992 3476 82044 3528
rect 83464 3476 83516 3528
rect 84844 3476 84896 3528
rect 86316 3476 86368 3528
rect 87696 3476 87748 3528
rect 92020 3476 92072 3528
rect 92204 3519 92256 3528
rect 92204 3485 92213 3519
rect 92213 3485 92247 3519
rect 92247 3485 92256 3519
rect 92204 3476 92256 3485
rect 96160 3476 96212 3528
rect 97724 3476 97776 3528
rect 98644 3476 98696 3528
rect 106004 3621 106013 3655
rect 106013 3621 106047 3655
rect 106047 3621 106056 3655
rect 106004 3612 106056 3621
rect 106096 3612 106148 3664
rect 107660 3612 107712 3664
rect 114928 3655 114980 3664
rect 114928 3621 114937 3655
rect 114937 3621 114971 3655
rect 114971 3621 114980 3655
rect 114928 3612 114980 3621
rect 114008 3544 114060 3596
rect 114100 3544 114152 3596
rect 99288 3476 99340 3528
rect 100300 3476 100352 3528
rect 105820 3519 105872 3528
rect 105820 3485 105829 3519
rect 105829 3485 105863 3519
rect 105863 3485 105872 3519
rect 105820 3476 105872 3485
rect 106280 3476 106332 3528
rect 112260 3519 112312 3528
rect 112260 3485 112269 3519
rect 112269 3485 112303 3519
rect 112303 3485 112312 3519
rect 112260 3476 112312 3485
rect 115204 3544 115256 3596
rect 116400 3587 116452 3596
rect 116400 3553 116409 3587
rect 116409 3553 116443 3587
rect 116443 3553 116452 3587
rect 116400 3544 116452 3553
rect 116124 3519 116176 3528
rect 65524 3408 65576 3460
rect 76196 3408 76248 3460
rect 88892 3408 88944 3460
rect 97632 3408 97684 3460
rect 99104 3408 99156 3460
rect 99564 3408 99616 3460
rect 63592 3340 63644 3392
rect 69112 3340 69164 3392
rect 76472 3340 76524 3392
rect 83096 3340 83148 3392
rect 83556 3383 83608 3392
rect 83556 3349 83565 3383
rect 83565 3349 83599 3383
rect 83599 3349 83608 3383
rect 83556 3340 83608 3349
rect 84936 3383 84988 3392
rect 84936 3349 84945 3383
rect 84945 3349 84979 3383
rect 84979 3349 84988 3383
rect 84936 3340 84988 3349
rect 86408 3383 86460 3392
rect 86408 3349 86417 3383
rect 86417 3349 86451 3383
rect 86451 3349 86460 3383
rect 86408 3340 86460 3349
rect 87788 3383 87840 3392
rect 87788 3349 87797 3383
rect 87797 3349 87831 3383
rect 87831 3349 87840 3383
rect 87788 3340 87840 3349
rect 91560 3383 91612 3392
rect 91560 3349 91569 3383
rect 91569 3349 91603 3383
rect 91603 3349 91612 3383
rect 91560 3340 91612 3349
rect 92388 3383 92440 3392
rect 92388 3349 92397 3383
rect 92397 3349 92431 3383
rect 92431 3349 92440 3383
rect 92388 3340 92440 3349
rect 96988 3340 97040 3392
rect 98092 3383 98144 3392
rect 98092 3349 98101 3383
rect 98101 3349 98135 3383
rect 98135 3349 98144 3383
rect 98092 3340 98144 3349
rect 99840 3383 99892 3392
rect 99840 3349 99849 3383
rect 99849 3349 99883 3383
rect 99883 3349 99892 3383
rect 99840 3340 99892 3349
rect 100576 3383 100628 3392
rect 100576 3349 100585 3383
rect 100585 3349 100619 3383
rect 100619 3349 100628 3383
rect 100576 3340 100628 3349
rect 100760 3340 100812 3392
rect 106004 3340 106056 3392
rect 106096 3340 106148 3392
rect 112076 3383 112128 3392
rect 112076 3349 112085 3383
rect 112085 3349 112119 3383
rect 112119 3349 112128 3383
rect 112076 3340 112128 3349
rect 114928 3408 114980 3460
rect 116124 3485 116133 3519
rect 116133 3485 116167 3519
rect 116167 3485 116176 3519
rect 116124 3476 116176 3485
rect 116308 3476 116360 3528
rect 116860 3408 116912 3460
rect 117136 3408 117188 3460
rect 117964 3340 118016 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 81014 3238 81066 3290
rect 81078 3238 81130 3290
rect 81142 3238 81194 3290
rect 81206 3238 81258 3290
rect 81270 3238 81322 3290
rect 111734 3238 111786 3290
rect 111798 3238 111850 3290
rect 111862 3238 111914 3290
rect 111926 3238 111978 3290
rect 111990 3238 112042 3290
rect 17040 3136 17092 3188
rect 65524 3136 65576 3188
rect 76656 3179 76708 3188
rect 54852 3000 54904 3052
rect 59176 3000 59228 3052
rect 59544 3000 59596 3052
rect 61384 3068 61436 3120
rect 76656 3145 76665 3179
rect 76665 3145 76699 3179
rect 76699 3145 76708 3179
rect 76656 3136 76708 3145
rect 78680 3179 78732 3188
rect 78680 3145 78689 3179
rect 78689 3145 78723 3179
rect 78723 3145 78732 3179
rect 78680 3136 78732 3145
rect 79600 3179 79652 3188
rect 79600 3145 79609 3179
rect 79609 3145 79643 3179
rect 79643 3145 79652 3179
rect 79600 3136 79652 3145
rect 81716 3179 81768 3188
rect 81716 3145 81725 3179
rect 81725 3145 81759 3179
rect 81759 3145 81768 3179
rect 81716 3136 81768 3145
rect 82820 3179 82872 3188
rect 82820 3145 82829 3179
rect 82829 3145 82863 3179
rect 82863 3145 82872 3179
rect 82820 3136 82872 3145
rect 85212 3179 85264 3188
rect 85212 3145 85221 3179
rect 85221 3145 85255 3179
rect 85255 3145 85264 3179
rect 85212 3136 85264 3145
rect 86684 3179 86736 3188
rect 86684 3145 86693 3179
rect 86693 3145 86727 3179
rect 86727 3145 86736 3179
rect 86684 3136 86736 3145
rect 61016 3000 61068 3052
rect 61660 3043 61712 3052
rect 61660 3009 61669 3043
rect 61669 3009 61703 3043
rect 61703 3009 61712 3043
rect 61660 3000 61712 3009
rect 63592 3043 63644 3052
rect 63592 3009 63601 3043
rect 63601 3009 63635 3043
rect 63635 3009 63644 3043
rect 63592 3000 63644 3009
rect 64880 3043 64932 3052
rect 64880 3009 64889 3043
rect 64889 3009 64923 3043
rect 64923 3009 64932 3043
rect 64880 3000 64932 3009
rect 51908 2864 51960 2916
rect 56692 2864 56744 2916
rect 64420 2932 64472 2984
rect 64972 2932 65024 2984
rect 65524 2975 65576 2984
rect 65524 2941 65533 2975
rect 65533 2941 65567 2975
rect 65567 2941 65576 2975
rect 70124 3068 70176 3120
rect 92572 3136 92624 3188
rect 93952 3136 94004 3188
rect 95976 3179 96028 3188
rect 95976 3145 95985 3179
rect 95985 3145 96019 3179
rect 96019 3145 96028 3179
rect 95976 3136 96028 3145
rect 96896 3136 96948 3188
rect 99288 3136 99340 3188
rect 102416 3179 102468 3188
rect 102416 3145 102425 3179
rect 102425 3145 102459 3179
rect 102459 3145 102468 3179
rect 102416 3136 102468 3145
rect 104440 3179 104492 3188
rect 104440 3145 104449 3179
rect 104449 3145 104483 3179
rect 104483 3145 104492 3179
rect 104440 3136 104492 3145
rect 106096 3179 106148 3188
rect 106096 3145 106105 3179
rect 106105 3145 106139 3179
rect 106139 3145 106148 3179
rect 106096 3136 106148 3145
rect 107108 3136 107160 3188
rect 108488 3179 108540 3188
rect 108488 3145 108497 3179
rect 108497 3145 108531 3179
rect 108531 3145 108540 3179
rect 108488 3136 108540 3145
rect 110788 3179 110840 3188
rect 66720 3000 66772 3052
rect 67364 3043 67416 3052
rect 67364 3009 67373 3043
rect 67373 3009 67407 3043
rect 67407 3009 67416 3043
rect 67364 3000 67416 3009
rect 69112 3043 69164 3052
rect 69112 3009 69121 3043
rect 69121 3009 69155 3043
rect 69155 3009 69164 3043
rect 69112 3000 69164 3009
rect 65524 2932 65576 2941
rect 56508 2796 56560 2848
rect 66168 2864 66220 2916
rect 61108 2796 61160 2848
rect 62120 2796 62172 2848
rect 63500 2796 63552 2848
rect 64972 2796 65024 2848
rect 66352 2796 66404 2848
rect 67732 2796 67784 2848
rect 69204 2796 69256 2848
rect 69572 2796 69624 2848
rect 88892 3111 88944 3120
rect 88892 3077 88901 3111
rect 88901 3077 88935 3111
rect 88935 3077 88944 3111
rect 88892 3068 88944 3077
rect 71688 3043 71740 3052
rect 71688 3009 71697 3043
rect 71697 3009 71731 3043
rect 71731 3009 71740 3043
rect 71688 3000 71740 3009
rect 73528 3043 73580 3052
rect 73528 3009 73537 3043
rect 73537 3009 73571 3043
rect 73571 3009 73580 3043
rect 73528 3000 73580 3009
rect 74908 3000 74960 3052
rect 76564 3043 76616 3052
rect 76564 3009 76573 3043
rect 76573 3009 76607 3043
rect 76607 3009 76616 3043
rect 76564 3000 76616 3009
rect 77760 3000 77812 3052
rect 78588 3043 78640 3052
rect 78588 3009 78597 3043
rect 78597 3009 78631 3043
rect 78631 3009 78640 3043
rect 78588 3000 78640 3009
rect 79508 3043 79560 3052
rect 79508 3009 79517 3043
rect 79517 3009 79551 3043
rect 79551 3009 79560 3043
rect 79508 3000 79560 3009
rect 80612 3000 80664 3052
rect 81624 3043 81676 3052
rect 81624 3009 81633 3043
rect 81633 3009 81667 3043
rect 81667 3009 81676 3043
rect 81624 3000 81676 3009
rect 82544 3043 82596 3052
rect 82544 3009 82553 3043
rect 82553 3009 82587 3043
rect 82587 3009 82596 3043
rect 82544 3000 82596 3009
rect 83740 3043 83792 3052
rect 83740 3009 83749 3043
rect 83749 3009 83783 3043
rect 83783 3009 83792 3043
rect 83740 3000 83792 3009
rect 85120 3043 85172 3052
rect 85120 3009 85129 3043
rect 85129 3009 85163 3043
rect 85163 3009 85172 3043
rect 85120 3000 85172 3009
rect 86592 3043 86644 3052
rect 86592 3009 86601 3043
rect 86601 3009 86635 3043
rect 86635 3009 86644 3043
rect 86592 3000 86644 3009
rect 70124 2864 70176 2916
rect 99656 3068 99708 3120
rect 100576 3068 100628 3120
rect 110788 3145 110797 3179
rect 110797 3145 110831 3179
rect 110831 3145 110840 3179
rect 110788 3136 110840 3145
rect 112168 3136 112220 3188
rect 114008 3136 114060 3188
rect 89168 3000 89220 3052
rect 90640 3000 90692 3052
rect 91468 3000 91520 3052
rect 92572 3043 92624 3052
rect 92572 3009 92581 3043
rect 92581 3009 92615 3043
rect 92615 3009 92624 3043
rect 92572 3000 92624 3009
rect 92664 3000 92716 3052
rect 89444 2932 89496 2984
rect 92296 2932 92348 2984
rect 92848 2932 92900 2984
rect 94872 3000 94924 3052
rect 95792 3043 95844 3052
rect 95792 3009 95801 3043
rect 95801 3009 95835 3043
rect 95835 3009 95844 3043
rect 95792 3000 95844 3009
rect 96252 3000 96304 3052
rect 97632 3043 97684 3052
rect 97632 3009 97641 3043
rect 97641 3009 97675 3043
rect 97675 3009 97684 3043
rect 97632 3000 97684 3009
rect 98644 3000 98696 3052
rect 99472 3043 99524 3052
rect 99472 3009 99481 3043
rect 99481 3009 99515 3043
rect 99515 3009 99524 3043
rect 99472 3000 99524 3009
rect 101220 3043 101272 3052
rect 99564 2932 99616 2984
rect 99748 2975 99800 2984
rect 99748 2941 99757 2975
rect 99757 2941 99791 2975
rect 99791 2941 99800 2975
rect 99748 2932 99800 2941
rect 101220 3009 101229 3043
rect 101229 3009 101263 3043
rect 101263 3009 101272 3043
rect 101220 3000 101272 3009
rect 102140 3000 102192 3052
rect 104256 3043 104308 3052
rect 100760 2932 100812 2984
rect 102048 2932 102100 2984
rect 104256 3009 104265 3043
rect 104265 3009 104299 3043
rect 104299 3009 104308 3043
rect 104256 3000 104308 3009
rect 104900 3000 104952 3052
rect 105268 3000 105320 3052
rect 106188 2975 106240 2984
rect 106188 2941 106197 2975
rect 106197 2941 106231 2975
rect 106231 2941 106240 2975
rect 106188 2932 106240 2941
rect 70584 2796 70636 2848
rect 72056 2796 72108 2848
rect 73528 2796 73580 2848
rect 75000 2839 75052 2848
rect 75000 2805 75009 2839
rect 75009 2805 75043 2839
rect 75043 2805 75052 2839
rect 75000 2796 75052 2805
rect 77668 2796 77720 2848
rect 81532 2796 81584 2848
rect 86868 2796 86920 2848
rect 89260 2796 89312 2848
rect 90548 2796 90600 2848
rect 91468 2839 91520 2848
rect 91468 2805 91477 2839
rect 91477 2805 91511 2839
rect 91511 2805 91520 2839
rect 91468 2796 91520 2805
rect 92940 2796 92992 2848
rect 95516 2796 95568 2848
rect 97908 2796 97960 2848
rect 98460 2839 98512 2848
rect 98460 2805 98469 2839
rect 98469 2805 98503 2839
rect 98503 2805 98512 2839
rect 98460 2796 98512 2805
rect 98644 2796 98696 2848
rect 102324 2796 102376 2848
rect 102968 2839 103020 2848
rect 102968 2805 102977 2839
rect 102977 2805 103011 2839
rect 103011 2805 103020 2839
rect 102968 2796 103020 2805
rect 105176 2796 105228 2848
rect 107752 3000 107804 3052
rect 108304 3043 108356 3052
rect 108304 3009 108313 3043
rect 108313 3009 108347 3043
rect 108347 3009 108356 3043
rect 108304 3000 108356 3009
rect 109040 3000 109092 3052
rect 110512 3000 110564 3052
rect 110696 3000 110748 3052
rect 112536 3043 112588 3052
rect 109960 2975 110012 2984
rect 109960 2941 109969 2975
rect 109969 2941 110003 2975
rect 110003 2941 110012 2975
rect 109960 2932 110012 2941
rect 107660 2839 107712 2848
rect 107660 2805 107669 2839
rect 107669 2805 107703 2839
rect 107703 2805 107712 2839
rect 107660 2796 107712 2805
rect 112536 3009 112545 3043
rect 112545 3009 112579 3043
rect 112579 3009 112588 3043
rect 112536 3000 112588 3009
rect 113456 3000 113508 3052
rect 115296 2932 115348 2984
rect 116216 3136 116268 3188
rect 116308 3000 116360 3052
rect 117780 3043 117832 3052
rect 117780 3009 117789 3043
rect 117789 3009 117823 3043
rect 117823 3009 117832 3043
rect 117780 3000 117832 3009
rect 115480 2932 115532 2984
rect 116400 2975 116452 2984
rect 116400 2941 116409 2975
rect 116409 2941 116443 2975
rect 116443 2941 116452 2975
rect 116400 2932 116452 2941
rect 117412 2864 117464 2916
rect 112628 2839 112680 2848
rect 112628 2805 112637 2839
rect 112637 2805 112671 2839
rect 112671 2805 112680 2839
rect 112628 2796 112680 2805
rect 113548 2839 113600 2848
rect 113548 2805 113557 2839
rect 113557 2805 113591 2839
rect 113591 2805 113600 2839
rect 113548 2796 113600 2805
rect 113640 2796 113692 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 96374 2694 96426 2746
rect 96438 2694 96490 2746
rect 96502 2694 96554 2746
rect 96566 2694 96618 2746
rect 96630 2694 96682 2746
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 17040 2567 17092 2576
rect 17040 2533 17049 2567
rect 17049 2533 17083 2567
rect 17083 2533 17092 2567
rect 17040 2524 17092 2533
rect 55864 2524 55916 2576
rect 35900 2456 35952 2508
rect 35992 2456 36044 2508
rect 45376 2456 45428 2508
rect 45468 2456 45520 2508
rect 55772 2456 55824 2508
rect 56140 2635 56192 2644
rect 56140 2601 56149 2635
rect 56149 2601 56183 2635
rect 56183 2601 56192 2635
rect 56140 2592 56192 2601
rect 57152 2635 57204 2644
rect 57152 2601 57161 2635
rect 57161 2601 57195 2635
rect 57195 2601 57204 2635
rect 57152 2592 57204 2601
rect 58256 2635 58308 2644
rect 58256 2601 58265 2635
rect 58265 2601 58299 2635
rect 58299 2601 58308 2635
rect 58256 2592 58308 2601
rect 58440 2592 58492 2644
rect 64144 2635 64196 2644
rect 56048 2524 56100 2576
rect 64144 2601 64153 2635
rect 64153 2601 64187 2635
rect 64187 2601 64196 2635
rect 64144 2592 64196 2601
rect 64880 2592 64932 2644
rect 65156 2635 65208 2644
rect 65156 2601 65165 2635
rect 65165 2601 65199 2635
rect 65199 2601 65208 2635
rect 65156 2592 65208 2601
rect 65248 2592 65300 2644
rect 74632 2635 74684 2644
rect 74632 2601 74641 2635
rect 74641 2601 74675 2635
rect 74675 2601 74684 2635
rect 74632 2592 74684 2601
rect 76564 2592 76616 2644
rect 78588 2592 78640 2644
rect 79508 2592 79560 2644
rect 79600 2592 79652 2644
rect 80888 2592 80940 2644
rect 81624 2592 81676 2644
rect 82544 2592 82596 2644
rect 83740 2592 83792 2644
rect 85120 2592 85172 2644
rect 86592 2592 86644 2644
rect 88340 2592 88392 2644
rect 88800 2635 88852 2644
rect 88800 2601 88809 2635
rect 88809 2601 88843 2635
rect 88843 2601 88852 2635
rect 88800 2592 88852 2601
rect 90824 2592 90876 2644
rect 92204 2592 92256 2644
rect 93124 2635 93176 2644
rect 93124 2601 93133 2635
rect 93133 2601 93167 2635
rect 93167 2601 93176 2635
rect 93124 2592 93176 2601
rect 93952 2635 94004 2644
rect 93952 2601 93961 2635
rect 93961 2601 93995 2635
rect 93995 2601 94004 2635
rect 93952 2592 94004 2601
rect 95792 2592 95844 2644
rect 96252 2592 96304 2644
rect 97908 2592 97960 2644
rect 100300 2635 100352 2644
rect 60280 2456 60332 2508
rect 60648 2456 60700 2508
rect 60832 2456 60884 2508
rect 61292 2456 61344 2508
rect 97540 2524 97592 2576
rect 97724 2567 97776 2576
rect 97724 2533 97733 2567
rect 97733 2533 97767 2567
rect 97767 2533 97776 2567
rect 97724 2524 97776 2533
rect 664 2252 716 2304
rect 2044 2252 2096 2304
rect 3516 2252 3568 2304
rect 4896 2252 4948 2304
rect 6368 2252 6420 2304
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 12164 2431 12216 2440
rect 12164 2397 12173 2431
rect 12173 2397 12207 2431
rect 12207 2397 12216 2431
rect 12164 2388 12216 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 22008 2388 22060 2440
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 7748 2252 7800 2304
rect 9220 2252 9272 2304
rect 10600 2252 10652 2304
rect 12072 2252 12124 2304
rect 13452 2252 13504 2304
rect 14924 2320 14976 2372
rect 15476 2363 15528 2372
rect 15476 2329 15485 2363
rect 15485 2329 15519 2363
rect 15519 2329 15528 2363
rect 15476 2320 15528 2329
rect 16304 2320 16356 2372
rect 17776 2320 17828 2372
rect 18328 2363 18380 2372
rect 18328 2329 18337 2363
rect 18337 2329 18371 2363
rect 18371 2329 18380 2363
rect 18328 2320 18380 2329
rect 19156 2320 19208 2372
rect 20628 2320 20680 2372
rect 19432 2252 19484 2304
rect 19984 2252 20036 2304
rect 23480 2320 23532 2372
rect 24952 2320 25004 2372
rect 25780 2388 25832 2440
rect 35716 2388 35768 2440
rect 35808 2388 35860 2440
rect 26240 2320 26292 2372
rect 26332 2320 26384 2372
rect 27712 2320 27764 2372
rect 29184 2320 29236 2372
rect 30012 2363 30064 2372
rect 30012 2329 30021 2363
rect 30021 2329 30055 2363
rect 30055 2329 30064 2363
rect 30012 2320 30064 2329
rect 30840 2363 30892 2372
rect 30840 2329 30849 2363
rect 30849 2329 30883 2363
rect 30883 2329 30892 2363
rect 30840 2320 30892 2329
rect 24768 2295 24820 2304
rect 24768 2261 24777 2295
rect 24777 2261 24811 2295
rect 24811 2261 24820 2295
rect 24768 2252 24820 2261
rect 25688 2295 25740 2304
rect 25688 2261 25697 2295
rect 25697 2261 25731 2295
rect 25731 2261 25740 2295
rect 27344 2295 27396 2304
rect 25688 2252 25740 2261
rect 27344 2261 27353 2295
rect 27353 2261 27387 2295
rect 27387 2261 27396 2295
rect 27344 2252 27396 2261
rect 31668 2252 31720 2304
rect 32036 2320 32088 2372
rect 32588 2363 32640 2372
rect 32588 2329 32597 2363
rect 32597 2329 32631 2363
rect 32631 2329 32640 2363
rect 32588 2320 32640 2329
rect 33416 2320 33468 2372
rect 33508 2320 33560 2372
rect 35164 2363 35216 2372
rect 35164 2329 35173 2363
rect 35173 2329 35207 2363
rect 35207 2329 35216 2363
rect 35164 2320 35216 2329
rect 37280 2320 37332 2372
rect 35532 2252 35584 2304
rect 36360 2252 36412 2304
rect 37740 2320 37792 2372
rect 39212 2320 39264 2372
rect 40592 2320 40644 2372
rect 42064 2320 42116 2372
rect 43444 2320 43496 2372
rect 44916 2320 44968 2372
rect 46296 2320 46348 2372
rect 47676 2320 47728 2372
rect 47768 2320 47820 2372
rect 37648 2295 37700 2304
rect 37648 2261 37657 2295
rect 37657 2261 37691 2295
rect 37691 2261 37700 2295
rect 37648 2252 37700 2261
rect 38568 2295 38620 2304
rect 38568 2261 38577 2295
rect 38577 2261 38611 2295
rect 38611 2261 38620 2295
rect 38568 2252 38620 2261
rect 40500 2252 40552 2304
rect 41144 2295 41196 2304
rect 41144 2261 41153 2295
rect 41153 2261 41187 2295
rect 41187 2261 41196 2295
rect 41144 2252 41196 2261
rect 42800 2295 42852 2304
rect 42800 2261 42809 2295
rect 42809 2261 42843 2295
rect 42843 2261 42852 2295
rect 42800 2252 42852 2261
rect 43904 2295 43956 2304
rect 43904 2261 43913 2295
rect 43913 2261 43947 2295
rect 43947 2261 43956 2295
rect 43904 2252 43956 2261
rect 45192 2295 45244 2304
rect 45192 2261 45201 2295
rect 45201 2261 45235 2295
rect 45235 2261 45244 2295
rect 45192 2252 45244 2261
rect 45376 2252 45428 2304
rect 49056 2320 49108 2372
rect 49148 2320 49200 2372
rect 49608 2252 49660 2304
rect 50620 2320 50672 2372
rect 51908 2320 51960 2372
rect 52000 2320 52052 2372
rect 53380 2320 53432 2372
rect 53472 2320 53524 2372
rect 55680 2252 55732 2304
rect 56140 2252 56192 2304
rect 56692 2320 56744 2372
rect 57704 2320 57756 2372
rect 59544 2363 59596 2372
rect 59544 2329 59553 2363
rect 59553 2329 59587 2363
rect 59587 2329 59596 2363
rect 59544 2320 59596 2329
rect 59912 2388 59964 2440
rect 62120 2431 62172 2440
rect 62120 2397 62129 2431
rect 62129 2397 62163 2431
rect 62163 2397 62172 2431
rect 62120 2388 62172 2397
rect 63408 2388 63460 2440
rect 64420 2388 64472 2440
rect 65524 2388 65576 2440
rect 66720 2431 66772 2440
rect 66720 2397 66729 2431
rect 66729 2397 66763 2431
rect 66763 2397 66772 2431
rect 66720 2388 66772 2397
rect 68284 2431 68336 2440
rect 68284 2397 68293 2431
rect 68293 2397 68327 2431
rect 68327 2397 68336 2431
rect 68284 2388 68336 2397
rect 69572 2431 69624 2440
rect 69572 2397 69581 2431
rect 69581 2397 69615 2431
rect 69615 2397 69624 2431
rect 69572 2388 69624 2397
rect 69664 2388 69716 2440
rect 72792 2431 72844 2440
rect 60188 2320 60240 2372
rect 61016 2363 61068 2372
rect 61016 2329 61025 2363
rect 61025 2329 61059 2363
rect 61059 2329 61068 2363
rect 61016 2320 61068 2329
rect 63132 2363 63184 2372
rect 63132 2329 63141 2363
rect 63141 2329 63175 2363
rect 63175 2329 63184 2363
rect 63132 2320 63184 2329
rect 63316 2320 63368 2372
rect 59636 2252 59688 2304
rect 59728 2252 59780 2304
rect 61936 2252 61988 2304
rect 62028 2252 62080 2304
rect 65156 2252 65208 2304
rect 66812 2295 66864 2304
rect 66812 2261 66821 2295
rect 66821 2261 66855 2295
rect 66855 2261 66864 2295
rect 66812 2252 66864 2261
rect 67456 2252 67508 2304
rect 69756 2320 69808 2372
rect 71688 2320 71740 2372
rect 72792 2397 72801 2431
rect 72801 2397 72835 2431
rect 72835 2397 72844 2431
rect 72792 2388 72844 2397
rect 73528 2431 73580 2440
rect 73528 2397 73537 2431
rect 73537 2397 73571 2431
rect 73571 2397 73580 2431
rect 73528 2388 73580 2397
rect 74816 2456 74868 2508
rect 75000 2456 75052 2508
rect 79232 2499 79284 2508
rect 79232 2465 79241 2499
rect 79241 2465 79275 2499
rect 79275 2465 79284 2499
rect 79232 2456 79284 2465
rect 81532 2499 81584 2508
rect 79416 2388 79468 2440
rect 73344 2252 73396 2304
rect 73436 2252 73488 2304
rect 73896 2320 73948 2372
rect 76104 2320 76156 2372
rect 76196 2320 76248 2372
rect 81532 2465 81541 2499
rect 81541 2465 81575 2499
rect 81575 2465 81584 2499
rect 81532 2456 81584 2465
rect 81440 2388 81492 2440
rect 83556 2456 83608 2508
rect 84936 2456 84988 2508
rect 85580 2456 85632 2508
rect 86408 2456 86460 2508
rect 74448 2252 74500 2304
rect 75000 2295 75052 2304
rect 75000 2261 75009 2295
rect 75009 2261 75043 2295
rect 75043 2261 75052 2295
rect 75000 2252 75052 2261
rect 76472 2252 76524 2304
rect 77576 2295 77628 2304
rect 77576 2261 77585 2295
rect 77585 2261 77619 2295
rect 77619 2261 77628 2295
rect 77576 2252 77628 2261
rect 77668 2295 77720 2304
rect 77668 2261 77677 2295
rect 77677 2261 77711 2295
rect 77711 2261 77720 2295
rect 79048 2295 79100 2304
rect 77668 2252 77720 2261
rect 79048 2261 79057 2295
rect 79057 2261 79091 2295
rect 79091 2261 79100 2295
rect 84108 2320 84160 2372
rect 79048 2252 79100 2261
rect 80520 2252 80572 2304
rect 83096 2295 83148 2304
rect 83096 2261 83105 2295
rect 83105 2261 83139 2295
rect 83139 2261 83148 2295
rect 83096 2252 83148 2261
rect 84016 2295 84068 2304
rect 84016 2261 84025 2295
rect 84025 2261 84059 2295
rect 84059 2261 84068 2295
rect 84016 2252 84068 2261
rect 85028 2388 85080 2440
rect 86868 2456 86920 2508
rect 87788 2456 87840 2508
rect 89260 2499 89312 2508
rect 89260 2465 89269 2499
rect 89269 2465 89303 2499
rect 89303 2465 89312 2499
rect 89260 2456 89312 2465
rect 90548 2499 90600 2508
rect 90548 2465 90557 2499
rect 90557 2465 90591 2499
rect 90591 2465 90600 2499
rect 90548 2456 90600 2465
rect 89444 2388 89496 2440
rect 91560 2456 91612 2508
rect 92296 2456 92348 2508
rect 95516 2499 95568 2508
rect 95516 2465 95525 2499
rect 95525 2465 95559 2499
rect 95559 2465 95568 2499
rect 95516 2456 95568 2465
rect 96988 2499 97040 2508
rect 92940 2431 92992 2440
rect 92940 2397 92949 2431
rect 92949 2397 92983 2431
rect 92983 2397 92992 2431
rect 92940 2388 92992 2397
rect 93492 2388 93544 2440
rect 96988 2465 96997 2499
rect 96997 2465 97031 2499
rect 97031 2465 97040 2499
rect 96988 2456 97040 2465
rect 98000 2456 98052 2508
rect 100300 2601 100309 2635
rect 100309 2601 100343 2635
rect 100343 2601 100352 2635
rect 100300 2592 100352 2601
rect 102140 2592 102192 2644
rect 104256 2592 104308 2644
rect 105820 2592 105872 2644
rect 108304 2592 108356 2644
rect 110512 2592 110564 2644
rect 114100 2592 114152 2644
rect 116584 2592 116636 2644
rect 99104 2567 99156 2576
rect 99104 2533 99113 2567
rect 99113 2533 99147 2567
rect 99147 2533 99156 2567
rect 99104 2524 99156 2533
rect 99564 2524 99616 2576
rect 99748 2524 99800 2576
rect 100300 2456 100352 2508
rect 100392 2456 100444 2508
rect 106188 2524 106240 2576
rect 102324 2499 102376 2508
rect 102324 2465 102333 2499
rect 102333 2465 102367 2499
rect 102367 2465 102376 2499
rect 103520 2499 103572 2508
rect 102324 2456 102376 2465
rect 103520 2465 103529 2499
rect 103529 2465 103563 2499
rect 103563 2465 103572 2499
rect 103520 2456 103572 2465
rect 102968 2388 103020 2440
rect 84292 2320 84344 2372
rect 85580 2252 85632 2304
rect 86592 2295 86644 2304
rect 86592 2261 86601 2295
rect 86601 2261 86635 2295
rect 86635 2261 86644 2295
rect 86592 2252 86644 2261
rect 87880 2295 87932 2304
rect 87880 2261 87889 2295
rect 87889 2261 87923 2295
rect 87923 2261 87932 2295
rect 87880 2252 87932 2261
rect 88340 2252 88392 2304
rect 90456 2295 90508 2304
rect 90456 2261 90465 2295
rect 90465 2261 90499 2295
rect 90499 2261 90508 2295
rect 90456 2252 90508 2261
rect 91928 2295 91980 2304
rect 91928 2261 91937 2295
rect 91937 2261 91971 2295
rect 91971 2261 91980 2295
rect 91928 2252 91980 2261
rect 95424 2295 95476 2304
rect 95424 2261 95433 2295
rect 95433 2261 95467 2295
rect 95467 2261 95476 2295
rect 95424 2252 95476 2261
rect 96896 2295 96948 2304
rect 96896 2261 96905 2295
rect 96905 2261 96939 2295
rect 96939 2261 96948 2295
rect 96896 2252 96948 2261
rect 98092 2295 98144 2304
rect 98092 2261 98101 2295
rect 98101 2261 98135 2295
rect 98135 2261 98144 2295
rect 98092 2252 98144 2261
rect 99472 2363 99524 2372
rect 99472 2329 99481 2363
rect 99481 2329 99515 2363
rect 99515 2329 99524 2363
rect 99472 2320 99524 2329
rect 103428 2320 103480 2372
rect 100668 2295 100720 2304
rect 100668 2261 100677 2295
rect 100677 2261 100711 2295
rect 100711 2261 100720 2295
rect 100668 2252 100720 2261
rect 100760 2252 100812 2304
rect 103244 2295 103296 2304
rect 103244 2261 103253 2295
rect 103253 2261 103287 2295
rect 103287 2261 103296 2295
rect 103244 2252 103296 2261
rect 105176 2456 105228 2508
rect 105452 2431 105504 2440
rect 105452 2397 105461 2431
rect 105461 2397 105495 2431
rect 105495 2397 105504 2431
rect 105452 2388 105504 2397
rect 107660 2456 107712 2508
rect 110696 2524 110748 2576
rect 115848 2524 115900 2576
rect 109960 2499 110012 2508
rect 109960 2465 109969 2499
rect 109969 2465 110003 2499
rect 110003 2465 110012 2499
rect 109960 2456 110012 2465
rect 110604 2456 110656 2508
rect 105728 2388 105780 2440
rect 109040 2388 109092 2440
rect 109132 2388 109184 2440
rect 112076 2456 112128 2508
rect 112628 2499 112680 2508
rect 112628 2465 112637 2499
rect 112637 2465 112671 2499
rect 112671 2465 112680 2499
rect 112628 2456 112680 2465
rect 113548 2456 113600 2508
rect 115388 2499 115440 2508
rect 115388 2465 115397 2499
rect 115397 2465 115431 2499
rect 115431 2465 115440 2499
rect 115388 2456 115440 2465
rect 115480 2499 115532 2508
rect 115480 2465 115489 2499
rect 115489 2465 115523 2499
rect 115523 2465 115532 2499
rect 115480 2456 115532 2465
rect 119160 2456 119212 2508
rect 116492 2431 116544 2440
rect 116492 2397 116501 2431
rect 116501 2397 116535 2431
rect 116535 2397 116544 2431
rect 116492 2388 116544 2397
rect 117596 2431 117648 2440
rect 117596 2397 117605 2431
rect 117605 2397 117639 2431
rect 117639 2397 117648 2431
rect 117596 2388 117648 2397
rect 106188 2320 106240 2372
rect 108672 2363 108724 2372
rect 108672 2329 108681 2363
rect 108681 2329 108715 2363
rect 108715 2329 108724 2363
rect 108672 2320 108724 2329
rect 112536 2320 112588 2372
rect 113640 2363 113692 2372
rect 113640 2329 113649 2363
rect 113649 2329 113683 2363
rect 113683 2329 113692 2363
rect 113640 2320 113692 2329
rect 116768 2363 116820 2372
rect 116768 2329 116777 2363
rect 116777 2329 116811 2363
rect 116811 2329 116820 2363
rect 116768 2320 116820 2329
rect 109776 2295 109828 2304
rect 109776 2261 109785 2295
rect 109785 2261 109819 2295
rect 109819 2261 109828 2295
rect 109776 2252 109828 2261
rect 111524 2295 111576 2304
rect 111524 2261 111533 2295
rect 111533 2261 111567 2295
rect 111567 2261 111576 2295
rect 111524 2252 111576 2261
rect 115296 2295 115348 2304
rect 115296 2261 115305 2295
rect 115305 2261 115339 2295
rect 115339 2261 115348 2295
rect 115296 2252 115348 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 81014 2150 81066 2202
rect 81078 2150 81130 2202
rect 81142 2150 81194 2202
rect 81206 2150 81258 2202
rect 81270 2150 81322 2202
rect 111734 2150 111786 2202
rect 111798 2150 111850 2202
rect 111862 2150 111914 2202
rect 111926 2150 111978 2202
rect 111990 2150 112042 2202
rect 2136 2048 2188 2100
rect 51080 2048 51132 2100
rect 3792 1980 3844 2032
rect 60188 2048 60240 2100
rect 60372 2048 60424 2100
rect 66812 2048 66864 2100
rect 66904 2048 66956 2100
rect 113640 2048 113692 2100
rect 51356 1980 51408 2032
rect 59820 1980 59872 2032
rect 24768 1912 24820 1964
rect 61936 1980 61988 2032
rect 111524 1980 111576 2032
rect 76012 1912 76064 1964
rect 76104 1912 76156 1964
rect 80520 1912 80572 1964
rect 80888 1912 80940 1964
rect 84752 1912 84804 1964
rect 103520 1912 103572 1964
rect 108672 1912 108724 1964
rect 19432 1844 19484 1896
rect 25780 1844 25832 1896
rect 26240 1844 26292 1896
rect 35624 1844 35676 1896
rect 27344 1776 27396 1828
rect 60740 1844 60792 1896
rect 60924 1844 60976 1896
rect 35808 1776 35860 1828
rect 79140 1776 79192 1828
rect 19984 1708 20036 1760
rect 79048 1708 79100 1760
rect 79324 1844 79376 1896
rect 79508 1844 79560 1896
rect 91468 1844 91520 1896
rect 100300 1844 100352 1896
rect 117596 1844 117648 1896
rect 87880 1776 87932 1828
rect 86592 1708 86644 1760
rect 10692 1640 10744 1692
rect 63316 1640 63368 1692
rect 66168 1640 66220 1692
rect 70216 1640 70268 1692
rect 70308 1640 70360 1692
rect 73896 1640 73948 1692
rect 73988 1640 74040 1692
rect 99472 1640 99524 1692
rect 12164 1572 12216 1624
rect 45560 1572 45612 1624
rect 45652 1572 45704 1624
rect 7840 1504 7892 1556
rect 51080 1504 51132 1556
rect 51264 1504 51316 1556
rect 60556 1504 60608 1556
rect 99380 1572 99432 1624
rect 61752 1504 61804 1556
rect 115296 1504 115348 1556
rect 14096 1436 14148 1488
rect 45652 1436 45704 1488
rect 45744 1436 45796 1488
rect 51172 1436 51224 1488
rect 51632 1436 51684 1488
rect 60464 1436 60516 1488
rect 61016 1436 61068 1488
rect 105268 1436 105320 1488
rect 7104 1368 7156 1420
rect 51264 1368 51316 1420
rect 45560 1300 45612 1352
rect 60740 1368 60792 1420
rect 61200 1368 61252 1420
rect 72792 1368 72844 1420
rect 72884 1368 72936 1420
rect 77576 1368 77628 1420
rect 77668 1368 77720 1420
rect 84016 1368 84068 1420
rect 84752 1368 84804 1420
rect 98460 1368 98512 1420
rect 99196 1368 99248 1420
rect 101220 1368 101272 1420
rect 56324 1300 56376 1352
rect 61752 1300 61804 1352
rect 65524 1300 65576 1352
rect 109776 1300 109828 1352
rect 35532 1232 35584 1284
rect 95424 1232 95476 1284
rect 45652 1164 45704 1216
rect 51632 1164 51684 1216
rect 61384 1164 61436 1216
rect 116768 1164 116820 1216
rect 38568 1096 38620 1148
rect 98092 1096 98144 1148
rect 41144 1028 41196 1080
rect 100668 1028 100720 1080
rect 32588 960 32640 1012
rect 91928 960 91980 1012
rect 31668 892 31720 944
rect 90456 892 90508 944
rect 43904 824 43956 876
rect 103244 824 103296 876
rect 30012 756 30064 808
rect 88340 756 88392 808
rect 37648 688 37700 740
rect 96896 688 96948 740
rect 42800 620 42852 672
rect 100760 620 100812 672
rect 18328 552 18380 604
rect 72884 552 72936 604
rect 15476 484 15528 536
rect 75000 484 75052 536
rect 49608 348 49660 400
rect 65524 348 65576 400
<< metal2 >>
rect 117134 39536 117190 39545
rect 117134 39471 117190 39480
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 65654 37564 65962 37584
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37488 65962 37508
rect 96374 37564 96682 37584
rect 96374 37562 96380 37564
rect 96436 37562 96460 37564
rect 96516 37562 96540 37564
rect 96596 37562 96620 37564
rect 96676 37562 96682 37564
rect 96436 37510 96438 37562
rect 96618 37510 96620 37562
rect 96374 37508 96380 37510
rect 96436 37508 96460 37510
rect 96516 37508 96540 37510
rect 96596 37508 96620 37510
rect 96676 37508 96682 37510
rect 96374 37488 96682 37508
rect 114928 37256 114980 37262
rect 114928 37198 114980 37204
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 81014 37020 81322 37040
rect 81014 37018 81020 37020
rect 81076 37018 81100 37020
rect 81156 37018 81180 37020
rect 81236 37018 81260 37020
rect 81316 37018 81322 37020
rect 81076 36966 81078 37018
rect 81258 36966 81260 37018
rect 81014 36964 81020 36966
rect 81076 36964 81100 36966
rect 81156 36964 81180 36966
rect 81236 36964 81260 36966
rect 81316 36964 81322 36966
rect 81014 36944 81322 36964
rect 111734 37020 112042 37040
rect 111734 37018 111740 37020
rect 111796 37018 111820 37020
rect 111876 37018 111900 37020
rect 111956 37018 111980 37020
rect 112036 37018 112042 37020
rect 111796 36966 111798 37018
rect 111978 36966 111980 37018
rect 111734 36964 111740 36966
rect 111796 36964 111820 36966
rect 111876 36964 111900 36966
rect 111956 36964 111980 36966
rect 112036 36964 112042 36966
rect 111734 36944 112042 36964
rect 98920 36780 98972 36786
rect 98920 36722 98972 36728
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 65654 36476 65962 36496
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36400 65962 36420
rect 96374 36476 96682 36496
rect 96374 36474 96380 36476
rect 96436 36474 96460 36476
rect 96516 36474 96540 36476
rect 96596 36474 96620 36476
rect 96676 36474 96682 36476
rect 96436 36422 96438 36474
rect 96618 36422 96620 36474
rect 96374 36420 96380 36422
rect 96436 36420 96460 36422
rect 96516 36420 96540 36422
rect 96596 36420 96620 36422
rect 96676 36420 96682 36422
rect 96374 36400 96682 36420
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 81014 35932 81322 35952
rect 81014 35930 81020 35932
rect 81076 35930 81100 35932
rect 81156 35930 81180 35932
rect 81236 35930 81260 35932
rect 81316 35930 81322 35932
rect 81076 35878 81078 35930
rect 81258 35878 81260 35930
rect 81014 35876 81020 35878
rect 81076 35876 81100 35878
rect 81156 35876 81180 35878
rect 81236 35876 81260 35878
rect 81316 35876 81322 35878
rect 81014 35856 81322 35876
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 65654 35388 65962 35408
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35312 65962 35332
rect 96374 35388 96682 35408
rect 96374 35386 96380 35388
rect 96436 35386 96460 35388
rect 96516 35386 96540 35388
rect 96596 35386 96620 35388
rect 96676 35386 96682 35388
rect 96436 35334 96438 35386
rect 96618 35334 96620 35386
rect 96374 35332 96380 35334
rect 96436 35332 96460 35334
rect 96516 35332 96540 35334
rect 96596 35332 96620 35334
rect 96676 35332 96682 35334
rect 96374 35312 96682 35332
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 81014 34844 81322 34864
rect 81014 34842 81020 34844
rect 81076 34842 81100 34844
rect 81156 34842 81180 34844
rect 81236 34842 81260 34844
rect 81316 34842 81322 34844
rect 81076 34790 81078 34842
rect 81258 34790 81260 34842
rect 81014 34788 81020 34790
rect 81076 34788 81100 34790
rect 81156 34788 81180 34790
rect 81236 34788 81260 34790
rect 81316 34788 81322 34790
rect 81014 34768 81322 34788
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 65654 34300 65962 34320
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34224 65962 34244
rect 96374 34300 96682 34320
rect 96374 34298 96380 34300
rect 96436 34298 96460 34300
rect 96516 34298 96540 34300
rect 96596 34298 96620 34300
rect 96676 34298 96682 34300
rect 96436 34246 96438 34298
rect 96618 34246 96620 34298
rect 96374 34244 96380 34246
rect 96436 34244 96460 34246
rect 96516 34244 96540 34246
rect 96596 34244 96620 34246
rect 96676 34244 96682 34246
rect 96374 34224 96682 34244
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 81014 33756 81322 33776
rect 81014 33754 81020 33756
rect 81076 33754 81100 33756
rect 81156 33754 81180 33756
rect 81236 33754 81260 33756
rect 81316 33754 81322 33756
rect 81076 33702 81078 33754
rect 81258 33702 81260 33754
rect 81014 33700 81020 33702
rect 81076 33700 81100 33702
rect 81156 33700 81180 33702
rect 81236 33700 81260 33702
rect 81316 33700 81322 33702
rect 81014 33680 81322 33700
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 65654 33212 65962 33232
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33136 65962 33156
rect 96374 33212 96682 33232
rect 96374 33210 96380 33212
rect 96436 33210 96460 33212
rect 96516 33210 96540 33212
rect 96596 33210 96620 33212
rect 96676 33210 96682 33212
rect 96436 33158 96438 33210
rect 96618 33158 96620 33210
rect 96374 33156 96380 33158
rect 96436 33156 96460 33158
rect 96516 33156 96540 33158
rect 96596 33156 96620 33158
rect 96676 33156 96682 33158
rect 96374 33136 96682 33156
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 81014 32668 81322 32688
rect 81014 32666 81020 32668
rect 81076 32666 81100 32668
rect 81156 32666 81180 32668
rect 81236 32666 81260 32668
rect 81316 32666 81322 32668
rect 81076 32614 81078 32666
rect 81258 32614 81260 32666
rect 81014 32612 81020 32614
rect 81076 32612 81100 32614
rect 81156 32612 81180 32614
rect 81236 32612 81260 32614
rect 81316 32612 81322 32614
rect 81014 32592 81322 32612
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 65654 32124 65962 32144
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32048 65962 32068
rect 96374 32124 96682 32144
rect 96374 32122 96380 32124
rect 96436 32122 96460 32124
rect 96516 32122 96540 32124
rect 96596 32122 96620 32124
rect 96676 32122 96682 32124
rect 96436 32070 96438 32122
rect 96618 32070 96620 32122
rect 96374 32068 96380 32070
rect 96436 32068 96460 32070
rect 96516 32068 96540 32070
rect 96596 32068 96620 32070
rect 96676 32068 96682 32070
rect 96374 32048 96682 32068
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 81014 31580 81322 31600
rect 81014 31578 81020 31580
rect 81076 31578 81100 31580
rect 81156 31578 81180 31580
rect 81236 31578 81260 31580
rect 81316 31578 81322 31580
rect 81076 31526 81078 31578
rect 81258 31526 81260 31578
rect 81014 31524 81020 31526
rect 81076 31524 81100 31526
rect 81156 31524 81180 31526
rect 81236 31524 81260 31526
rect 81316 31524 81322 31526
rect 81014 31504 81322 31524
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 65654 31036 65962 31056
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30960 65962 30980
rect 96374 31036 96682 31056
rect 96374 31034 96380 31036
rect 96436 31034 96460 31036
rect 96516 31034 96540 31036
rect 96596 31034 96620 31036
rect 96676 31034 96682 31036
rect 96436 30982 96438 31034
rect 96618 30982 96620 31034
rect 96374 30980 96380 30982
rect 96436 30980 96460 30982
rect 96516 30980 96540 30982
rect 96596 30980 96620 30982
rect 96676 30980 96682 30982
rect 96374 30960 96682 30980
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 81014 30492 81322 30512
rect 81014 30490 81020 30492
rect 81076 30490 81100 30492
rect 81156 30490 81180 30492
rect 81236 30490 81260 30492
rect 81316 30490 81322 30492
rect 81076 30438 81078 30490
rect 81258 30438 81260 30490
rect 81014 30436 81020 30438
rect 81076 30436 81100 30438
rect 81156 30436 81180 30438
rect 81236 30436 81260 30438
rect 81316 30436 81322 30438
rect 81014 30416 81322 30436
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 65654 29948 65962 29968
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29872 65962 29892
rect 96374 29948 96682 29968
rect 96374 29946 96380 29948
rect 96436 29946 96460 29948
rect 96516 29946 96540 29948
rect 96596 29946 96620 29948
rect 96676 29946 96682 29948
rect 96436 29894 96438 29946
rect 96618 29894 96620 29946
rect 96374 29892 96380 29894
rect 96436 29892 96460 29894
rect 96516 29892 96540 29894
rect 96596 29892 96620 29894
rect 96676 29892 96682 29894
rect 96374 29872 96682 29892
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 81014 29404 81322 29424
rect 81014 29402 81020 29404
rect 81076 29402 81100 29404
rect 81156 29402 81180 29404
rect 81236 29402 81260 29404
rect 81316 29402 81322 29404
rect 81076 29350 81078 29402
rect 81258 29350 81260 29402
rect 81014 29348 81020 29350
rect 81076 29348 81100 29350
rect 81156 29348 81180 29350
rect 81236 29348 81260 29350
rect 81316 29348 81322 29350
rect 81014 29328 81322 29348
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 65654 28860 65962 28880
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28784 65962 28804
rect 96374 28860 96682 28880
rect 96374 28858 96380 28860
rect 96436 28858 96460 28860
rect 96516 28858 96540 28860
rect 96596 28858 96620 28860
rect 96676 28858 96682 28860
rect 96436 28806 96438 28858
rect 96618 28806 96620 28858
rect 96374 28804 96380 28806
rect 96436 28804 96460 28806
rect 96516 28804 96540 28806
rect 96596 28804 96620 28806
rect 96676 28804 96682 28806
rect 96374 28784 96682 28804
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 81014 28316 81322 28336
rect 81014 28314 81020 28316
rect 81076 28314 81100 28316
rect 81156 28314 81180 28316
rect 81236 28314 81260 28316
rect 81316 28314 81322 28316
rect 81076 28262 81078 28314
rect 81258 28262 81260 28314
rect 81014 28260 81020 28262
rect 81076 28260 81100 28262
rect 81156 28260 81180 28262
rect 81236 28260 81260 28262
rect 81316 28260 81322 28262
rect 81014 28240 81322 28260
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 65654 27772 65962 27792
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27696 65962 27716
rect 96374 27772 96682 27792
rect 96374 27770 96380 27772
rect 96436 27770 96460 27772
rect 96516 27770 96540 27772
rect 96596 27770 96620 27772
rect 96676 27770 96682 27772
rect 96436 27718 96438 27770
rect 96618 27718 96620 27770
rect 96374 27716 96380 27718
rect 96436 27716 96460 27718
rect 96516 27716 96540 27718
rect 96596 27716 96620 27718
rect 96676 27716 96682 27718
rect 96374 27696 96682 27716
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 81014 27228 81322 27248
rect 81014 27226 81020 27228
rect 81076 27226 81100 27228
rect 81156 27226 81180 27228
rect 81236 27226 81260 27228
rect 81316 27226 81322 27228
rect 81076 27174 81078 27226
rect 81258 27174 81260 27226
rect 81014 27172 81020 27174
rect 81076 27172 81100 27174
rect 81156 27172 81180 27174
rect 81236 27172 81260 27174
rect 81316 27172 81322 27174
rect 81014 27152 81322 27172
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 65654 26684 65962 26704
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26608 65962 26628
rect 96374 26684 96682 26704
rect 96374 26682 96380 26684
rect 96436 26682 96460 26684
rect 96516 26682 96540 26684
rect 96596 26682 96620 26684
rect 96676 26682 96682 26684
rect 96436 26630 96438 26682
rect 96618 26630 96620 26682
rect 96374 26628 96380 26630
rect 96436 26628 96460 26630
rect 96516 26628 96540 26630
rect 96596 26628 96620 26630
rect 96676 26628 96682 26630
rect 96374 26608 96682 26628
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 81014 26140 81322 26160
rect 81014 26138 81020 26140
rect 81076 26138 81100 26140
rect 81156 26138 81180 26140
rect 81236 26138 81260 26140
rect 81316 26138 81322 26140
rect 81076 26086 81078 26138
rect 81258 26086 81260 26138
rect 81014 26084 81020 26086
rect 81076 26084 81100 26086
rect 81156 26084 81180 26086
rect 81236 26084 81260 26086
rect 81316 26084 81322 26086
rect 81014 26064 81322 26084
rect 98092 25900 98144 25906
rect 98092 25842 98144 25848
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 65654 25596 65962 25616
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25520 65962 25540
rect 96374 25596 96682 25616
rect 96374 25594 96380 25596
rect 96436 25594 96460 25596
rect 96516 25594 96540 25596
rect 96596 25594 96620 25596
rect 96676 25594 96682 25596
rect 96436 25542 96438 25594
rect 96618 25542 96620 25594
rect 96374 25540 96380 25542
rect 96436 25540 96460 25542
rect 96516 25540 96540 25542
rect 96596 25540 96620 25542
rect 96676 25540 96682 25542
rect 96374 25520 96682 25540
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 81014 25052 81322 25072
rect 81014 25050 81020 25052
rect 81076 25050 81100 25052
rect 81156 25050 81180 25052
rect 81236 25050 81260 25052
rect 81316 25050 81322 25052
rect 81076 24998 81078 25050
rect 81258 24998 81260 25050
rect 81014 24996 81020 24998
rect 81076 24996 81100 24998
rect 81156 24996 81180 24998
rect 81236 24996 81260 24998
rect 81316 24996 81322 24998
rect 81014 24976 81322 24996
rect 96896 24812 96948 24818
rect 96896 24754 96948 24760
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 65654 24508 65962 24528
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24432 65962 24452
rect 96374 24508 96682 24528
rect 96374 24506 96380 24508
rect 96436 24506 96460 24508
rect 96516 24506 96540 24508
rect 96596 24506 96620 24508
rect 96676 24506 96682 24508
rect 96436 24454 96438 24506
rect 96618 24454 96620 24506
rect 96374 24452 96380 24454
rect 96436 24452 96460 24454
rect 96516 24452 96540 24454
rect 96596 24452 96620 24454
rect 96676 24452 96682 24454
rect 96374 24432 96682 24452
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 81014 23964 81322 23984
rect 81014 23962 81020 23964
rect 81076 23962 81100 23964
rect 81156 23962 81180 23964
rect 81236 23962 81260 23964
rect 81316 23962 81322 23964
rect 81076 23910 81078 23962
rect 81258 23910 81260 23962
rect 81014 23908 81020 23910
rect 81076 23908 81100 23910
rect 81156 23908 81180 23910
rect 81236 23908 81260 23910
rect 81316 23908 81322 23910
rect 81014 23888 81322 23908
rect 95976 23724 96028 23730
rect 95976 23666 96028 23672
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 65654 23420 65962 23440
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23344 65962 23364
rect 93124 23112 93176 23118
rect 93124 23054 93176 23060
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 81014 22876 81322 22896
rect 81014 22874 81020 22876
rect 81076 22874 81100 22876
rect 81156 22874 81180 22876
rect 81236 22874 81260 22876
rect 81316 22874 81322 22876
rect 81076 22822 81078 22874
rect 81258 22822 81260 22874
rect 81014 22820 81020 22822
rect 81076 22820 81100 22822
rect 81156 22820 81180 22822
rect 81236 22820 81260 22822
rect 81316 22820 81322 22822
rect 81014 22800 81322 22820
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 65654 22332 65962 22352
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22256 65962 22276
rect 92388 21888 92440 21894
rect 92388 21830 92440 21836
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 81014 21788 81322 21808
rect 81014 21786 81020 21788
rect 81076 21786 81100 21788
rect 81156 21786 81180 21788
rect 81236 21786 81260 21788
rect 81316 21786 81322 21788
rect 81076 21734 81078 21786
rect 81258 21734 81260 21786
rect 81014 21732 81020 21734
rect 81076 21732 81100 21734
rect 81156 21732 81180 21734
rect 81236 21732 81260 21734
rect 81316 21732 81322 21734
rect 81014 21712 81322 21732
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 65654 21244 65962 21264
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21168 65962 21188
rect 91008 20936 91060 20942
rect 91008 20878 91060 20884
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 81014 20700 81322 20720
rect 81014 20698 81020 20700
rect 81076 20698 81100 20700
rect 81156 20698 81180 20700
rect 81236 20698 81260 20700
rect 81316 20698 81322 20700
rect 81076 20646 81078 20698
rect 81258 20646 81260 20698
rect 81014 20644 81020 20646
rect 81076 20644 81100 20646
rect 81156 20644 81180 20646
rect 81236 20644 81260 20646
rect 81316 20644 81322 20646
rect 81014 20624 81322 20644
rect 89444 20460 89496 20466
rect 89444 20402 89496 20408
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 65654 20156 65962 20176
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20080 65962 20100
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 81014 19612 81322 19632
rect 81014 19610 81020 19612
rect 81076 19610 81100 19612
rect 81156 19610 81180 19612
rect 81236 19610 81260 19612
rect 81316 19610 81322 19612
rect 81076 19558 81078 19610
rect 81258 19558 81260 19610
rect 81014 19556 81020 19558
rect 81076 19556 81100 19558
rect 81156 19556 81180 19558
rect 81236 19556 81260 19558
rect 81316 19556 81322 19558
rect 81014 19536 81322 19556
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 65654 19068 65962 19088
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 18992 65962 19012
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 81014 18524 81322 18544
rect 81014 18522 81020 18524
rect 81076 18522 81100 18524
rect 81156 18522 81180 18524
rect 81236 18522 81260 18524
rect 81316 18522 81322 18524
rect 81076 18470 81078 18522
rect 81258 18470 81260 18522
rect 81014 18468 81020 18470
rect 81076 18468 81100 18470
rect 81156 18468 81180 18470
rect 81236 18468 81260 18470
rect 81316 18468 81322 18470
rect 81014 18448 81322 18468
rect 86684 18080 86736 18086
rect 86684 18022 86736 18028
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 65654 17980 65962 18000
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17904 65962 17924
rect 85212 17672 85264 17678
rect 85212 17614 85264 17620
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 81014 17436 81322 17456
rect 81014 17434 81020 17436
rect 81076 17434 81100 17436
rect 81156 17434 81180 17436
rect 81236 17434 81260 17436
rect 81316 17434 81322 17436
rect 81076 17382 81078 17434
rect 81258 17382 81260 17434
rect 81014 17380 81020 17382
rect 81076 17380 81100 17382
rect 81156 17380 81180 17382
rect 81236 17380 81260 17382
rect 81316 17380 81322 17382
rect 81014 17360 81322 17380
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 65654 16892 65962 16912
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16816 65962 16836
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 81014 16348 81322 16368
rect 81014 16346 81020 16348
rect 81076 16346 81100 16348
rect 81156 16346 81180 16348
rect 81236 16346 81260 16348
rect 81316 16346 81322 16348
rect 81076 16294 81078 16346
rect 81258 16294 81260 16346
rect 81014 16292 81020 16294
rect 81076 16292 81100 16294
rect 81156 16292 81180 16294
rect 81236 16292 81260 16294
rect 81316 16292 81322 16294
rect 81014 16272 81322 16292
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 65654 15804 65962 15824
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15728 65962 15748
rect 82820 15496 82872 15502
rect 82820 15438 82872 15444
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 81014 15260 81322 15280
rect 81014 15258 81020 15260
rect 81076 15258 81100 15260
rect 81156 15258 81180 15260
rect 81236 15258 81260 15260
rect 81316 15258 81322 15260
rect 81076 15206 81078 15258
rect 81258 15206 81260 15258
rect 81014 15204 81020 15206
rect 81076 15204 81100 15206
rect 81156 15204 81180 15206
rect 81236 15204 81260 15206
rect 81316 15204 81322 15206
rect 81014 15184 81322 15204
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 65654 14716 65962 14736
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14640 65962 14660
rect 81716 14408 81768 14414
rect 81716 14350 81768 14356
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 81014 14172 81322 14192
rect 81014 14170 81020 14172
rect 81076 14170 81100 14172
rect 81156 14170 81180 14172
rect 81236 14170 81260 14172
rect 81316 14170 81322 14172
rect 81076 14118 81078 14170
rect 81258 14118 81260 14170
rect 81014 14116 81020 14118
rect 81076 14116 81100 14118
rect 81156 14116 81180 14118
rect 81236 14116 81260 14118
rect 81316 14116 81322 14118
rect 81014 14096 81322 14116
rect 79600 13932 79652 13938
rect 79600 13874 79652 13880
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 65654 13628 65962 13648
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13552 65962 13572
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 78680 12844 78732 12850
rect 78680 12786 78732 12792
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 65654 12540 65962 12560
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12464 65962 12484
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 76656 11552 76708 11558
rect 76656 11494 76708 11500
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 65654 11452 65962 11472
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11376 65962 11396
rect 76104 11144 76156 11150
rect 76104 11086 76156 11092
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 65654 10364 65962 10384
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10288 65962 10308
rect 76116 10266 76144 11086
rect 76104 10260 76156 10266
rect 76104 10202 76156 10208
rect 74632 10056 74684 10062
rect 74632 9998 74684 10004
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 65654 9276 65962 9296
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9200 65962 9220
rect 73528 8832 73580 8838
rect 73528 8774 73580 8780
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 65654 8188 65962 8208
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8112 65962 8132
rect 71688 7744 71740 7750
rect 71688 7686 71740 7692
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 65654 7100 65962 7120
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7024 65962 7044
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 65654 6012 65962 6032
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5936 65962 5956
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 65654 4924 65962 4944
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4848 65962 4868
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 58256 4276 58308 4282
rect 58256 4218 58308 4224
rect 25688 4208 25740 4214
rect 25688 4150 25740 4156
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 17052 2582 17080 3130
rect 17040 2576 17092 2582
rect 17040 2518 17092 2524
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 664 2304 716 2310
rect 664 2246 716 2252
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 676 800 704 2246
rect 2056 800 2084 2246
rect 2148 2106 2176 2382
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 2136 2100 2188 2106
rect 2136 2042 2188 2048
rect 3528 800 3556 2246
rect 3804 2038 3832 2382
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 3792 2032 3844 2038
rect 3792 1974 3844 1980
rect 4908 800 4936 2246
rect 6380 800 6408 2246
rect 7116 1426 7144 2246
rect 7104 1420 7156 1426
rect 7104 1362 7156 1368
rect 7760 800 7788 2246
rect 7852 1562 7880 2382
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 7840 1556 7892 1562
rect 7840 1498 7892 1504
rect 9232 800 9260 2246
rect 10612 800 10640 2246
rect 10704 1698 10732 2382
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 10692 1692 10744 1698
rect 10692 1634 10744 1640
rect 12084 800 12112 2246
rect 12176 1630 12204 2382
rect 13452 2304 13504 2310
rect 13452 2246 13504 2252
rect 12164 1624 12216 1630
rect 12164 1566 12216 1572
rect 13464 800 13492 2246
rect 14108 1494 14136 2382
rect 14924 2372 14976 2378
rect 14924 2314 14976 2320
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 19156 2372 19208 2378
rect 19156 2314 19208 2320
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 14096 1488 14148 1494
rect 14096 1430 14148 1436
rect 14936 800 14964 2314
rect 662 0 718 800
rect 2042 0 2098 800
rect 3514 0 3570 800
rect 4894 0 4950 800
rect 6366 0 6422 800
rect 7746 0 7802 800
rect 9218 0 9274 800
rect 10598 0 10654 800
rect 12070 0 12126 800
rect 13450 0 13506 800
rect 14922 0 14978 800
rect 15488 542 15516 2314
rect 16316 800 16344 2314
rect 17788 800 17816 2314
rect 15476 536 15528 542
rect 15476 478 15528 484
rect 16302 0 16358 800
rect 17774 0 17830 800
rect 18340 610 18368 2314
rect 19168 800 19196 2314
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19444 1902 19472 2246
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19432 1896 19484 1902
rect 19432 1838 19484 1844
rect 19996 1766 20024 2246
rect 19984 1760 20036 1766
rect 19984 1702 20036 1708
rect 20640 800 20668 2314
rect 22020 800 22048 2382
rect 23480 2372 23532 2378
rect 24952 2372 25004 2378
rect 23480 2314 23532 2320
rect 24872 2332 24952 2360
rect 23492 800 23520 2314
rect 24768 2304 24820 2310
rect 24768 2246 24820 2252
rect 24780 1970 24808 2246
rect 24768 1964 24820 1970
rect 24768 1906 24820 1912
rect 24872 800 24900 2332
rect 24952 2314 25004 2320
rect 25700 2310 25728 4150
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 57152 3664 57204 3670
rect 57152 3606 57204 3612
rect 45192 3596 45244 3602
rect 45192 3538 45244 3544
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35898 2544 35954 2553
rect 35898 2479 35900 2488
rect 35952 2479 35954 2488
rect 35992 2508 36044 2514
rect 35900 2450 35952 2456
rect 35992 2450 36044 2456
rect 25780 2440 25832 2446
rect 35716 2440 35768 2446
rect 25780 2382 25832 2388
rect 35714 2408 35716 2417
rect 35808 2440 35860 2446
rect 35768 2408 35770 2417
rect 25688 2304 25740 2310
rect 25688 2246 25740 2252
rect 25792 1902 25820 2382
rect 26240 2372 26292 2378
rect 26240 2314 26292 2320
rect 26332 2372 26384 2378
rect 26332 2314 26384 2320
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 29184 2372 29236 2378
rect 29184 2314 29236 2320
rect 30012 2372 30064 2378
rect 30012 2314 30064 2320
rect 30840 2372 30892 2378
rect 30840 2314 30892 2320
rect 32036 2372 32088 2378
rect 32036 2314 32088 2320
rect 32588 2372 32640 2378
rect 32588 2314 32640 2320
rect 33416 2372 33468 2378
rect 33416 2314 33468 2320
rect 33508 2372 33560 2378
rect 33508 2314 33560 2320
rect 35164 2372 35216 2378
rect 36004 2417 36032 2450
rect 35808 2382 35860 2388
rect 35990 2408 36046 2417
rect 35714 2343 35770 2352
rect 35164 2314 35216 2320
rect 26252 1902 26280 2314
rect 25780 1896 25832 1902
rect 25780 1838 25832 1844
rect 26240 1896 26292 1902
rect 26240 1838 26292 1844
rect 26344 800 26372 2314
rect 27344 2304 27396 2310
rect 27344 2246 27396 2252
rect 27356 1834 27384 2246
rect 27344 1828 27396 1834
rect 27344 1770 27396 1776
rect 27724 800 27752 2314
rect 29196 800 29224 2314
rect 30024 814 30052 2314
rect 30852 1170 30880 2314
rect 31668 2304 31720 2310
rect 31668 2246 31720 2252
rect 30668 1142 30880 1170
rect 30012 808 30064 814
rect 18328 604 18380 610
rect 18328 546 18380 552
rect 19154 0 19210 800
rect 20626 0 20682 800
rect 22006 0 22062 800
rect 23478 0 23534 800
rect 24858 0 24914 800
rect 26330 0 26386 800
rect 27710 0 27766 800
rect 29182 0 29238 800
rect 30668 800 30696 1142
rect 31680 950 31708 2246
rect 31668 944 31720 950
rect 31668 886 31720 892
rect 32048 800 32076 2314
rect 32600 1018 32628 2314
rect 33428 1873 33456 2314
rect 33414 1864 33470 1873
rect 33414 1799 33470 1808
rect 32588 1012 32640 1018
rect 32588 954 32640 960
rect 33520 800 33548 2314
rect 34900 870 35020 898
rect 34900 800 34928 870
rect 30012 750 30064 756
rect 30654 0 30710 800
rect 32034 0 32090 800
rect 33506 0 33562 800
rect 34886 0 34942 800
rect 34992 762 35020 870
rect 35176 762 35204 2314
rect 35532 2304 35584 2310
rect 35820 2258 35848 2382
rect 35990 2343 36046 2352
rect 37280 2372 37332 2378
rect 37280 2314 37332 2320
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 39212 2372 39264 2378
rect 39212 2314 39264 2320
rect 40592 2372 40644 2378
rect 40592 2314 40644 2320
rect 42064 2372 42116 2378
rect 42064 2314 42116 2320
rect 43444 2372 43496 2378
rect 43444 2314 43496 2320
rect 44916 2372 44968 2378
rect 44916 2314 44968 2320
rect 35532 2246 35584 2252
rect 35544 1290 35572 2246
rect 35636 2230 35848 2258
rect 36360 2304 36412 2310
rect 37292 2281 37320 2314
rect 37648 2304 37700 2310
rect 36360 2246 36412 2252
rect 37278 2272 37334 2281
rect 35636 1902 35664 2230
rect 35624 1896 35676 1902
rect 35624 1838 35676 1844
rect 35806 1864 35862 1873
rect 35806 1799 35808 1808
rect 35860 1799 35862 1808
rect 35808 1770 35860 1776
rect 35532 1284 35584 1290
rect 35532 1226 35584 1232
rect 36372 800 36400 2246
rect 37648 2246 37700 2252
rect 37278 2207 37334 2216
rect 34992 734 35204 762
rect 36358 0 36414 800
rect 37660 746 37688 2246
rect 37752 800 37780 2314
rect 38568 2304 38620 2310
rect 38568 2246 38620 2252
rect 38580 1154 38608 2246
rect 38568 1148 38620 1154
rect 38568 1090 38620 1096
rect 39224 800 39252 2314
rect 40500 2304 40552 2310
rect 40500 2246 40552 2252
rect 40512 1737 40540 2246
rect 40498 1728 40554 1737
rect 40498 1663 40554 1672
rect 40604 800 40632 2314
rect 41144 2304 41196 2310
rect 41144 2246 41196 2252
rect 41156 1086 41184 2246
rect 41144 1080 41196 1086
rect 41144 1022 41196 1028
rect 42076 800 42104 2314
rect 42800 2304 42852 2310
rect 42800 2246 42852 2252
rect 37648 740 37700 746
rect 37648 682 37700 688
rect 37738 0 37794 800
rect 39210 0 39266 800
rect 40590 0 40646 800
rect 42062 0 42118 800
rect 42812 678 42840 2246
rect 43456 800 43484 2314
rect 43904 2304 43956 2310
rect 43904 2246 43956 2252
rect 43916 882 43944 2246
rect 43904 876 43956 882
rect 43904 818 43956 824
rect 44928 800 44956 2314
rect 45204 2310 45232 3538
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 54852 3052 54904 3058
rect 54852 2994 54904 3000
rect 51908 2916 51960 2922
rect 51908 2858 51960 2864
rect 45466 2544 45522 2553
rect 45376 2508 45428 2514
rect 45466 2479 45468 2488
rect 45376 2450 45428 2456
rect 45520 2479 45522 2488
rect 45468 2450 45520 2456
rect 45388 2417 45416 2450
rect 45374 2408 45430 2417
rect 45374 2343 45430 2352
rect 45742 2408 45798 2417
rect 49054 2408 49110 2417
rect 45742 2343 45798 2352
rect 46296 2372 46348 2378
rect 45192 2304 45244 2310
rect 45376 2304 45428 2310
rect 45192 2246 45244 2252
rect 45374 2272 45376 2281
rect 45428 2272 45430 2281
rect 45374 2207 45430 2216
rect 45650 1728 45706 1737
rect 45650 1663 45706 1672
rect 45664 1630 45692 1663
rect 45560 1624 45612 1630
rect 45560 1566 45612 1572
rect 45652 1624 45704 1630
rect 45652 1566 45704 1572
rect 45572 1358 45600 1566
rect 45756 1494 45784 2343
rect 46296 2314 46348 2320
rect 47676 2372 47728 2378
rect 47676 2314 47728 2320
rect 47768 2372 47820 2378
rect 51920 2378 51948 2858
rect 53378 2408 53434 2417
rect 49054 2343 49056 2352
rect 47768 2314 47820 2320
rect 49108 2343 49110 2352
rect 49148 2372 49200 2378
rect 49056 2314 49108 2320
rect 49148 2314 49200 2320
rect 50620 2372 50672 2378
rect 50620 2314 50672 2320
rect 51908 2372 51960 2378
rect 51908 2314 51960 2320
rect 52000 2372 52052 2378
rect 53378 2343 53380 2352
rect 52000 2314 52052 2320
rect 53432 2343 53434 2352
rect 53472 2372 53524 2378
rect 53380 2314 53432 2320
rect 53472 2314 53524 2320
rect 45652 1488 45704 1494
rect 45652 1430 45704 1436
rect 45744 1488 45796 1494
rect 45744 1430 45796 1436
rect 45560 1352 45612 1358
rect 45560 1294 45612 1300
rect 45664 1222 45692 1430
rect 45652 1216 45704 1222
rect 45652 1158 45704 1164
rect 46308 800 46336 2314
rect 47688 1601 47716 2314
rect 47674 1592 47730 1601
rect 47674 1527 47730 1536
rect 47780 800 47808 2314
rect 49160 800 49188 2314
rect 49608 2304 49660 2310
rect 49608 2246 49660 2252
rect 42800 672 42852 678
rect 42800 614 42852 620
rect 43442 0 43498 800
rect 44914 0 44970 800
rect 46294 0 46350 800
rect 47766 0 47822 800
rect 49146 0 49202 800
rect 49620 406 49648 2246
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 50632 800 50660 2314
rect 51080 2100 51132 2106
rect 51080 2042 51132 2048
rect 51092 2009 51120 2042
rect 51356 2032 51408 2038
rect 51078 2000 51134 2009
rect 51356 1974 51408 1980
rect 51078 1935 51134 1944
rect 51078 1864 51134 1873
rect 51078 1799 51134 1808
rect 51092 1562 51120 1799
rect 51170 1728 51226 1737
rect 51170 1663 51226 1672
rect 51080 1556 51132 1562
rect 51080 1498 51132 1504
rect 51184 1494 51212 1663
rect 51262 1592 51318 1601
rect 51262 1527 51264 1536
rect 51316 1527 51318 1536
rect 51264 1498 51316 1504
rect 51172 1488 51224 1494
rect 51368 1442 51396 1974
rect 51172 1430 51224 1436
rect 51276 1426 51396 1442
rect 51632 1488 51684 1494
rect 51632 1430 51684 1436
rect 51264 1420 51396 1426
rect 51316 1414 51396 1420
rect 51264 1362 51316 1368
rect 51644 1222 51672 1430
rect 51632 1216 51684 1222
rect 51632 1158 51684 1164
rect 52012 800 52040 2314
rect 53484 800 53512 2314
rect 54864 800 54892 2994
rect 56692 2916 56744 2922
rect 56692 2858 56744 2864
rect 56508 2848 56560 2854
rect 56508 2790 56560 2796
rect 56140 2644 56192 2650
rect 56140 2586 56192 2592
rect 55864 2576 55916 2582
rect 55770 2544 55826 2553
rect 56048 2576 56100 2582
rect 55916 2524 56048 2530
rect 55864 2518 56100 2524
rect 55876 2502 56088 2518
rect 55770 2479 55772 2488
rect 55824 2479 55826 2488
rect 55772 2450 55824 2456
rect 56152 2310 56180 2586
rect 56520 2394 56548 2790
rect 56704 2689 56732 2858
rect 56690 2680 56746 2689
rect 57164 2650 57192 3606
rect 58268 2650 58296 4218
rect 67364 4140 67416 4146
rect 67364 4082 67416 4088
rect 63132 4072 63184 4078
rect 63132 4014 63184 4020
rect 61660 3732 61712 3738
rect 61660 3674 61712 3680
rect 61384 3120 61436 3126
rect 61384 3062 61436 3068
rect 59176 3052 59228 3058
rect 59176 2994 59228 3000
rect 59544 3052 59596 3058
rect 59544 2994 59596 3000
rect 61016 3052 61068 3058
rect 61016 2994 61068 3000
rect 56690 2615 56746 2624
rect 57152 2644 57204 2650
rect 57152 2586 57204 2592
rect 58256 2644 58308 2650
rect 58256 2586 58308 2592
rect 58440 2644 58492 2650
rect 58440 2586 58492 2592
rect 58452 2553 58480 2586
rect 58438 2544 58494 2553
rect 58438 2479 58494 2488
rect 56336 2366 56548 2394
rect 56692 2372 56744 2378
rect 55680 2304 55732 2310
rect 55678 2272 55680 2281
rect 56140 2304 56192 2310
rect 55732 2272 55734 2281
rect 56140 2246 56192 2252
rect 55678 2207 55734 2216
rect 56336 1358 56364 2366
rect 56692 2314 56744 2320
rect 57704 2372 57756 2378
rect 57704 2314 57756 2320
rect 56704 2122 56732 2314
rect 56520 2094 56732 2122
rect 56324 1352 56376 1358
rect 56324 1294 56376 1300
rect 56520 1034 56548 2094
rect 56336 1006 56548 1034
rect 56336 800 56364 1006
rect 57716 800 57744 2314
rect 59188 800 59216 2994
rect 59556 2378 59584 2994
rect 59818 2816 59874 2825
rect 59818 2751 59874 2760
rect 59634 2408 59690 2417
rect 59544 2372 59596 2378
rect 59634 2343 59690 2352
rect 59544 2314 59596 2320
rect 59648 2310 59676 2343
rect 59636 2304 59688 2310
rect 59728 2304 59780 2310
rect 59636 2246 59688 2252
rect 59726 2272 59728 2281
rect 59780 2272 59782 2281
rect 59726 2207 59782 2216
rect 59832 2038 59860 2751
rect 60278 2544 60334 2553
rect 60278 2479 60280 2488
rect 60332 2479 60334 2488
rect 60648 2508 60700 2514
rect 60280 2450 60332 2456
rect 60832 2508 60884 2514
rect 60648 2450 60700 2456
rect 60752 2468 60832 2496
rect 59912 2440 59964 2446
rect 59912 2382 59964 2388
rect 59820 2032 59872 2038
rect 59924 2009 59952 2382
rect 60188 2372 60240 2378
rect 60660 2360 60688 2450
rect 60188 2314 60240 2320
rect 60568 2332 60688 2360
rect 60200 2281 60228 2314
rect 60186 2272 60242 2281
rect 60186 2207 60242 2216
rect 60188 2100 60240 2106
rect 60188 2042 60240 2048
rect 60372 2100 60424 2106
rect 60372 2042 60424 2048
rect 59820 1974 59872 1980
rect 59910 2000 59966 2009
rect 59910 1935 59966 1944
rect 60200 1873 60228 2042
rect 60384 2009 60412 2042
rect 60370 2000 60426 2009
rect 60370 1935 60426 1944
rect 60186 1864 60242 1873
rect 60186 1799 60242 1808
rect 60568 1737 60596 2332
rect 60752 2281 60780 2468
rect 60832 2450 60884 2456
rect 61028 2378 61056 2994
rect 61108 2848 61160 2854
rect 61108 2790 61160 2796
rect 61016 2372 61068 2378
rect 61016 2314 61068 2320
rect 60738 2272 60794 2281
rect 60738 2207 60794 2216
rect 60740 1896 60792 1902
rect 60924 1896 60976 1902
rect 60792 1844 60924 1850
rect 60740 1838 60976 1844
rect 60752 1822 60964 1838
rect 60554 1728 60610 1737
rect 60554 1663 60610 1672
rect 60568 1562 60872 1578
rect 60556 1556 60872 1562
rect 60608 1550 60872 1556
rect 60556 1498 60608 1504
rect 60464 1488 60516 1494
rect 60844 1476 60872 1550
rect 61016 1488 61068 1494
rect 60464 1430 60516 1436
rect 60738 1456 60794 1465
rect 60476 1329 60504 1430
rect 60844 1448 61016 1476
rect 61016 1430 61068 1436
rect 60738 1391 60740 1400
rect 60792 1391 60794 1400
rect 60740 1362 60792 1368
rect 60462 1320 60518 1329
rect 60462 1255 60518 1264
rect 61120 898 61148 2790
rect 61290 2680 61346 2689
rect 61290 2615 61346 2624
rect 61304 2514 61332 2615
rect 61292 2508 61344 2514
rect 61292 2450 61344 2456
rect 61200 1420 61252 1426
rect 61200 1362 61252 1368
rect 61212 1329 61240 1362
rect 61198 1320 61254 1329
rect 61198 1255 61254 1264
rect 61396 1222 61424 3062
rect 61672 3058 61700 3674
rect 63144 3534 63172 4014
rect 64972 3936 65024 3942
rect 64972 3878 65024 3884
rect 63132 3528 63184 3534
rect 63132 3470 63184 3476
rect 61660 3052 61712 3058
rect 61660 2994 61712 3000
rect 62120 2848 62172 2854
rect 62120 2790 62172 2796
rect 62132 2446 62160 2790
rect 62120 2440 62172 2446
rect 62120 2382 62172 2388
rect 63144 2378 63172 3470
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 63604 3058 63632 3334
rect 63592 3052 63644 3058
rect 63592 2994 63644 3000
rect 64880 3052 64932 3058
rect 64880 2994 64932 3000
rect 64420 2984 64472 2990
rect 64420 2926 64472 2932
rect 63500 2848 63552 2854
rect 63500 2790 63552 2796
rect 63408 2440 63460 2446
rect 63408 2382 63460 2388
rect 63132 2372 63184 2378
rect 63132 2314 63184 2320
rect 63316 2372 63368 2378
rect 63316 2314 63368 2320
rect 61936 2304 61988 2310
rect 61936 2246 61988 2252
rect 62028 2304 62080 2310
rect 62028 2246 62080 2252
rect 61948 2038 61976 2246
rect 61936 2032 61988 2038
rect 61936 1974 61988 1980
rect 61752 1556 61804 1562
rect 61752 1498 61804 1504
rect 61764 1358 61792 1498
rect 61752 1352 61804 1358
rect 61752 1294 61804 1300
rect 61384 1216 61436 1222
rect 61384 1158 61436 1164
rect 60660 870 60780 898
rect 60660 800 60688 870
rect 49608 400 49660 406
rect 49608 342 49660 348
rect 50618 0 50674 800
rect 51998 0 52054 800
rect 53470 0 53526 800
rect 54850 0 54906 800
rect 56322 0 56378 800
rect 57702 0 57758 800
rect 59174 0 59230 800
rect 60646 0 60702 800
rect 60752 762 60780 870
rect 61028 870 61148 898
rect 61028 762 61056 870
rect 62040 800 62068 2246
rect 63328 1698 63356 2314
rect 63420 1873 63448 2382
rect 63406 1864 63462 1873
rect 63406 1799 63462 1808
rect 63316 1692 63368 1698
rect 63316 1634 63368 1640
rect 63512 800 63540 2790
rect 64144 2644 64196 2650
rect 64144 2586 64196 2592
rect 64156 2553 64184 2586
rect 64142 2544 64198 2553
rect 64142 2479 64198 2488
rect 64432 2446 64460 2926
rect 64892 2650 64920 2994
rect 64984 2990 65012 3878
rect 65654 3836 65962 3856
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3760 65962 3780
rect 65524 3460 65576 3466
rect 65524 3402 65576 3408
rect 65536 3194 65564 3402
rect 65524 3188 65576 3194
rect 65524 3130 65576 3136
rect 67376 3058 67404 4082
rect 68836 4004 68888 4010
rect 68836 3946 68888 3952
rect 68848 3534 68876 3946
rect 68284 3528 68336 3534
rect 68284 3470 68336 3476
rect 68836 3528 68888 3534
rect 68836 3470 68888 3476
rect 66720 3052 66772 3058
rect 66720 2994 66772 3000
rect 67364 3052 67416 3058
rect 67364 2994 67416 3000
rect 64972 2984 65024 2990
rect 65524 2984 65576 2990
rect 64972 2926 65024 2932
rect 65246 2952 65302 2961
rect 65524 2926 65576 2932
rect 65246 2887 65302 2896
rect 64972 2848 65024 2854
rect 64972 2790 65024 2796
rect 65154 2816 65210 2825
rect 64880 2644 64932 2650
rect 64880 2586 64932 2592
rect 64420 2440 64472 2446
rect 64420 2382 64472 2388
rect 64984 1442 65012 2790
rect 65154 2751 65210 2760
rect 65168 2650 65196 2751
rect 65260 2650 65288 2887
rect 65156 2644 65208 2650
rect 65156 2586 65208 2592
rect 65248 2644 65300 2650
rect 65248 2586 65300 2592
rect 65168 2310 65196 2586
rect 65536 2446 65564 2926
rect 66168 2916 66220 2922
rect 66168 2858 66220 2864
rect 65654 2748 65962 2768
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2672 65962 2692
rect 65524 2440 65576 2446
rect 65524 2382 65576 2388
rect 65156 2304 65208 2310
rect 65156 2246 65208 2252
rect 66180 1698 66208 2858
rect 66352 2848 66404 2854
rect 66352 2790 66404 2796
rect 66168 1692 66220 1698
rect 66168 1634 66220 1640
rect 64892 1414 65012 1442
rect 64892 800 64920 1414
rect 65524 1352 65576 1358
rect 65524 1294 65576 1300
rect 60752 734 61056 762
rect 62026 0 62082 800
rect 63498 0 63554 800
rect 64878 0 64934 800
rect 65536 406 65564 1294
rect 66364 800 66392 2790
rect 66732 2446 66760 2994
rect 67732 2848 67784 2854
rect 67732 2790 67784 2796
rect 66720 2440 66772 2446
rect 66720 2382 66772 2388
rect 66902 2408 66958 2417
rect 66902 2343 66958 2352
rect 66812 2304 66864 2310
rect 66812 2246 66864 2252
rect 66824 2106 66852 2246
rect 66916 2106 66944 2343
rect 67456 2304 67508 2310
rect 67454 2272 67456 2281
rect 67508 2272 67510 2281
rect 67454 2207 67510 2216
rect 66812 2100 66864 2106
rect 66812 2042 66864 2048
rect 66904 2100 66956 2106
rect 66904 2042 66956 2048
rect 67744 800 67772 2790
rect 68296 2446 68324 3470
rect 69112 3392 69164 3398
rect 69112 3334 69164 3340
rect 69124 3058 69152 3334
rect 70124 3120 70176 3126
rect 70124 3062 70176 3068
rect 69112 3052 69164 3058
rect 69112 2994 69164 3000
rect 70136 2922 70164 3062
rect 71700 3058 71728 7686
rect 73540 3058 73568 8774
rect 71688 3052 71740 3058
rect 73528 3052 73580 3058
rect 71688 2994 71740 3000
rect 73356 3012 73528 3040
rect 70124 2916 70176 2922
rect 70124 2858 70176 2864
rect 69204 2848 69256 2854
rect 69204 2790 69256 2796
rect 69572 2848 69624 2854
rect 69572 2790 69624 2796
rect 70584 2848 70636 2854
rect 70584 2790 70636 2796
rect 68284 2440 68336 2446
rect 68284 2382 68336 2388
rect 69216 800 69244 2790
rect 69584 2446 69612 2790
rect 69572 2440 69624 2446
rect 69572 2382 69624 2388
rect 69664 2440 69716 2446
rect 69664 2382 69716 2388
rect 69676 2145 69704 2382
rect 69756 2372 69808 2378
rect 69756 2314 69808 2320
rect 69662 2136 69718 2145
rect 69662 2071 69718 2080
rect 69768 1465 69796 2314
rect 70306 2000 70362 2009
rect 70306 1935 70362 1944
rect 70214 1728 70270 1737
rect 70320 1698 70348 1935
rect 70214 1663 70216 1672
rect 70268 1663 70270 1672
rect 70308 1692 70360 1698
rect 70216 1634 70268 1640
rect 70308 1634 70360 1640
rect 69754 1456 69810 1465
rect 69754 1391 69810 1400
rect 70596 800 70624 2790
rect 71700 2378 71728 2994
rect 72056 2848 72108 2854
rect 72056 2790 72108 2796
rect 71688 2372 71740 2378
rect 71688 2314 71740 2320
rect 72068 800 72096 2790
rect 72792 2440 72844 2446
rect 72792 2382 72844 2388
rect 72804 1426 72832 2382
rect 73356 2310 73384 3012
rect 73528 2994 73580 3000
rect 73528 2848 73580 2854
rect 73528 2790 73580 2796
rect 73540 2446 73568 2790
rect 74644 2650 74672 9998
rect 76288 3528 76340 3534
rect 76288 3470 76340 3476
rect 76196 3460 76248 3466
rect 76196 3402 76248 3408
rect 74908 3052 74960 3058
rect 74908 2994 74960 3000
rect 74632 2644 74684 2650
rect 74632 2586 74684 2592
rect 74816 2508 74868 2514
rect 74816 2450 74868 2456
rect 73528 2440 73580 2446
rect 74828 2417 74856 2450
rect 73528 2382 73580 2388
rect 74814 2408 74870 2417
rect 73896 2372 73948 2378
rect 74814 2343 74870 2352
rect 73896 2314 73948 2320
rect 73344 2304 73396 2310
rect 73344 2246 73396 2252
rect 73436 2304 73488 2310
rect 73436 2246 73488 2252
rect 72792 1420 72844 1426
rect 72792 1362 72844 1368
rect 72884 1420 72936 1426
rect 72884 1362 72936 1368
rect 65524 400 65576 406
rect 65524 342 65576 348
rect 66350 0 66406 800
rect 67730 0 67786 800
rect 69202 0 69258 800
rect 70582 0 70638 800
rect 72054 0 72110 800
rect 72896 610 72924 1362
rect 73448 800 73476 2246
rect 73908 1698 73936 2314
rect 74448 2304 74500 2310
rect 74446 2272 74448 2281
rect 74500 2272 74502 2281
rect 74446 2207 74502 2216
rect 73986 1728 74042 1737
rect 73896 1692 73948 1698
rect 73986 1663 73988 1672
rect 73896 1634 73948 1640
rect 74040 1663 74042 1672
rect 73988 1634 74040 1640
rect 74920 800 74948 2994
rect 75000 2848 75052 2854
rect 75000 2790 75052 2796
rect 75012 2514 75040 2790
rect 75000 2508 75052 2514
rect 75000 2450 75052 2456
rect 76208 2378 76236 3402
rect 76104 2372 76156 2378
rect 76104 2314 76156 2320
rect 76196 2372 76248 2378
rect 76196 2314 76248 2320
rect 75000 2304 75052 2310
rect 75000 2246 75052 2252
rect 72884 604 72936 610
rect 72884 546 72936 552
rect 73434 0 73490 800
rect 74906 0 74962 800
rect 75012 542 75040 2246
rect 76116 1970 76144 2314
rect 76012 1964 76064 1970
rect 76012 1906 76064 1912
rect 76104 1964 76156 1970
rect 76104 1906 76156 1912
rect 76024 1465 76052 1906
rect 76010 1456 76066 1465
rect 76010 1391 76066 1400
rect 76300 800 76328 3470
rect 76472 3392 76524 3398
rect 76472 3334 76524 3340
rect 76484 2310 76512 3334
rect 76668 3194 76696 11494
rect 78692 3194 78720 12786
rect 79612 3194 79640 13874
rect 81014 13084 81322 13104
rect 81014 13082 81020 13084
rect 81076 13082 81100 13084
rect 81156 13082 81180 13084
rect 81236 13082 81260 13084
rect 81316 13082 81322 13084
rect 81076 13030 81078 13082
rect 81258 13030 81260 13082
rect 81014 13028 81020 13030
rect 81076 13028 81100 13030
rect 81156 13028 81180 13030
rect 81236 13028 81260 13030
rect 81316 13028 81322 13030
rect 81014 13008 81322 13028
rect 81014 11996 81322 12016
rect 81014 11994 81020 11996
rect 81076 11994 81100 11996
rect 81156 11994 81180 11996
rect 81236 11994 81260 11996
rect 81316 11994 81322 11996
rect 81076 11942 81078 11994
rect 81258 11942 81260 11994
rect 81014 11940 81020 11942
rect 81076 11940 81100 11942
rect 81156 11940 81180 11942
rect 81236 11940 81260 11942
rect 81316 11940 81322 11942
rect 81014 11920 81322 11940
rect 81014 10908 81322 10928
rect 81014 10906 81020 10908
rect 81076 10906 81100 10908
rect 81156 10906 81180 10908
rect 81236 10906 81260 10908
rect 81316 10906 81322 10908
rect 81076 10854 81078 10906
rect 81258 10854 81260 10906
rect 81014 10852 81020 10854
rect 81076 10852 81100 10854
rect 81156 10852 81180 10854
rect 81236 10852 81260 10854
rect 81316 10852 81322 10854
rect 81014 10832 81322 10852
rect 81014 9820 81322 9840
rect 81014 9818 81020 9820
rect 81076 9818 81100 9820
rect 81156 9818 81180 9820
rect 81236 9818 81260 9820
rect 81316 9818 81322 9820
rect 81076 9766 81078 9818
rect 81258 9766 81260 9818
rect 81014 9764 81020 9766
rect 81076 9764 81100 9766
rect 81156 9764 81180 9766
rect 81236 9764 81260 9766
rect 81316 9764 81322 9766
rect 81014 9744 81322 9764
rect 81014 8732 81322 8752
rect 81014 8730 81020 8732
rect 81076 8730 81100 8732
rect 81156 8730 81180 8732
rect 81236 8730 81260 8732
rect 81316 8730 81322 8732
rect 81076 8678 81078 8730
rect 81258 8678 81260 8730
rect 81014 8676 81020 8678
rect 81076 8676 81100 8678
rect 81156 8676 81180 8678
rect 81236 8676 81260 8678
rect 81316 8676 81322 8678
rect 81014 8656 81322 8676
rect 81014 7644 81322 7664
rect 81014 7642 81020 7644
rect 81076 7642 81100 7644
rect 81156 7642 81180 7644
rect 81236 7642 81260 7644
rect 81316 7642 81322 7644
rect 81076 7590 81078 7642
rect 81258 7590 81260 7642
rect 81014 7588 81020 7590
rect 81076 7588 81100 7590
rect 81156 7588 81180 7590
rect 81236 7588 81260 7590
rect 81316 7588 81322 7590
rect 81014 7568 81322 7588
rect 81014 6556 81322 6576
rect 81014 6554 81020 6556
rect 81076 6554 81100 6556
rect 81156 6554 81180 6556
rect 81236 6554 81260 6556
rect 81316 6554 81322 6556
rect 81076 6502 81078 6554
rect 81258 6502 81260 6554
rect 81014 6500 81020 6502
rect 81076 6500 81100 6502
rect 81156 6500 81180 6502
rect 81236 6500 81260 6502
rect 81316 6500 81322 6502
rect 81014 6480 81322 6500
rect 81014 5468 81322 5488
rect 81014 5466 81020 5468
rect 81076 5466 81100 5468
rect 81156 5466 81180 5468
rect 81236 5466 81260 5468
rect 81316 5466 81322 5468
rect 81076 5414 81078 5466
rect 81258 5414 81260 5466
rect 81014 5412 81020 5414
rect 81076 5412 81100 5414
rect 81156 5412 81180 5414
rect 81236 5412 81260 5414
rect 81316 5412 81322 5414
rect 81014 5392 81322 5412
rect 81014 4380 81322 4400
rect 81014 4378 81020 4380
rect 81076 4378 81100 4380
rect 81156 4378 81180 4380
rect 81236 4378 81260 4380
rect 81316 4378 81322 4380
rect 81076 4326 81078 4378
rect 81258 4326 81260 4378
rect 81014 4324 81020 4326
rect 81076 4324 81100 4326
rect 81156 4324 81180 4326
rect 81236 4324 81260 4326
rect 81316 4324 81322 4326
rect 81014 4304 81322 4324
rect 81014 3292 81322 3312
rect 81014 3290 81020 3292
rect 81076 3290 81100 3292
rect 81156 3290 81180 3292
rect 81236 3290 81260 3292
rect 81316 3290 81322 3292
rect 81076 3238 81078 3290
rect 81258 3238 81260 3290
rect 81014 3236 81020 3238
rect 81076 3236 81100 3238
rect 81156 3236 81180 3238
rect 81236 3236 81260 3238
rect 81316 3236 81322 3238
rect 81014 3216 81322 3236
rect 81728 3194 81756 14350
rect 81992 3528 82044 3534
rect 81992 3470 82044 3476
rect 76656 3188 76708 3194
rect 76656 3130 76708 3136
rect 78680 3188 78732 3194
rect 78680 3130 78732 3136
rect 79600 3188 79652 3194
rect 79600 3130 79652 3136
rect 81716 3188 81768 3194
rect 81716 3130 81768 3136
rect 76564 3052 76616 3058
rect 76564 2994 76616 3000
rect 77760 3052 77812 3058
rect 77760 2994 77812 3000
rect 78588 3052 78640 3058
rect 78588 2994 78640 3000
rect 79508 3052 79560 3058
rect 79508 2994 79560 3000
rect 80612 3052 80664 3058
rect 80612 2994 80664 3000
rect 81624 3052 81676 3058
rect 81624 2994 81676 3000
rect 76576 2650 76604 2994
rect 77668 2848 77720 2854
rect 77668 2790 77720 2796
rect 76564 2644 76616 2650
rect 76564 2586 76616 2592
rect 77680 2310 77708 2790
rect 76472 2304 76524 2310
rect 76472 2246 76524 2252
rect 77576 2304 77628 2310
rect 77576 2246 77628 2252
rect 77668 2304 77720 2310
rect 77668 2246 77720 2252
rect 77588 1426 77616 2246
rect 77666 1456 77722 1465
rect 77576 1420 77628 1426
rect 77666 1391 77668 1400
rect 77576 1362 77628 1368
rect 77720 1391 77722 1400
rect 77668 1362 77720 1368
rect 77772 800 77800 2994
rect 78600 2650 78628 2994
rect 79520 2650 79548 2994
rect 78588 2644 78640 2650
rect 78588 2586 78640 2592
rect 79508 2644 79560 2650
rect 79508 2586 79560 2592
rect 79600 2644 79652 2650
rect 79600 2586 79652 2592
rect 79612 2530 79640 2586
rect 79244 2514 79640 2530
rect 79232 2508 79640 2514
rect 79284 2502 79640 2508
rect 79232 2450 79284 2456
rect 79416 2440 79468 2446
rect 79416 2382 79468 2388
rect 79048 2304 79100 2310
rect 79048 2246 79100 2252
rect 79060 1766 79088 2246
rect 79324 1896 79376 1902
rect 79152 1844 79324 1850
rect 79152 1838 79376 1844
rect 79152 1834 79364 1838
rect 79140 1828 79364 1834
rect 79192 1822 79364 1828
rect 79140 1770 79192 1776
rect 79048 1760 79100 1766
rect 79048 1702 79100 1708
rect 79152 870 79272 898
rect 79152 800 79180 870
rect 75000 536 75052 542
rect 75000 478 75052 484
rect 76286 0 76342 800
rect 77758 0 77814 800
rect 79138 0 79194 800
rect 79244 762 79272 870
rect 79428 762 79456 2382
rect 80520 2304 80572 2310
rect 79506 2272 79562 2281
rect 80520 2246 80572 2252
rect 79506 2207 79562 2216
rect 79520 1902 79548 2207
rect 80532 1970 80560 2246
rect 80520 1964 80572 1970
rect 80520 1906 80572 1912
rect 79508 1896 79560 1902
rect 79508 1838 79560 1844
rect 80624 800 80652 2994
rect 81532 2848 81584 2854
rect 81532 2790 81584 2796
rect 80888 2644 80940 2650
rect 80888 2586 80940 2592
rect 80900 1970 80928 2586
rect 81544 2514 81572 2790
rect 81636 2650 81664 2994
rect 81624 2644 81676 2650
rect 81624 2586 81676 2592
rect 81532 2508 81584 2514
rect 81532 2450 81584 2456
rect 81440 2440 81492 2446
rect 81438 2408 81440 2417
rect 81492 2408 81494 2417
rect 81438 2343 81494 2352
rect 81014 2204 81322 2224
rect 81014 2202 81020 2204
rect 81076 2202 81100 2204
rect 81156 2202 81180 2204
rect 81236 2202 81260 2204
rect 81316 2202 81322 2204
rect 81076 2150 81078 2202
rect 81258 2150 81260 2202
rect 81014 2148 81020 2150
rect 81076 2148 81100 2150
rect 81156 2148 81180 2150
rect 81236 2148 81260 2150
rect 81316 2148 81322 2150
rect 81014 2128 81322 2148
rect 80888 1964 80940 1970
rect 80888 1906 80940 1912
rect 82004 800 82032 3470
rect 82832 3194 82860 15438
rect 85028 4208 85080 4214
rect 85028 4150 85080 4156
rect 83464 3528 83516 3534
rect 83464 3470 83516 3476
rect 84844 3528 84896 3534
rect 84844 3470 84896 3476
rect 83096 3392 83148 3398
rect 83096 3334 83148 3340
rect 82820 3188 82872 3194
rect 82820 3130 82872 3136
rect 82544 3052 82596 3058
rect 82544 2994 82596 3000
rect 82556 2650 82584 2994
rect 82544 2644 82596 2650
rect 82544 2586 82596 2592
rect 83108 2310 83136 3334
rect 83096 2304 83148 2310
rect 83096 2246 83148 2252
rect 83476 800 83504 3470
rect 83556 3392 83608 3398
rect 83556 3334 83608 3340
rect 83568 2514 83596 3334
rect 83740 3052 83792 3058
rect 83740 2994 83792 3000
rect 83752 2650 83780 2994
rect 83740 2644 83792 2650
rect 83740 2586 83792 2592
rect 83556 2508 83608 2514
rect 83556 2450 83608 2456
rect 84120 2378 84332 2394
rect 84108 2372 84344 2378
rect 84160 2366 84292 2372
rect 84108 2314 84160 2320
rect 84292 2314 84344 2320
rect 84016 2304 84068 2310
rect 84016 2246 84068 2252
rect 84028 1426 84056 2246
rect 84752 1964 84804 1970
rect 84752 1906 84804 1912
rect 84764 1426 84792 1906
rect 84016 1420 84068 1426
rect 84016 1362 84068 1368
rect 84752 1420 84804 1426
rect 84752 1362 84804 1368
rect 84856 800 84884 3470
rect 84936 3392 84988 3398
rect 84936 3334 84988 3340
rect 84948 2514 84976 3334
rect 84936 2508 84988 2514
rect 84936 2450 84988 2456
rect 85040 2446 85068 4150
rect 85224 3194 85252 17614
rect 86316 3528 86368 3534
rect 86316 3470 86368 3476
rect 85212 3188 85264 3194
rect 85212 3130 85264 3136
rect 85120 3052 85172 3058
rect 85120 2994 85172 3000
rect 85132 2650 85160 2994
rect 85120 2644 85172 2650
rect 85120 2586 85172 2592
rect 85580 2508 85632 2514
rect 85580 2450 85632 2456
rect 85028 2440 85080 2446
rect 85028 2382 85080 2388
rect 85592 2310 85620 2450
rect 85580 2304 85632 2310
rect 85580 2246 85632 2252
rect 86328 800 86356 3470
rect 86408 3392 86460 3398
rect 86408 3334 86460 3340
rect 86420 2514 86448 3334
rect 86696 3194 86724 18022
rect 89456 12986 89484 20402
rect 89444 12980 89496 12986
rect 89444 12922 89496 12928
rect 88800 12844 88852 12850
rect 88800 12786 88852 12792
rect 88340 6316 88392 6322
rect 88340 6258 88392 6264
rect 87696 3528 87748 3534
rect 87696 3470 87748 3476
rect 86684 3188 86736 3194
rect 86684 3130 86736 3136
rect 86592 3052 86644 3058
rect 86592 2994 86644 3000
rect 86604 2650 86632 2994
rect 86868 2848 86920 2854
rect 86868 2790 86920 2796
rect 86592 2644 86644 2650
rect 86592 2586 86644 2592
rect 86880 2514 86908 2790
rect 86408 2508 86460 2514
rect 86408 2450 86460 2456
rect 86868 2508 86920 2514
rect 86868 2450 86920 2456
rect 86592 2304 86644 2310
rect 86592 2246 86644 2252
rect 86604 1766 86632 2246
rect 86592 1760 86644 1766
rect 86592 1702 86644 1708
rect 87708 800 87736 3470
rect 87788 3392 87840 3398
rect 87788 3334 87840 3340
rect 87800 2514 87828 3334
rect 88352 2650 88380 6258
rect 88812 2650 88840 12786
rect 91020 6458 91048 20878
rect 91008 6452 91060 6458
rect 91008 6394 91060 6400
rect 90824 6316 90876 6322
rect 90824 6258 90876 6264
rect 88892 3460 88944 3466
rect 88892 3402 88944 3408
rect 88904 3126 88932 3402
rect 88892 3120 88944 3126
rect 88892 3062 88944 3068
rect 89168 3052 89220 3058
rect 89168 2994 89220 3000
rect 90640 3052 90692 3058
rect 90640 2994 90692 3000
rect 88340 2644 88392 2650
rect 88340 2586 88392 2592
rect 88800 2644 88852 2650
rect 88800 2586 88852 2592
rect 87788 2508 87840 2514
rect 87788 2450 87840 2456
rect 87880 2304 87932 2310
rect 87880 2246 87932 2252
rect 88340 2304 88392 2310
rect 88340 2246 88392 2252
rect 87892 1834 87920 2246
rect 87880 1828 87932 1834
rect 87880 1770 87932 1776
rect 88352 814 88380 2246
rect 88340 808 88392 814
rect 79244 734 79456 762
rect 80610 0 80666 800
rect 81990 0 82046 800
rect 83462 0 83518 800
rect 84842 0 84898 800
rect 86314 0 86370 800
rect 87694 0 87750 800
rect 89180 800 89208 2994
rect 89444 2984 89496 2990
rect 89444 2926 89496 2932
rect 89260 2848 89312 2854
rect 89260 2790 89312 2796
rect 89272 2514 89300 2790
rect 89260 2508 89312 2514
rect 89260 2450 89312 2456
rect 89456 2446 89484 2926
rect 90548 2848 90600 2854
rect 90548 2790 90600 2796
rect 90560 2514 90588 2790
rect 90548 2508 90600 2514
rect 90548 2450 90600 2456
rect 89444 2440 89496 2446
rect 89444 2382 89496 2388
rect 90456 2304 90508 2310
rect 90456 2246 90508 2252
rect 90468 950 90496 2246
rect 90456 944 90508 950
rect 90456 886 90508 892
rect 90652 800 90680 2994
rect 90836 2650 90864 6258
rect 92020 3528 92072 3534
rect 92020 3470 92072 3476
rect 92204 3528 92256 3534
rect 92204 3470 92256 3476
rect 91560 3392 91612 3398
rect 91560 3334 91612 3340
rect 91468 3052 91520 3058
rect 91468 2994 91520 3000
rect 91480 2854 91508 2994
rect 91468 2848 91520 2854
rect 91468 2790 91520 2796
rect 90824 2644 90876 2650
rect 90824 2586 90876 2592
rect 91480 1902 91508 2790
rect 91572 2514 91600 3334
rect 91560 2508 91612 2514
rect 91560 2450 91612 2456
rect 91928 2304 91980 2310
rect 91928 2246 91980 2252
rect 91468 1896 91520 1902
rect 91468 1838 91520 1844
rect 91940 1018 91968 2246
rect 91928 1012 91980 1018
rect 91928 954 91980 960
rect 92032 800 92060 3470
rect 92216 2650 92244 3470
rect 92400 3398 92428 21830
rect 92388 3392 92440 3398
rect 92388 3334 92440 3340
rect 92572 3188 92624 3194
rect 92624 3148 92704 3176
rect 92572 3130 92624 3136
rect 92676 3058 92704 3148
rect 92572 3052 92624 3058
rect 92572 2994 92624 3000
rect 92664 3052 92716 3058
rect 92664 2994 92716 3000
rect 92296 2984 92348 2990
rect 92296 2926 92348 2932
rect 92584 2938 92612 2994
rect 92848 2984 92900 2990
rect 92584 2932 92848 2938
rect 92584 2926 92900 2932
rect 92204 2644 92256 2650
rect 92204 2586 92256 2592
rect 92308 2514 92336 2926
rect 92584 2910 92888 2926
rect 92940 2848 92992 2854
rect 92940 2790 92992 2796
rect 92296 2508 92348 2514
rect 92296 2450 92348 2456
rect 92952 2446 92980 2790
rect 93136 2650 93164 23054
rect 95988 3194 96016 23666
rect 96374 23420 96682 23440
rect 96374 23418 96380 23420
rect 96436 23418 96460 23420
rect 96516 23418 96540 23420
rect 96596 23418 96620 23420
rect 96676 23418 96682 23420
rect 96436 23366 96438 23418
rect 96618 23366 96620 23418
rect 96374 23364 96380 23366
rect 96436 23364 96460 23366
rect 96516 23364 96540 23366
rect 96596 23364 96620 23366
rect 96676 23364 96682 23366
rect 96374 23344 96682 23364
rect 96374 22332 96682 22352
rect 96374 22330 96380 22332
rect 96436 22330 96460 22332
rect 96516 22330 96540 22332
rect 96596 22330 96620 22332
rect 96676 22330 96682 22332
rect 96436 22278 96438 22330
rect 96618 22278 96620 22330
rect 96374 22276 96380 22278
rect 96436 22276 96460 22278
rect 96516 22276 96540 22278
rect 96596 22276 96620 22278
rect 96676 22276 96682 22278
rect 96374 22256 96682 22276
rect 96374 21244 96682 21264
rect 96374 21242 96380 21244
rect 96436 21242 96460 21244
rect 96516 21242 96540 21244
rect 96596 21242 96620 21244
rect 96676 21242 96682 21244
rect 96436 21190 96438 21242
rect 96618 21190 96620 21242
rect 96374 21188 96380 21190
rect 96436 21188 96460 21190
rect 96516 21188 96540 21190
rect 96596 21188 96620 21190
rect 96676 21188 96682 21190
rect 96374 21168 96682 21188
rect 96374 20156 96682 20176
rect 96374 20154 96380 20156
rect 96436 20154 96460 20156
rect 96516 20154 96540 20156
rect 96596 20154 96620 20156
rect 96676 20154 96682 20156
rect 96436 20102 96438 20154
rect 96618 20102 96620 20154
rect 96374 20100 96380 20102
rect 96436 20100 96460 20102
rect 96516 20100 96540 20102
rect 96596 20100 96620 20102
rect 96676 20100 96682 20102
rect 96374 20080 96682 20100
rect 96374 19068 96682 19088
rect 96374 19066 96380 19068
rect 96436 19066 96460 19068
rect 96516 19066 96540 19068
rect 96596 19066 96620 19068
rect 96676 19066 96682 19068
rect 96436 19014 96438 19066
rect 96618 19014 96620 19066
rect 96374 19012 96380 19014
rect 96436 19012 96460 19014
rect 96516 19012 96540 19014
rect 96596 19012 96620 19014
rect 96676 19012 96682 19014
rect 96374 18992 96682 19012
rect 96374 17980 96682 18000
rect 96374 17978 96380 17980
rect 96436 17978 96460 17980
rect 96516 17978 96540 17980
rect 96596 17978 96620 17980
rect 96676 17978 96682 17980
rect 96436 17926 96438 17978
rect 96618 17926 96620 17978
rect 96374 17924 96380 17926
rect 96436 17924 96460 17926
rect 96516 17924 96540 17926
rect 96596 17924 96620 17926
rect 96676 17924 96682 17926
rect 96374 17904 96682 17924
rect 96374 16892 96682 16912
rect 96374 16890 96380 16892
rect 96436 16890 96460 16892
rect 96516 16890 96540 16892
rect 96596 16890 96620 16892
rect 96676 16890 96682 16892
rect 96436 16838 96438 16890
rect 96618 16838 96620 16890
rect 96374 16836 96380 16838
rect 96436 16836 96460 16838
rect 96516 16836 96540 16838
rect 96596 16836 96620 16838
rect 96676 16836 96682 16838
rect 96374 16816 96682 16836
rect 96374 15804 96682 15824
rect 96374 15802 96380 15804
rect 96436 15802 96460 15804
rect 96516 15802 96540 15804
rect 96596 15802 96620 15804
rect 96676 15802 96682 15804
rect 96436 15750 96438 15802
rect 96618 15750 96620 15802
rect 96374 15748 96380 15750
rect 96436 15748 96460 15750
rect 96516 15748 96540 15750
rect 96596 15748 96620 15750
rect 96676 15748 96682 15750
rect 96374 15728 96682 15748
rect 96374 14716 96682 14736
rect 96374 14714 96380 14716
rect 96436 14714 96460 14716
rect 96516 14714 96540 14716
rect 96596 14714 96620 14716
rect 96676 14714 96682 14716
rect 96436 14662 96438 14714
rect 96618 14662 96620 14714
rect 96374 14660 96380 14662
rect 96436 14660 96460 14662
rect 96516 14660 96540 14662
rect 96596 14660 96620 14662
rect 96676 14660 96682 14662
rect 96374 14640 96682 14660
rect 96374 13628 96682 13648
rect 96374 13626 96380 13628
rect 96436 13626 96460 13628
rect 96516 13626 96540 13628
rect 96596 13626 96620 13628
rect 96676 13626 96682 13628
rect 96436 13574 96438 13626
rect 96618 13574 96620 13626
rect 96374 13572 96380 13574
rect 96436 13572 96460 13574
rect 96516 13572 96540 13574
rect 96596 13572 96620 13574
rect 96676 13572 96682 13574
rect 96374 13552 96682 13572
rect 96374 12540 96682 12560
rect 96374 12538 96380 12540
rect 96436 12538 96460 12540
rect 96516 12538 96540 12540
rect 96596 12538 96620 12540
rect 96676 12538 96682 12540
rect 96436 12486 96438 12538
rect 96618 12486 96620 12538
rect 96374 12484 96380 12486
rect 96436 12484 96460 12486
rect 96516 12484 96540 12486
rect 96596 12484 96620 12486
rect 96676 12484 96682 12486
rect 96374 12464 96682 12484
rect 96374 11452 96682 11472
rect 96374 11450 96380 11452
rect 96436 11450 96460 11452
rect 96516 11450 96540 11452
rect 96596 11450 96620 11452
rect 96676 11450 96682 11452
rect 96436 11398 96438 11450
rect 96618 11398 96620 11450
rect 96374 11396 96380 11398
rect 96436 11396 96460 11398
rect 96516 11396 96540 11398
rect 96596 11396 96620 11398
rect 96676 11396 96682 11398
rect 96374 11376 96682 11396
rect 96374 10364 96682 10384
rect 96374 10362 96380 10364
rect 96436 10362 96460 10364
rect 96516 10362 96540 10364
rect 96596 10362 96620 10364
rect 96676 10362 96682 10364
rect 96436 10310 96438 10362
rect 96618 10310 96620 10362
rect 96374 10308 96380 10310
rect 96436 10308 96460 10310
rect 96516 10308 96540 10310
rect 96596 10308 96620 10310
rect 96676 10308 96682 10310
rect 96374 10288 96682 10308
rect 96374 9276 96682 9296
rect 96374 9274 96380 9276
rect 96436 9274 96460 9276
rect 96516 9274 96540 9276
rect 96596 9274 96620 9276
rect 96676 9274 96682 9276
rect 96436 9222 96438 9274
rect 96618 9222 96620 9274
rect 96374 9220 96380 9222
rect 96436 9220 96460 9222
rect 96516 9220 96540 9222
rect 96596 9220 96620 9222
rect 96676 9220 96682 9222
rect 96374 9200 96682 9220
rect 96374 8188 96682 8208
rect 96374 8186 96380 8188
rect 96436 8186 96460 8188
rect 96516 8186 96540 8188
rect 96596 8186 96620 8188
rect 96676 8186 96682 8188
rect 96436 8134 96438 8186
rect 96618 8134 96620 8186
rect 96374 8132 96380 8134
rect 96436 8132 96460 8134
rect 96516 8132 96540 8134
rect 96596 8132 96620 8134
rect 96676 8132 96682 8134
rect 96374 8112 96682 8132
rect 96374 7100 96682 7120
rect 96374 7098 96380 7100
rect 96436 7098 96460 7100
rect 96516 7098 96540 7100
rect 96596 7098 96620 7100
rect 96676 7098 96682 7100
rect 96436 7046 96438 7098
rect 96618 7046 96620 7098
rect 96374 7044 96380 7046
rect 96436 7044 96460 7046
rect 96516 7044 96540 7046
rect 96596 7044 96620 7046
rect 96676 7044 96682 7046
rect 96374 7024 96682 7044
rect 96374 6012 96682 6032
rect 96374 6010 96380 6012
rect 96436 6010 96460 6012
rect 96516 6010 96540 6012
rect 96596 6010 96620 6012
rect 96676 6010 96682 6012
rect 96436 5958 96438 6010
rect 96618 5958 96620 6010
rect 96374 5956 96380 5958
rect 96436 5956 96460 5958
rect 96516 5956 96540 5958
rect 96596 5956 96620 5958
rect 96676 5956 96682 5958
rect 96374 5936 96682 5956
rect 96374 4924 96682 4944
rect 96374 4922 96380 4924
rect 96436 4922 96460 4924
rect 96516 4922 96540 4924
rect 96596 4922 96620 4924
rect 96676 4922 96682 4924
rect 96436 4870 96438 4922
rect 96618 4870 96620 4922
rect 96374 4868 96380 4870
rect 96436 4868 96460 4870
rect 96516 4868 96540 4870
rect 96596 4868 96620 4870
rect 96676 4868 96682 4870
rect 96374 4848 96682 4868
rect 96374 3836 96682 3856
rect 96374 3834 96380 3836
rect 96436 3834 96460 3836
rect 96516 3834 96540 3836
rect 96596 3834 96620 3836
rect 96676 3834 96682 3836
rect 96436 3782 96438 3834
rect 96618 3782 96620 3834
rect 96374 3780 96380 3782
rect 96436 3780 96460 3782
rect 96516 3780 96540 3782
rect 96596 3780 96620 3782
rect 96676 3780 96682 3782
rect 96374 3760 96682 3780
rect 96160 3528 96212 3534
rect 96160 3470 96212 3476
rect 93952 3188 94004 3194
rect 93952 3130 94004 3136
rect 95976 3188 96028 3194
rect 95976 3130 96028 3136
rect 93964 2650 93992 3130
rect 94872 3052 94924 3058
rect 94872 2994 94924 3000
rect 95792 3052 95844 3058
rect 95792 2994 95844 3000
rect 93124 2644 93176 2650
rect 93124 2586 93176 2592
rect 93952 2644 94004 2650
rect 93952 2586 94004 2592
rect 92940 2440 92992 2446
rect 92940 2382 92992 2388
rect 93492 2440 93544 2446
rect 93492 2382 93544 2388
rect 93504 800 93532 2382
rect 94884 800 94912 2994
rect 95516 2848 95568 2854
rect 95516 2790 95568 2796
rect 95528 2514 95556 2790
rect 95804 2650 95832 2994
rect 95792 2644 95844 2650
rect 95792 2586 95844 2592
rect 95516 2508 95568 2514
rect 95516 2450 95568 2456
rect 95424 2304 95476 2310
rect 95424 2246 95476 2252
rect 95436 1290 95464 2246
rect 96172 1850 96200 3470
rect 96908 3194 96936 24754
rect 97540 4480 97592 4486
rect 97540 4422 97592 4428
rect 97552 4282 97580 4422
rect 97540 4276 97592 4282
rect 97540 4218 97592 4224
rect 98000 4276 98052 4282
rect 98000 4218 98052 4224
rect 97908 4140 97960 4146
rect 97908 4082 97960 4088
rect 97724 3528 97776 3534
rect 97724 3470 97776 3476
rect 97632 3460 97684 3466
rect 97632 3402 97684 3408
rect 96988 3392 97040 3398
rect 96988 3334 97040 3340
rect 96896 3188 96948 3194
rect 96896 3130 96948 3136
rect 96252 3052 96304 3058
rect 96252 2994 96304 3000
rect 96264 2650 96292 2994
rect 96374 2748 96682 2768
rect 96374 2746 96380 2748
rect 96436 2746 96460 2748
rect 96516 2746 96540 2748
rect 96596 2746 96620 2748
rect 96676 2746 96682 2748
rect 96436 2694 96438 2746
rect 96618 2694 96620 2746
rect 96374 2692 96380 2694
rect 96436 2692 96460 2694
rect 96516 2692 96540 2694
rect 96596 2692 96620 2694
rect 96676 2692 96682 2694
rect 96374 2672 96682 2692
rect 96252 2644 96304 2650
rect 96252 2586 96304 2592
rect 97000 2514 97028 3334
rect 97644 3097 97672 3402
rect 97630 3088 97686 3097
rect 97630 3023 97632 3032
rect 97684 3023 97686 3032
rect 97632 2994 97684 3000
rect 97736 2582 97764 3470
rect 97920 2938 97948 4082
rect 97828 2910 97948 2938
rect 97540 2576 97592 2582
rect 97540 2518 97592 2524
rect 97724 2576 97776 2582
rect 97724 2518 97776 2524
rect 96988 2508 97040 2514
rect 96988 2450 97040 2456
rect 97552 2417 97580 2518
rect 97538 2408 97594 2417
rect 97538 2343 97594 2352
rect 96896 2304 96948 2310
rect 96896 2246 96948 2252
rect 96172 1822 96384 1850
rect 95424 1284 95476 1290
rect 95424 1226 95476 1232
rect 96356 800 96384 1822
rect 88340 750 88392 756
rect 89166 0 89222 800
rect 90638 0 90694 800
rect 92018 0 92074 800
rect 93490 0 93546 800
rect 94870 0 94926 800
rect 96342 0 96398 800
rect 96908 746 96936 2246
rect 97828 2122 97856 2910
rect 97908 2848 97960 2854
rect 97908 2790 97960 2796
rect 97920 2650 97948 2790
rect 97908 2644 97960 2650
rect 97908 2586 97960 2592
rect 98012 2514 98040 4218
rect 98104 3398 98132 25842
rect 98932 3670 98960 36722
rect 111734 35932 112042 35952
rect 111734 35930 111740 35932
rect 111796 35930 111820 35932
rect 111876 35930 111900 35932
rect 111956 35930 111980 35932
rect 112036 35930 112042 35932
rect 111796 35878 111798 35930
rect 111978 35878 111980 35930
rect 111734 35876 111740 35878
rect 111796 35876 111820 35878
rect 111876 35876 111900 35878
rect 111956 35876 111980 35878
rect 112036 35876 112042 35878
rect 111734 35856 112042 35876
rect 111734 34844 112042 34864
rect 111734 34842 111740 34844
rect 111796 34842 111820 34844
rect 111876 34842 111900 34844
rect 111956 34842 111980 34844
rect 112036 34842 112042 34844
rect 111796 34790 111798 34842
rect 111978 34790 111980 34842
rect 111734 34788 111740 34790
rect 111796 34788 111820 34790
rect 111876 34788 111900 34790
rect 111956 34788 111980 34790
rect 112036 34788 112042 34790
rect 111734 34768 112042 34788
rect 112168 33992 112220 33998
rect 112168 33934 112220 33940
rect 111734 33756 112042 33776
rect 111734 33754 111740 33756
rect 111796 33754 111820 33756
rect 111876 33754 111900 33756
rect 111956 33754 111980 33756
rect 112036 33754 112042 33756
rect 111796 33702 111798 33754
rect 111978 33702 111980 33754
rect 111734 33700 111740 33702
rect 111796 33700 111820 33702
rect 111876 33700 111900 33702
rect 111956 33700 111980 33702
rect 112036 33700 112042 33702
rect 111734 33680 112042 33700
rect 110788 33516 110840 33522
rect 110788 33458 110840 33464
rect 108488 32428 108540 32434
rect 108488 32370 108540 32376
rect 107108 31340 107160 31346
rect 107108 31282 107160 31288
rect 106004 30252 106056 30258
rect 106004 30194 106056 30200
rect 104440 29640 104492 29646
rect 104440 29582 104492 29588
rect 102416 28552 102468 28558
rect 102416 28494 102468 28500
rect 100576 27464 100628 27470
rect 100576 27406 100628 27412
rect 99840 26988 99892 26994
rect 99840 26930 99892 26936
rect 98644 3664 98696 3670
rect 98644 3606 98696 3612
rect 98920 3664 98972 3670
rect 98920 3606 98972 3612
rect 98656 3534 98684 3606
rect 98736 3596 98788 3602
rect 98736 3538 98788 3544
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 98092 3392 98144 3398
rect 98092 3334 98144 3340
rect 98644 3052 98696 3058
rect 98644 2994 98696 3000
rect 98656 2854 98684 2994
rect 98460 2848 98512 2854
rect 98460 2790 98512 2796
rect 98644 2848 98696 2854
rect 98644 2790 98696 2796
rect 98472 2689 98500 2790
rect 98458 2680 98514 2689
rect 98458 2615 98514 2624
rect 98000 2508 98052 2514
rect 98000 2450 98052 2456
rect 98092 2304 98144 2310
rect 98092 2246 98144 2252
rect 97736 2094 97856 2122
rect 97736 800 97764 2094
rect 98104 1154 98132 2246
rect 98472 1426 98500 2615
rect 98748 2553 98776 3538
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99104 3460 99156 3466
rect 99104 3402 99156 3408
rect 99116 2582 99144 3402
rect 99300 3194 99328 3470
rect 99564 3460 99616 3466
rect 99564 3402 99616 3408
rect 99288 3188 99340 3194
rect 99288 3130 99340 3136
rect 99472 3052 99524 3058
rect 99472 2994 99524 3000
rect 99104 2576 99156 2582
rect 98734 2544 98790 2553
rect 99484 2530 99512 2994
rect 99576 2990 99604 3402
rect 99852 3398 99880 26930
rect 100392 4276 100444 4282
rect 100392 4218 100444 4224
rect 100300 3528 100352 3534
rect 100300 3470 100352 3476
rect 99840 3392 99892 3398
rect 99840 3334 99892 3340
rect 99654 3224 99710 3233
rect 99654 3159 99710 3168
rect 99668 3126 99696 3159
rect 99656 3120 99708 3126
rect 99656 3062 99708 3068
rect 99564 2984 99616 2990
rect 99564 2926 99616 2932
rect 99748 2984 99800 2990
rect 99748 2926 99800 2932
rect 99562 2680 99618 2689
rect 99562 2615 99618 2624
rect 99576 2582 99604 2615
rect 99760 2582 99788 2926
rect 100312 2650 100340 3470
rect 100300 2644 100352 2650
rect 100300 2586 100352 2592
rect 99104 2518 99156 2524
rect 98734 2479 98790 2488
rect 99392 2502 99512 2530
rect 99564 2576 99616 2582
rect 99564 2518 99616 2524
rect 99748 2576 99800 2582
rect 99748 2518 99800 2524
rect 100404 2514 100432 4218
rect 100588 3398 100616 27406
rect 100852 4140 100904 4146
rect 100852 4082 100904 4088
rect 100864 4026 100892 4082
rect 100680 3998 100892 4026
rect 100576 3392 100628 3398
rect 100576 3334 100628 3340
rect 100574 3224 100630 3233
rect 100574 3159 100630 3168
rect 100588 3126 100616 3159
rect 100576 3120 100628 3126
rect 100576 3062 100628 3068
rect 100680 2774 100708 3998
rect 100760 3392 100812 3398
rect 100760 3334 100812 3340
rect 100772 3097 100800 3334
rect 102428 3194 102456 28494
rect 104164 4480 104216 4486
rect 104164 4422 104216 4428
rect 104176 4282 104204 4422
rect 104164 4276 104216 4282
rect 104164 4218 104216 4224
rect 104452 3194 104480 29582
rect 106016 3670 106044 30194
rect 106004 3664 106056 3670
rect 106004 3606 106056 3612
rect 106096 3664 106148 3670
rect 106096 3606 106148 3612
rect 105820 3528 105872 3534
rect 106108 3482 106136 3606
rect 105820 3470 105872 3476
rect 102416 3188 102468 3194
rect 102416 3130 102468 3136
rect 104440 3188 104492 3194
rect 104440 3130 104492 3136
rect 100758 3088 100814 3097
rect 100758 3023 100814 3032
rect 101220 3052 101272 3058
rect 100772 2990 100800 3023
rect 101220 2994 101272 3000
rect 102140 3052 102192 3058
rect 102140 2994 102192 3000
rect 104256 3052 104308 3058
rect 104256 2994 104308 3000
rect 104900 3052 104952 3058
rect 104900 2994 104952 3000
rect 105268 3052 105320 3058
rect 105268 2994 105320 3000
rect 100760 2984 100812 2990
rect 100760 2926 100812 2932
rect 100588 2746 100708 2774
rect 100300 2508 100352 2514
rect 99392 1630 99420 2502
rect 100300 2450 100352 2456
rect 100392 2508 100444 2514
rect 100392 2450 100444 2456
rect 99472 2372 99524 2378
rect 99472 2314 99524 2320
rect 99484 1698 99512 2314
rect 100312 1902 100340 2450
rect 100300 1896 100352 1902
rect 100300 1838 100352 1844
rect 99472 1692 99524 1698
rect 99472 1634 99524 1640
rect 99380 1624 99432 1630
rect 99380 1566 99432 1572
rect 98460 1420 98512 1426
rect 98460 1362 98512 1368
rect 99196 1420 99248 1426
rect 99196 1362 99248 1368
rect 98092 1148 98144 1154
rect 98092 1090 98144 1096
rect 99208 800 99236 1362
rect 100588 800 100616 2746
rect 100668 2304 100720 2310
rect 100668 2246 100720 2252
rect 100760 2304 100812 2310
rect 100760 2246 100812 2252
rect 100680 1086 100708 2246
rect 100668 1080 100720 1086
rect 100668 1022 100720 1028
rect 96896 740 96948 746
rect 96896 682 96948 688
rect 97722 0 97778 800
rect 99194 0 99250 800
rect 100574 0 100630 800
rect 100772 678 100800 2246
rect 101232 1426 101260 2994
rect 102048 2984 102100 2990
rect 102048 2926 102100 2932
rect 101220 1420 101272 1426
rect 101220 1362 101272 1368
rect 102060 800 102088 2926
rect 102152 2650 102180 2994
rect 102324 2848 102376 2854
rect 102324 2790 102376 2796
rect 102968 2848 103020 2854
rect 102968 2790 103020 2796
rect 102140 2644 102192 2650
rect 102140 2586 102192 2592
rect 102336 2514 102364 2790
rect 102324 2508 102376 2514
rect 102324 2450 102376 2456
rect 102980 2446 103008 2790
rect 104268 2650 104296 2994
rect 104256 2644 104308 2650
rect 104256 2586 104308 2592
rect 103520 2508 103572 2514
rect 103520 2450 103572 2456
rect 102968 2440 103020 2446
rect 102968 2382 103020 2388
rect 103428 2372 103480 2378
rect 103428 2314 103480 2320
rect 103244 2304 103296 2310
rect 103244 2246 103296 2252
rect 103256 882 103284 2246
rect 103244 876 103296 882
rect 103244 818 103296 824
rect 103440 800 103468 2314
rect 103532 1970 103560 2450
rect 103520 1964 103572 1970
rect 103520 1906 103572 1912
rect 104912 800 104940 2994
rect 105176 2848 105228 2854
rect 105176 2790 105228 2796
rect 105188 2514 105216 2790
rect 105176 2508 105228 2514
rect 105176 2450 105228 2456
rect 105280 1494 105308 2994
rect 105832 2650 105860 3470
rect 106016 3454 106136 3482
rect 106280 3528 106332 3534
rect 106280 3470 106332 3476
rect 106016 3398 106044 3454
rect 106004 3392 106056 3398
rect 106004 3334 106056 3340
rect 106096 3392 106148 3398
rect 106096 3334 106148 3340
rect 106108 3194 106136 3334
rect 106096 3188 106148 3194
rect 106096 3130 106148 3136
rect 106188 2984 106240 2990
rect 106188 2926 106240 2932
rect 105820 2644 105872 2650
rect 105820 2586 105872 2592
rect 106200 2582 106228 2926
rect 106188 2576 106240 2582
rect 105450 2544 105506 2553
rect 106188 2518 106240 2524
rect 105450 2479 105506 2488
rect 105464 2446 105492 2479
rect 105452 2440 105504 2446
rect 105728 2440 105780 2446
rect 105452 2382 105504 2388
rect 105726 2408 105728 2417
rect 105780 2408 105782 2417
rect 106200 2378 106228 2518
rect 105726 2343 105782 2352
rect 106188 2372 106240 2378
rect 106188 2314 106240 2320
rect 105268 1488 105320 1494
rect 105268 1430 105320 1436
rect 106292 800 106320 3470
rect 107120 3194 107148 31282
rect 107660 9920 107712 9926
rect 107660 9862 107712 9868
rect 107672 3670 107700 9862
rect 107660 3664 107712 3670
rect 107660 3606 107712 3612
rect 108500 3194 108528 32370
rect 110800 3194 110828 33458
rect 111734 32668 112042 32688
rect 111734 32666 111740 32668
rect 111796 32666 111820 32668
rect 111876 32666 111900 32668
rect 111956 32666 111980 32668
rect 112036 32666 112042 32668
rect 111796 32614 111798 32666
rect 111978 32614 111980 32666
rect 111734 32612 111740 32614
rect 111796 32612 111820 32614
rect 111876 32612 111900 32614
rect 111956 32612 111980 32614
rect 112036 32612 112042 32614
rect 111734 32592 112042 32612
rect 111734 31580 112042 31600
rect 111734 31578 111740 31580
rect 111796 31578 111820 31580
rect 111876 31578 111900 31580
rect 111956 31578 111980 31580
rect 112036 31578 112042 31580
rect 111796 31526 111798 31578
rect 111978 31526 111980 31578
rect 111734 31524 111740 31526
rect 111796 31524 111820 31526
rect 111876 31524 111900 31526
rect 111956 31524 111980 31526
rect 112036 31524 112042 31526
rect 111734 31504 112042 31524
rect 111734 30492 112042 30512
rect 111734 30490 111740 30492
rect 111796 30490 111820 30492
rect 111876 30490 111900 30492
rect 111956 30490 111980 30492
rect 112036 30490 112042 30492
rect 111796 30438 111798 30490
rect 111978 30438 111980 30490
rect 111734 30436 111740 30438
rect 111796 30436 111820 30438
rect 111876 30436 111900 30438
rect 111956 30436 111980 30438
rect 112036 30436 112042 30438
rect 111734 30416 112042 30436
rect 111734 29404 112042 29424
rect 111734 29402 111740 29404
rect 111796 29402 111820 29404
rect 111876 29402 111900 29404
rect 111956 29402 111980 29404
rect 112036 29402 112042 29404
rect 111796 29350 111798 29402
rect 111978 29350 111980 29402
rect 111734 29348 111740 29350
rect 111796 29348 111820 29350
rect 111876 29348 111900 29350
rect 111956 29348 111980 29350
rect 112036 29348 112042 29350
rect 111734 29328 112042 29348
rect 111734 28316 112042 28336
rect 111734 28314 111740 28316
rect 111796 28314 111820 28316
rect 111876 28314 111900 28316
rect 111956 28314 111980 28316
rect 112036 28314 112042 28316
rect 111796 28262 111798 28314
rect 111978 28262 111980 28314
rect 111734 28260 111740 28262
rect 111796 28260 111820 28262
rect 111876 28260 111900 28262
rect 111956 28260 111980 28262
rect 112036 28260 112042 28262
rect 111734 28240 112042 28260
rect 111734 27228 112042 27248
rect 111734 27226 111740 27228
rect 111796 27226 111820 27228
rect 111876 27226 111900 27228
rect 111956 27226 111980 27228
rect 112036 27226 112042 27228
rect 111796 27174 111798 27226
rect 111978 27174 111980 27226
rect 111734 27172 111740 27174
rect 111796 27172 111820 27174
rect 111876 27172 111900 27174
rect 111956 27172 111980 27174
rect 112036 27172 112042 27174
rect 111734 27152 112042 27172
rect 111734 26140 112042 26160
rect 111734 26138 111740 26140
rect 111796 26138 111820 26140
rect 111876 26138 111900 26140
rect 111956 26138 111980 26140
rect 112036 26138 112042 26140
rect 111796 26086 111798 26138
rect 111978 26086 111980 26138
rect 111734 26084 111740 26086
rect 111796 26084 111820 26086
rect 111876 26084 111900 26086
rect 111956 26084 111980 26086
rect 112036 26084 112042 26086
rect 111734 26064 112042 26084
rect 111734 25052 112042 25072
rect 111734 25050 111740 25052
rect 111796 25050 111820 25052
rect 111876 25050 111900 25052
rect 111956 25050 111980 25052
rect 112036 25050 112042 25052
rect 111796 24998 111798 25050
rect 111978 24998 111980 25050
rect 111734 24996 111740 24998
rect 111796 24996 111820 24998
rect 111876 24996 111900 24998
rect 111956 24996 111980 24998
rect 112036 24996 112042 24998
rect 111734 24976 112042 24996
rect 111734 23964 112042 23984
rect 111734 23962 111740 23964
rect 111796 23962 111820 23964
rect 111876 23962 111900 23964
rect 111956 23962 111980 23964
rect 112036 23962 112042 23964
rect 111796 23910 111798 23962
rect 111978 23910 111980 23962
rect 111734 23908 111740 23910
rect 111796 23908 111820 23910
rect 111876 23908 111900 23910
rect 111956 23908 111980 23910
rect 112036 23908 112042 23910
rect 111734 23888 112042 23908
rect 111734 22876 112042 22896
rect 111734 22874 111740 22876
rect 111796 22874 111820 22876
rect 111876 22874 111900 22876
rect 111956 22874 111980 22876
rect 112036 22874 112042 22876
rect 111796 22822 111798 22874
rect 111978 22822 111980 22874
rect 111734 22820 111740 22822
rect 111796 22820 111820 22822
rect 111876 22820 111900 22822
rect 111956 22820 111980 22822
rect 112036 22820 112042 22822
rect 111734 22800 112042 22820
rect 111734 21788 112042 21808
rect 111734 21786 111740 21788
rect 111796 21786 111820 21788
rect 111876 21786 111900 21788
rect 111956 21786 111980 21788
rect 112036 21786 112042 21788
rect 111796 21734 111798 21786
rect 111978 21734 111980 21786
rect 111734 21732 111740 21734
rect 111796 21732 111820 21734
rect 111876 21732 111900 21734
rect 111956 21732 111980 21734
rect 112036 21732 112042 21734
rect 111734 21712 112042 21732
rect 111734 20700 112042 20720
rect 111734 20698 111740 20700
rect 111796 20698 111820 20700
rect 111876 20698 111900 20700
rect 111956 20698 111980 20700
rect 112036 20698 112042 20700
rect 111796 20646 111798 20698
rect 111978 20646 111980 20698
rect 111734 20644 111740 20646
rect 111796 20644 111820 20646
rect 111876 20644 111900 20646
rect 111956 20644 111980 20646
rect 112036 20644 112042 20646
rect 111734 20624 112042 20644
rect 111734 19612 112042 19632
rect 111734 19610 111740 19612
rect 111796 19610 111820 19612
rect 111876 19610 111900 19612
rect 111956 19610 111980 19612
rect 112036 19610 112042 19612
rect 111796 19558 111798 19610
rect 111978 19558 111980 19610
rect 111734 19556 111740 19558
rect 111796 19556 111820 19558
rect 111876 19556 111900 19558
rect 111956 19556 111980 19558
rect 112036 19556 112042 19558
rect 111734 19536 112042 19556
rect 111734 18524 112042 18544
rect 111734 18522 111740 18524
rect 111796 18522 111820 18524
rect 111876 18522 111900 18524
rect 111956 18522 111980 18524
rect 112036 18522 112042 18524
rect 111796 18470 111798 18522
rect 111978 18470 111980 18522
rect 111734 18468 111740 18470
rect 111796 18468 111820 18470
rect 111876 18468 111900 18470
rect 111956 18468 111980 18470
rect 112036 18468 112042 18470
rect 111734 18448 112042 18468
rect 111734 17436 112042 17456
rect 111734 17434 111740 17436
rect 111796 17434 111820 17436
rect 111876 17434 111900 17436
rect 111956 17434 111980 17436
rect 112036 17434 112042 17436
rect 111796 17382 111798 17434
rect 111978 17382 111980 17434
rect 111734 17380 111740 17382
rect 111796 17380 111820 17382
rect 111876 17380 111900 17382
rect 111956 17380 111980 17382
rect 112036 17380 112042 17382
rect 111734 17360 112042 17380
rect 111734 16348 112042 16368
rect 111734 16346 111740 16348
rect 111796 16346 111820 16348
rect 111876 16346 111900 16348
rect 111956 16346 111980 16348
rect 112036 16346 112042 16348
rect 111796 16294 111798 16346
rect 111978 16294 111980 16346
rect 111734 16292 111740 16294
rect 111796 16292 111820 16294
rect 111876 16292 111900 16294
rect 111956 16292 111980 16294
rect 112036 16292 112042 16294
rect 111734 16272 112042 16292
rect 111734 15260 112042 15280
rect 111734 15258 111740 15260
rect 111796 15258 111820 15260
rect 111876 15258 111900 15260
rect 111956 15258 111980 15260
rect 112036 15258 112042 15260
rect 111796 15206 111798 15258
rect 111978 15206 111980 15258
rect 111734 15204 111740 15206
rect 111796 15204 111820 15206
rect 111876 15204 111900 15206
rect 111956 15204 111980 15206
rect 112036 15204 112042 15206
rect 111734 15184 112042 15204
rect 111734 14172 112042 14192
rect 111734 14170 111740 14172
rect 111796 14170 111820 14172
rect 111876 14170 111900 14172
rect 111956 14170 111980 14172
rect 112036 14170 112042 14172
rect 111796 14118 111798 14170
rect 111978 14118 111980 14170
rect 111734 14116 111740 14118
rect 111796 14116 111820 14118
rect 111876 14116 111900 14118
rect 111956 14116 111980 14118
rect 112036 14116 112042 14118
rect 111734 14096 112042 14116
rect 111734 13084 112042 13104
rect 111734 13082 111740 13084
rect 111796 13082 111820 13084
rect 111876 13082 111900 13084
rect 111956 13082 111980 13084
rect 112036 13082 112042 13084
rect 111796 13030 111798 13082
rect 111978 13030 111980 13082
rect 111734 13028 111740 13030
rect 111796 13028 111820 13030
rect 111876 13028 111900 13030
rect 111956 13028 111980 13030
rect 112036 13028 112042 13030
rect 111734 13008 112042 13028
rect 111734 11996 112042 12016
rect 111734 11994 111740 11996
rect 111796 11994 111820 11996
rect 111876 11994 111900 11996
rect 111956 11994 111980 11996
rect 112036 11994 112042 11996
rect 111796 11942 111798 11994
rect 111978 11942 111980 11994
rect 111734 11940 111740 11942
rect 111796 11940 111820 11942
rect 111876 11940 111900 11942
rect 111956 11940 111980 11942
rect 112036 11940 112042 11942
rect 111734 11920 112042 11940
rect 111734 10908 112042 10928
rect 111734 10906 111740 10908
rect 111796 10906 111820 10908
rect 111876 10906 111900 10908
rect 111956 10906 111980 10908
rect 112036 10906 112042 10908
rect 111796 10854 111798 10906
rect 111978 10854 111980 10906
rect 111734 10852 111740 10854
rect 111796 10852 111820 10854
rect 111876 10852 111900 10854
rect 111956 10852 111980 10854
rect 112036 10852 112042 10854
rect 111734 10832 112042 10852
rect 111734 9820 112042 9840
rect 111734 9818 111740 9820
rect 111796 9818 111820 9820
rect 111876 9818 111900 9820
rect 111956 9818 111980 9820
rect 112036 9818 112042 9820
rect 111796 9766 111798 9818
rect 111978 9766 111980 9818
rect 111734 9764 111740 9766
rect 111796 9764 111820 9766
rect 111876 9764 111900 9766
rect 111956 9764 111980 9766
rect 112036 9764 112042 9766
rect 111734 9744 112042 9764
rect 111734 8732 112042 8752
rect 111734 8730 111740 8732
rect 111796 8730 111820 8732
rect 111876 8730 111900 8732
rect 111956 8730 111980 8732
rect 112036 8730 112042 8732
rect 111796 8678 111798 8730
rect 111978 8678 111980 8730
rect 111734 8676 111740 8678
rect 111796 8676 111820 8678
rect 111876 8676 111900 8678
rect 111956 8676 111980 8678
rect 112036 8676 112042 8678
rect 111734 8656 112042 8676
rect 111734 7644 112042 7664
rect 111734 7642 111740 7644
rect 111796 7642 111820 7644
rect 111876 7642 111900 7644
rect 111956 7642 111980 7644
rect 112036 7642 112042 7644
rect 111796 7590 111798 7642
rect 111978 7590 111980 7642
rect 111734 7588 111740 7590
rect 111796 7588 111820 7590
rect 111876 7588 111900 7590
rect 111956 7588 111980 7590
rect 112036 7588 112042 7590
rect 111734 7568 112042 7588
rect 111734 6556 112042 6576
rect 111734 6554 111740 6556
rect 111796 6554 111820 6556
rect 111876 6554 111900 6556
rect 111956 6554 111980 6556
rect 112036 6554 112042 6556
rect 111796 6502 111798 6554
rect 111978 6502 111980 6554
rect 111734 6500 111740 6502
rect 111796 6500 111820 6502
rect 111876 6500 111900 6502
rect 111956 6500 111980 6502
rect 112036 6500 112042 6502
rect 111734 6480 112042 6500
rect 111734 5468 112042 5488
rect 111734 5466 111740 5468
rect 111796 5466 111820 5468
rect 111876 5466 111900 5468
rect 111956 5466 111980 5468
rect 112036 5466 112042 5468
rect 111796 5414 111798 5466
rect 111978 5414 111980 5466
rect 111734 5412 111740 5414
rect 111796 5412 111820 5414
rect 111876 5412 111900 5414
rect 111956 5412 111980 5414
rect 112036 5412 112042 5414
rect 111734 5392 112042 5412
rect 111734 4380 112042 4400
rect 111734 4378 111740 4380
rect 111796 4378 111820 4380
rect 111876 4378 111900 4380
rect 111956 4378 111980 4380
rect 112036 4378 112042 4380
rect 111796 4326 111798 4378
rect 111978 4326 111980 4378
rect 111734 4324 111740 4326
rect 111796 4324 111820 4326
rect 111876 4324 111900 4326
rect 111956 4324 111980 4326
rect 112036 4324 112042 4326
rect 111734 4304 112042 4324
rect 111708 4004 111760 4010
rect 111708 3946 111760 3952
rect 111524 3936 111576 3942
rect 111720 3890 111748 3946
rect 111576 3884 111748 3890
rect 111524 3878 111748 3884
rect 111536 3862 111748 3878
rect 112076 3392 112128 3398
rect 112076 3334 112128 3340
rect 111734 3292 112042 3312
rect 111734 3290 111740 3292
rect 111796 3290 111820 3292
rect 111876 3290 111900 3292
rect 111956 3290 111980 3292
rect 112036 3290 112042 3292
rect 111796 3238 111798 3290
rect 111978 3238 111980 3290
rect 111734 3236 111740 3238
rect 111796 3236 111820 3238
rect 111876 3236 111900 3238
rect 111956 3236 111980 3238
rect 112036 3236 112042 3238
rect 111734 3216 112042 3236
rect 107108 3188 107160 3194
rect 107108 3130 107160 3136
rect 108488 3188 108540 3194
rect 108488 3130 108540 3136
rect 110788 3188 110840 3194
rect 110788 3130 110840 3136
rect 107752 3052 107804 3058
rect 107752 2994 107804 3000
rect 108304 3052 108356 3058
rect 108304 2994 108356 3000
rect 109040 3052 109092 3058
rect 109040 2994 109092 3000
rect 110512 3052 110564 3058
rect 110512 2994 110564 3000
rect 110696 3052 110748 3058
rect 110696 2994 110748 3000
rect 107660 2848 107712 2854
rect 107660 2790 107712 2796
rect 107672 2514 107700 2790
rect 107660 2508 107712 2514
rect 107660 2450 107712 2456
rect 107764 800 107792 2994
rect 108316 2650 108344 2994
rect 108304 2644 108356 2650
rect 108304 2586 108356 2592
rect 109052 2446 109080 2994
rect 109960 2984 110012 2990
rect 109960 2926 110012 2932
rect 109972 2514 110000 2926
rect 110524 2650 110552 2994
rect 110512 2644 110564 2650
rect 110512 2586 110564 2592
rect 110708 2582 110736 2994
rect 110696 2576 110748 2582
rect 110696 2518 110748 2524
rect 112088 2514 112116 3334
rect 112180 3194 112208 33934
rect 114744 4208 114796 4214
rect 114744 4150 114796 4156
rect 113364 4072 113416 4078
rect 113364 4014 113416 4020
rect 113376 3738 113404 4014
rect 114756 3942 114784 4150
rect 114836 4140 114888 4146
rect 114836 4082 114888 4088
rect 114744 3936 114796 3942
rect 114744 3878 114796 3884
rect 113272 3732 113324 3738
rect 113272 3674 113324 3680
rect 113364 3732 113416 3738
rect 113364 3674 113416 3680
rect 112260 3528 112312 3534
rect 112260 3470 112312 3476
rect 112168 3188 112220 3194
rect 112168 3130 112220 3136
rect 109960 2508 110012 2514
rect 109960 2450 110012 2456
rect 110604 2508 110656 2514
rect 110604 2450 110656 2456
rect 112076 2508 112128 2514
rect 112076 2450 112128 2456
rect 109040 2440 109092 2446
rect 109040 2382 109092 2388
rect 109132 2440 109184 2446
rect 109132 2382 109184 2388
rect 108672 2372 108724 2378
rect 108672 2314 108724 2320
rect 108684 1970 108712 2314
rect 108672 1964 108724 1970
rect 108672 1906 108724 1912
rect 109144 800 109172 2382
rect 109776 2304 109828 2310
rect 109776 2246 109828 2252
rect 109788 1358 109816 2246
rect 109776 1352 109828 1358
rect 109776 1294 109828 1300
rect 110616 800 110644 2450
rect 111524 2304 111576 2310
rect 111524 2246 111576 2252
rect 111536 2038 111564 2246
rect 111734 2204 112042 2224
rect 111734 2202 111740 2204
rect 111796 2202 111820 2204
rect 111876 2202 111900 2204
rect 111956 2202 111980 2204
rect 112036 2202 112042 2204
rect 111796 2150 111798 2202
rect 111978 2150 111980 2202
rect 111734 2148 111740 2150
rect 111796 2148 111820 2150
rect 111876 2148 111900 2150
rect 111956 2148 111980 2150
rect 112036 2148 112042 2150
rect 111734 2128 112042 2148
rect 111524 2032 111576 2038
rect 111524 1974 111576 1980
rect 111996 836 112116 864
rect 111996 800 112024 836
rect 100760 672 100812 678
rect 100760 614 100812 620
rect 102046 0 102102 800
rect 103426 0 103482 800
rect 104898 0 104954 800
rect 106278 0 106334 800
rect 107750 0 107806 800
rect 109130 0 109186 800
rect 110602 0 110658 800
rect 111982 0 112038 800
rect 112088 762 112116 836
rect 112272 762 112300 3470
rect 113284 3210 113312 3674
rect 114008 3596 114060 3602
rect 114008 3538 114060 3544
rect 114100 3596 114152 3602
rect 114100 3538 114152 3544
rect 113284 3182 113680 3210
rect 114020 3194 114048 3538
rect 112536 3052 112588 3058
rect 112536 2994 112588 3000
rect 113456 3052 113508 3058
rect 113456 2994 113508 3000
rect 112548 2378 112576 2994
rect 112628 2848 112680 2854
rect 112628 2790 112680 2796
rect 112640 2514 112668 2790
rect 112628 2508 112680 2514
rect 112628 2450 112680 2456
rect 112536 2372 112588 2378
rect 112536 2314 112588 2320
rect 113468 800 113496 2994
rect 113652 2854 113680 3182
rect 114008 3188 114060 3194
rect 114008 3130 114060 3136
rect 113548 2848 113600 2854
rect 113548 2790 113600 2796
rect 113640 2848 113692 2854
rect 113640 2790 113692 2796
rect 113560 2514 113588 2790
rect 114112 2650 114140 3538
rect 114100 2644 114152 2650
rect 114100 2586 114152 2592
rect 113548 2508 113600 2514
rect 113548 2450 113600 2456
rect 113640 2372 113692 2378
rect 113640 2314 113692 2320
rect 113652 2106 113680 2314
rect 113640 2100 113692 2106
rect 113640 2042 113692 2048
rect 114848 800 114876 4082
rect 114940 3670 114968 37198
rect 117148 36922 117176 39471
rect 117226 38584 117282 38593
rect 117226 38519 117282 38528
rect 117240 37466 117268 38519
rect 118054 37632 118110 37641
rect 118054 37567 118110 37576
rect 118068 37466 118096 37567
rect 117228 37460 117280 37466
rect 117228 37402 117280 37408
rect 118056 37460 118108 37466
rect 118056 37402 118108 37408
rect 117596 37256 117648 37262
rect 117596 37198 117648 37204
rect 117136 36916 117188 36922
rect 117136 36858 117188 36864
rect 117412 19168 117464 19174
rect 117412 19110 117464 19116
rect 116860 7200 116912 7206
rect 116860 7142 116912 7148
rect 116308 5568 116360 5574
rect 116308 5510 116360 5516
rect 116216 4616 116268 4622
rect 116216 4558 116268 4564
rect 115296 4480 115348 4486
rect 115296 4422 115348 4428
rect 114928 3664 114980 3670
rect 114928 3606 114980 3612
rect 115204 3596 115256 3602
rect 115204 3538 115256 3544
rect 115216 3482 115244 3538
rect 114940 3466 115244 3482
rect 114928 3460 115244 3466
rect 114980 3454 115244 3460
rect 114928 3402 114980 3408
rect 115308 2990 115336 4422
rect 116124 4276 116176 4282
rect 116124 4218 116176 4224
rect 115848 4140 115900 4146
rect 115848 4082 115900 4088
rect 115388 3936 115440 3942
rect 115388 3878 115440 3884
rect 115296 2984 115348 2990
rect 115296 2926 115348 2932
rect 115400 2514 115428 3878
rect 115480 2984 115532 2990
rect 115480 2926 115532 2932
rect 115492 2514 115520 2926
rect 115860 2582 115888 4082
rect 116136 3534 116164 4218
rect 116124 3528 116176 3534
rect 116124 3470 116176 3476
rect 116228 3194 116256 4558
rect 116320 3534 116348 5510
rect 116584 4140 116636 4146
rect 116584 4082 116636 4088
rect 116676 4140 116728 4146
rect 116676 4082 116728 4088
rect 116400 3596 116452 3602
rect 116400 3538 116452 3544
rect 116308 3528 116360 3534
rect 116308 3470 116360 3476
rect 116216 3188 116268 3194
rect 116216 3130 116268 3136
rect 116308 3052 116360 3058
rect 116308 2994 116360 3000
rect 115848 2576 115900 2582
rect 115848 2518 115900 2524
rect 115388 2508 115440 2514
rect 115388 2450 115440 2456
rect 115480 2508 115532 2514
rect 115480 2450 115532 2456
rect 115296 2304 115348 2310
rect 115296 2246 115348 2252
rect 115308 1562 115336 2246
rect 115296 1556 115348 1562
rect 115296 1498 115348 1504
rect 116320 800 116348 2994
rect 116412 2990 116440 3538
rect 116400 2984 116452 2990
rect 116400 2926 116452 2932
rect 116596 2650 116624 4082
rect 116688 3942 116716 4082
rect 116676 3936 116728 3942
rect 116676 3878 116728 3884
rect 116872 3466 116900 7142
rect 117424 6322 117452 19110
rect 117504 16448 117556 16454
rect 117504 16390 117556 16396
rect 117412 6316 117464 6322
rect 117412 6258 117464 6264
rect 117516 6202 117544 16390
rect 117424 6174 117544 6202
rect 117228 4208 117280 4214
rect 117228 4150 117280 4156
rect 116860 3460 116912 3466
rect 116860 3402 116912 3408
rect 117136 3460 117188 3466
rect 117136 3402 117188 3408
rect 116584 2644 116636 2650
rect 116584 2586 116636 2592
rect 116492 2440 116544 2446
rect 116492 2382 116544 2388
rect 112088 734 112300 762
rect 113454 0 113510 800
rect 114834 0 114890 800
rect 116306 0 116362 800
rect 116504 513 116532 2382
rect 116768 2372 116820 2378
rect 116768 2314 116820 2320
rect 116780 1222 116808 2314
rect 117148 2281 117176 3402
rect 117240 3233 117268 4150
rect 117226 3224 117282 3233
rect 117226 3159 117282 3168
rect 117424 2922 117452 6174
rect 117504 6112 117556 6118
rect 117504 6054 117556 6060
rect 117516 4282 117544 6054
rect 117608 4826 117636 37198
rect 118424 36780 118476 36786
rect 118424 36722 118476 36728
rect 118054 36680 118110 36689
rect 118054 36615 118056 36624
rect 118108 36615 118110 36624
rect 118056 36586 118108 36592
rect 118148 36168 118200 36174
rect 118148 36110 118200 36116
rect 118056 36032 118108 36038
rect 118056 35974 118108 35980
rect 118068 35737 118096 35974
rect 118054 35728 118110 35737
rect 118054 35663 118110 35672
rect 117688 35080 117740 35086
rect 117688 35022 117740 35028
rect 117700 16574 117728 35022
rect 118056 34944 118108 34950
rect 118056 34886 118108 34892
rect 118068 34785 118096 34886
rect 118054 34776 118110 34785
rect 118054 34711 118110 34720
rect 118054 33960 118110 33969
rect 118054 33895 118110 33904
rect 118068 33862 118096 33895
rect 118056 33856 118108 33862
rect 118056 33798 118108 33804
rect 118056 33312 118108 33318
rect 118056 33254 118108 33260
rect 118068 33017 118096 33254
rect 118054 33008 118110 33017
rect 118054 32943 118110 32952
rect 118056 32224 118108 32230
rect 118056 32166 118108 32172
rect 118068 32065 118096 32166
rect 118054 32056 118110 32065
rect 118054 31991 118110 32000
rect 118056 31136 118108 31142
rect 118054 31104 118056 31113
rect 118108 31104 118110 31113
rect 118054 31039 118110 31048
rect 118054 30152 118110 30161
rect 118054 30087 118056 30096
rect 118108 30087 118110 30096
rect 118056 30058 118108 30064
rect 118056 29504 118108 29510
rect 118056 29446 118108 29452
rect 118068 29209 118096 29446
rect 118054 29200 118110 29209
rect 118054 29135 118110 29144
rect 118056 28416 118108 28422
rect 118054 28384 118056 28393
rect 118108 28384 118110 28393
rect 118054 28319 118110 28328
rect 118054 27432 118110 27441
rect 118054 27367 118110 27376
rect 118068 27334 118096 27367
rect 118056 27328 118108 27334
rect 118056 27270 118108 27276
rect 118056 26784 118108 26790
rect 118056 26726 118108 26732
rect 118068 26489 118096 26726
rect 118054 26480 118110 26489
rect 118054 26415 118110 26424
rect 118056 25696 118108 25702
rect 118056 25638 118108 25644
rect 118068 25537 118096 25638
rect 118054 25528 118110 25537
rect 118054 25463 118110 25472
rect 118056 24608 118108 24614
rect 118054 24576 118056 24585
rect 118108 24576 118110 24585
rect 118054 24511 118110 24520
rect 118054 23624 118110 23633
rect 118054 23559 118056 23568
rect 118108 23559 118110 23568
rect 118056 23530 118108 23536
rect 118056 22976 118108 22982
rect 118056 22918 118108 22924
rect 118068 22817 118096 22918
rect 118054 22808 118110 22817
rect 118054 22743 118110 22752
rect 118056 21888 118108 21894
rect 118054 21856 118056 21865
rect 118108 21856 118110 21865
rect 118054 21791 118110 21800
rect 118054 20904 118110 20913
rect 118054 20839 118110 20848
rect 118068 20806 118096 20839
rect 118056 20800 118108 20806
rect 118056 20742 118108 20748
rect 118056 20256 118108 20262
rect 118056 20198 118108 20204
rect 118068 19961 118096 20198
rect 118054 19952 118110 19961
rect 118054 19887 118110 19896
rect 118056 19168 118108 19174
rect 118056 19110 118108 19116
rect 118068 19009 118096 19110
rect 118054 19000 118110 19009
rect 118054 18935 118110 18944
rect 118056 18080 118108 18086
rect 118054 18048 118056 18057
rect 118108 18048 118110 18057
rect 118054 17983 118110 17992
rect 118056 17536 118108 17542
rect 118056 17478 118108 17484
rect 118068 17241 118096 17478
rect 118054 17232 118110 17241
rect 118054 17167 118110 17176
rect 117700 16546 118004 16574
rect 117780 9988 117832 9994
rect 117780 9930 117832 9936
rect 117792 9761 117820 9930
rect 117778 9752 117834 9761
rect 117778 9687 117834 9696
rect 117780 8900 117832 8906
rect 117780 8842 117832 8848
rect 117792 8809 117820 8842
rect 117778 8800 117834 8809
rect 117778 8735 117834 8744
rect 117778 7848 117834 7857
rect 117778 7783 117780 7792
rect 117832 7783 117834 7792
rect 117780 7754 117832 7760
rect 117780 7404 117832 7410
rect 117780 7346 117832 7352
rect 117792 6905 117820 7346
rect 117778 6896 117834 6905
rect 117778 6831 117834 6840
rect 117780 6316 117832 6322
rect 117780 6258 117832 6264
rect 117792 6089 117820 6258
rect 117778 6080 117834 6089
rect 117778 6015 117834 6024
rect 117688 5704 117740 5710
rect 117688 5646 117740 5652
rect 117596 4820 117648 4826
rect 117596 4762 117648 4768
rect 117504 4276 117556 4282
rect 117504 4218 117556 4224
rect 117412 2916 117464 2922
rect 117412 2858 117464 2864
rect 117596 2440 117648 2446
rect 117596 2382 117648 2388
rect 117134 2272 117190 2281
rect 117134 2207 117190 2216
rect 117608 1902 117636 2382
rect 117596 1896 117648 1902
rect 117596 1838 117648 1844
rect 116768 1216 116820 1222
rect 116768 1158 116820 1164
rect 117700 800 117728 5646
rect 117780 5228 117832 5234
rect 117780 5170 117832 5176
rect 117792 5137 117820 5170
rect 117778 5128 117834 5137
rect 117778 5063 117834 5072
rect 117872 5024 117924 5030
rect 117872 4966 117924 4972
rect 117780 4548 117832 4554
rect 117780 4490 117832 4496
rect 117792 4185 117820 4490
rect 117778 4176 117834 4185
rect 117778 4111 117834 4120
rect 117884 4078 117912 4966
rect 117872 4072 117924 4078
rect 117872 4014 117924 4020
rect 117976 3398 118004 16546
rect 118056 16448 118108 16454
rect 118056 16390 118108 16396
rect 118068 16289 118096 16390
rect 118054 16280 118110 16289
rect 118054 16215 118110 16224
rect 118056 15360 118108 15366
rect 118054 15328 118056 15337
rect 118108 15328 118110 15337
rect 118054 15263 118110 15272
rect 118054 14376 118110 14385
rect 118054 14311 118110 14320
rect 118068 14278 118096 14311
rect 118056 14272 118108 14278
rect 118056 14214 118108 14220
rect 118056 13728 118108 13734
rect 118056 13670 118108 13676
rect 118068 13433 118096 13670
rect 118054 13424 118110 13433
rect 118054 13359 118110 13368
rect 118056 12640 118108 12646
rect 118056 12582 118108 12588
rect 118068 12481 118096 12582
rect 118054 12472 118110 12481
rect 118054 12407 118110 12416
rect 118054 11656 118110 11665
rect 118054 11591 118056 11600
rect 118108 11591 118110 11600
rect 118056 11562 118108 11568
rect 118056 11280 118108 11286
rect 118056 11222 118108 11228
rect 118068 10713 118096 11222
rect 118054 10704 118110 10713
rect 118054 10639 118110 10648
rect 118160 4146 118188 36110
rect 118148 4140 118200 4146
rect 118148 4082 118200 4088
rect 118436 3942 118464 36722
rect 118424 3936 118476 3942
rect 118424 3878 118476 3884
rect 117964 3392 118016 3398
rect 117964 3334 118016 3340
rect 117780 3052 117832 3058
rect 117780 2994 117832 3000
rect 117792 1329 117820 2994
rect 119160 2508 119212 2514
rect 119160 2450 119212 2456
rect 117778 1320 117834 1329
rect 117778 1255 117834 1264
rect 119172 800 119200 2450
rect 116490 504 116546 513
rect 116490 439 116546 448
rect 117686 0 117742 800
rect 119158 0 119214 800
<< via2 >>
rect 117134 39480 117190 39536
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 96380 37562 96436 37564
rect 96460 37562 96516 37564
rect 96540 37562 96596 37564
rect 96620 37562 96676 37564
rect 96380 37510 96426 37562
rect 96426 37510 96436 37562
rect 96460 37510 96490 37562
rect 96490 37510 96502 37562
rect 96502 37510 96516 37562
rect 96540 37510 96554 37562
rect 96554 37510 96566 37562
rect 96566 37510 96596 37562
rect 96620 37510 96630 37562
rect 96630 37510 96676 37562
rect 96380 37508 96436 37510
rect 96460 37508 96516 37510
rect 96540 37508 96596 37510
rect 96620 37508 96676 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 81020 37018 81076 37020
rect 81100 37018 81156 37020
rect 81180 37018 81236 37020
rect 81260 37018 81316 37020
rect 81020 36966 81066 37018
rect 81066 36966 81076 37018
rect 81100 36966 81130 37018
rect 81130 36966 81142 37018
rect 81142 36966 81156 37018
rect 81180 36966 81194 37018
rect 81194 36966 81206 37018
rect 81206 36966 81236 37018
rect 81260 36966 81270 37018
rect 81270 36966 81316 37018
rect 81020 36964 81076 36966
rect 81100 36964 81156 36966
rect 81180 36964 81236 36966
rect 81260 36964 81316 36966
rect 111740 37018 111796 37020
rect 111820 37018 111876 37020
rect 111900 37018 111956 37020
rect 111980 37018 112036 37020
rect 111740 36966 111786 37018
rect 111786 36966 111796 37018
rect 111820 36966 111850 37018
rect 111850 36966 111862 37018
rect 111862 36966 111876 37018
rect 111900 36966 111914 37018
rect 111914 36966 111926 37018
rect 111926 36966 111956 37018
rect 111980 36966 111990 37018
rect 111990 36966 112036 37018
rect 111740 36964 111796 36966
rect 111820 36964 111876 36966
rect 111900 36964 111956 36966
rect 111980 36964 112036 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 96380 36474 96436 36476
rect 96460 36474 96516 36476
rect 96540 36474 96596 36476
rect 96620 36474 96676 36476
rect 96380 36422 96426 36474
rect 96426 36422 96436 36474
rect 96460 36422 96490 36474
rect 96490 36422 96502 36474
rect 96502 36422 96516 36474
rect 96540 36422 96554 36474
rect 96554 36422 96566 36474
rect 96566 36422 96596 36474
rect 96620 36422 96630 36474
rect 96630 36422 96676 36474
rect 96380 36420 96436 36422
rect 96460 36420 96516 36422
rect 96540 36420 96596 36422
rect 96620 36420 96676 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 81020 35930 81076 35932
rect 81100 35930 81156 35932
rect 81180 35930 81236 35932
rect 81260 35930 81316 35932
rect 81020 35878 81066 35930
rect 81066 35878 81076 35930
rect 81100 35878 81130 35930
rect 81130 35878 81142 35930
rect 81142 35878 81156 35930
rect 81180 35878 81194 35930
rect 81194 35878 81206 35930
rect 81206 35878 81236 35930
rect 81260 35878 81270 35930
rect 81270 35878 81316 35930
rect 81020 35876 81076 35878
rect 81100 35876 81156 35878
rect 81180 35876 81236 35878
rect 81260 35876 81316 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 96380 35386 96436 35388
rect 96460 35386 96516 35388
rect 96540 35386 96596 35388
rect 96620 35386 96676 35388
rect 96380 35334 96426 35386
rect 96426 35334 96436 35386
rect 96460 35334 96490 35386
rect 96490 35334 96502 35386
rect 96502 35334 96516 35386
rect 96540 35334 96554 35386
rect 96554 35334 96566 35386
rect 96566 35334 96596 35386
rect 96620 35334 96630 35386
rect 96630 35334 96676 35386
rect 96380 35332 96436 35334
rect 96460 35332 96516 35334
rect 96540 35332 96596 35334
rect 96620 35332 96676 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 81020 34842 81076 34844
rect 81100 34842 81156 34844
rect 81180 34842 81236 34844
rect 81260 34842 81316 34844
rect 81020 34790 81066 34842
rect 81066 34790 81076 34842
rect 81100 34790 81130 34842
rect 81130 34790 81142 34842
rect 81142 34790 81156 34842
rect 81180 34790 81194 34842
rect 81194 34790 81206 34842
rect 81206 34790 81236 34842
rect 81260 34790 81270 34842
rect 81270 34790 81316 34842
rect 81020 34788 81076 34790
rect 81100 34788 81156 34790
rect 81180 34788 81236 34790
rect 81260 34788 81316 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 96380 34298 96436 34300
rect 96460 34298 96516 34300
rect 96540 34298 96596 34300
rect 96620 34298 96676 34300
rect 96380 34246 96426 34298
rect 96426 34246 96436 34298
rect 96460 34246 96490 34298
rect 96490 34246 96502 34298
rect 96502 34246 96516 34298
rect 96540 34246 96554 34298
rect 96554 34246 96566 34298
rect 96566 34246 96596 34298
rect 96620 34246 96630 34298
rect 96630 34246 96676 34298
rect 96380 34244 96436 34246
rect 96460 34244 96516 34246
rect 96540 34244 96596 34246
rect 96620 34244 96676 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 81020 33754 81076 33756
rect 81100 33754 81156 33756
rect 81180 33754 81236 33756
rect 81260 33754 81316 33756
rect 81020 33702 81066 33754
rect 81066 33702 81076 33754
rect 81100 33702 81130 33754
rect 81130 33702 81142 33754
rect 81142 33702 81156 33754
rect 81180 33702 81194 33754
rect 81194 33702 81206 33754
rect 81206 33702 81236 33754
rect 81260 33702 81270 33754
rect 81270 33702 81316 33754
rect 81020 33700 81076 33702
rect 81100 33700 81156 33702
rect 81180 33700 81236 33702
rect 81260 33700 81316 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 96380 33210 96436 33212
rect 96460 33210 96516 33212
rect 96540 33210 96596 33212
rect 96620 33210 96676 33212
rect 96380 33158 96426 33210
rect 96426 33158 96436 33210
rect 96460 33158 96490 33210
rect 96490 33158 96502 33210
rect 96502 33158 96516 33210
rect 96540 33158 96554 33210
rect 96554 33158 96566 33210
rect 96566 33158 96596 33210
rect 96620 33158 96630 33210
rect 96630 33158 96676 33210
rect 96380 33156 96436 33158
rect 96460 33156 96516 33158
rect 96540 33156 96596 33158
rect 96620 33156 96676 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 81020 32666 81076 32668
rect 81100 32666 81156 32668
rect 81180 32666 81236 32668
rect 81260 32666 81316 32668
rect 81020 32614 81066 32666
rect 81066 32614 81076 32666
rect 81100 32614 81130 32666
rect 81130 32614 81142 32666
rect 81142 32614 81156 32666
rect 81180 32614 81194 32666
rect 81194 32614 81206 32666
rect 81206 32614 81236 32666
rect 81260 32614 81270 32666
rect 81270 32614 81316 32666
rect 81020 32612 81076 32614
rect 81100 32612 81156 32614
rect 81180 32612 81236 32614
rect 81260 32612 81316 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 96380 32122 96436 32124
rect 96460 32122 96516 32124
rect 96540 32122 96596 32124
rect 96620 32122 96676 32124
rect 96380 32070 96426 32122
rect 96426 32070 96436 32122
rect 96460 32070 96490 32122
rect 96490 32070 96502 32122
rect 96502 32070 96516 32122
rect 96540 32070 96554 32122
rect 96554 32070 96566 32122
rect 96566 32070 96596 32122
rect 96620 32070 96630 32122
rect 96630 32070 96676 32122
rect 96380 32068 96436 32070
rect 96460 32068 96516 32070
rect 96540 32068 96596 32070
rect 96620 32068 96676 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 81020 31578 81076 31580
rect 81100 31578 81156 31580
rect 81180 31578 81236 31580
rect 81260 31578 81316 31580
rect 81020 31526 81066 31578
rect 81066 31526 81076 31578
rect 81100 31526 81130 31578
rect 81130 31526 81142 31578
rect 81142 31526 81156 31578
rect 81180 31526 81194 31578
rect 81194 31526 81206 31578
rect 81206 31526 81236 31578
rect 81260 31526 81270 31578
rect 81270 31526 81316 31578
rect 81020 31524 81076 31526
rect 81100 31524 81156 31526
rect 81180 31524 81236 31526
rect 81260 31524 81316 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 96380 31034 96436 31036
rect 96460 31034 96516 31036
rect 96540 31034 96596 31036
rect 96620 31034 96676 31036
rect 96380 30982 96426 31034
rect 96426 30982 96436 31034
rect 96460 30982 96490 31034
rect 96490 30982 96502 31034
rect 96502 30982 96516 31034
rect 96540 30982 96554 31034
rect 96554 30982 96566 31034
rect 96566 30982 96596 31034
rect 96620 30982 96630 31034
rect 96630 30982 96676 31034
rect 96380 30980 96436 30982
rect 96460 30980 96516 30982
rect 96540 30980 96596 30982
rect 96620 30980 96676 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 81020 30490 81076 30492
rect 81100 30490 81156 30492
rect 81180 30490 81236 30492
rect 81260 30490 81316 30492
rect 81020 30438 81066 30490
rect 81066 30438 81076 30490
rect 81100 30438 81130 30490
rect 81130 30438 81142 30490
rect 81142 30438 81156 30490
rect 81180 30438 81194 30490
rect 81194 30438 81206 30490
rect 81206 30438 81236 30490
rect 81260 30438 81270 30490
rect 81270 30438 81316 30490
rect 81020 30436 81076 30438
rect 81100 30436 81156 30438
rect 81180 30436 81236 30438
rect 81260 30436 81316 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 96380 29946 96436 29948
rect 96460 29946 96516 29948
rect 96540 29946 96596 29948
rect 96620 29946 96676 29948
rect 96380 29894 96426 29946
rect 96426 29894 96436 29946
rect 96460 29894 96490 29946
rect 96490 29894 96502 29946
rect 96502 29894 96516 29946
rect 96540 29894 96554 29946
rect 96554 29894 96566 29946
rect 96566 29894 96596 29946
rect 96620 29894 96630 29946
rect 96630 29894 96676 29946
rect 96380 29892 96436 29894
rect 96460 29892 96516 29894
rect 96540 29892 96596 29894
rect 96620 29892 96676 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 81020 29402 81076 29404
rect 81100 29402 81156 29404
rect 81180 29402 81236 29404
rect 81260 29402 81316 29404
rect 81020 29350 81066 29402
rect 81066 29350 81076 29402
rect 81100 29350 81130 29402
rect 81130 29350 81142 29402
rect 81142 29350 81156 29402
rect 81180 29350 81194 29402
rect 81194 29350 81206 29402
rect 81206 29350 81236 29402
rect 81260 29350 81270 29402
rect 81270 29350 81316 29402
rect 81020 29348 81076 29350
rect 81100 29348 81156 29350
rect 81180 29348 81236 29350
rect 81260 29348 81316 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 96380 28858 96436 28860
rect 96460 28858 96516 28860
rect 96540 28858 96596 28860
rect 96620 28858 96676 28860
rect 96380 28806 96426 28858
rect 96426 28806 96436 28858
rect 96460 28806 96490 28858
rect 96490 28806 96502 28858
rect 96502 28806 96516 28858
rect 96540 28806 96554 28858
rect 96554 28806 96566 28858
rect 96566 28806 96596 28858
rect 96620 28806 96630 28858
rect 96630 28806 96676 28858
rect 96380 28804 96436 28806
rect 96460 28804 96516 28806
rect 96540 28804 96596 28806
rect 96620 28804 96676 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 81020 28314 81076 28316
rect 81100 28314 81156 28316
rect 81180 28314 81236 28316
rect 81260 28314 81316 28316
rect 81020 28262 81066 28314
rect 81066 28262 81076 28314
rect 81100 28262 81130 28314
rect 81130 28262 81142 28314
rect 81142 28262 81156 28314
rect 81180 28262 81194 28314
rect 81194 28262 81206 28314
rect 81206 28262 81236 28314
rect 81260 28262 81270 28314
rect 81270 28262 81316 28314
rect 81020 28260 81076 28262
rect 81100 28260 81156 28262
rect 81180 28260 81236 28262
rect 81260 28260 81316 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 96380 27770 96436 27772
rect 96460 27770 96516 27772
rect 96540 27770 96596 27772
rect 96620 27770 96676 27772
rect 96380 27718 96426 27770
rect 96426 27718 96436 27770
rect 96460 27718 96490 27770
rect 96490 27718 96502 27770
rect 96502 27718 96516 27770
rect 96540 27718 96554 27770
rect 96554 27718 96566 27770
rect 96566 27718 96596 27770
rect 96620 27718 96630 27770
rect 96630 27718 96676 27770
rect 96380 27716 96436 27718
rect 96460 27716 96516 27718
rect 96540 27716 96596 27718
rect 96620 27716 96676 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 81020 27226 81076 27228
rect 81100 27226 81156 27228
rect 81180 27226 81236 27228
rect 81260 27226 81316 27228
rect 81020 27174 81066 27226
rect 81066 27174 81076 27226
rect 81100 27174 81130 27226
rect 81130 27174 81142 27226
rect 81142 27174 81156 27226
rect 81180 27174 81194 27226
rect 81194 27174 81206 27226
rect 81206 27174 81236 27226
rect 81260 27174 81270 27226
rect 81270 27174 81316 27226
rect 81020 27172 81076 27174
rect 81100 27172 81156 27174
rect 81180 27172 81236 27174
rect 81260 27172 81316 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 96380 26682 96436 26684
rect 96460 26682 96516 26684
rect 96540 26682 96596 26684
rect 96620 26682 96676 26684
rect 96380 26630 96426 26682
rect 96426 26630 96436 26682
rect 96460 26630 96490 26682
rect 96490 26630 96502 26682
rect 96502 26630 96516 26682
rect 96540 26630 96554 26682
rect 96554 26630 96566 26682
rect 96566 26630 96596 26682
rect 96620 26630 96630 26682
rect 96630 26630 96676 26682
rect 96380 26628 96436 26630
rect 96460 26628 96516 26630
rect 96540 26628 96596 26630
rect 96620 26628 96676 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 81020 26138 81076 26140
rect 81100 26138 81156 26140
rect 81180 26138 81236 26140
rect 81260 26138 81316 26140
rect 81020 26086 81066 26138
rect 81066 26086 81076 26138
rect 81100 26086 81130 26138
rect 81130 26086 81142 26138
rect 81142 26086 81156 26138
rect 81180 26086 81194 26138
rect 81194 26086 81206 26138
rect 81206 26086 81236 26138
rect 81260 26086 81270 26138
rect 81270 26086 81316 26138
rect 81020 26084 81076 26086
rect 81100 26084 81156 26086
rect 81180 26084 81236 26086
rect 81260 26084 81316 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 96380 25594 96436 25596
rect 96460 25594 96516 25596
rect 96540 25594 96596 25596
rect 96620 25594 96676 25596
rect 96380 25542 96426 25594
rect 96426 25542 96436 25594
rect 96460 25542 96490 25594
rect 96490 25542 96502 25594
rect 96502 25542 96516 25594
rect 96540 25542 96554 25594
rect 96554 25542 96566 25594
rect 96566 25542 96596 25594
rect 96620 25542 96630 25594
rect 96630 25542 96676 25594
rect 96380 25540 96436 25542
rect 96460 25540 96516 25542
rect 96540 25540 96596 25542
rect 96620 25540 96676 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 81020 25050 81076 25052
rect 81100 25050 81156 25052
rect 81180 25050 81236 25052
rect 81260 25050 81316 25052
rect 81020 24998 81066 25050
rect 81066 24998 81076 25050
rect 81100 24998 81130 25050
rect 81130 24998 81142 25050
rect 81142 24998 81156 25050
rect 81180 24998 81194 25050
rect 81194 24998 81206 25050
rect 81206 24998 81236 25050
rect 81260 24998 81270 25050
rect 81270 24998 81316 25050
rect 81020 24996 81076 24998
rect 81100 24996 81156 24998
rect 81180 24996 81236 24998
rect 81260 24996 81316 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 96380 24506 96436 24508
rect 96460 24506 96516 24508
rect 96540 24506 96596 24508
rect 96620 24506 96676 24508
rect 96380 24454 96426 24506
rect 96426 24454 96436 24506
rect 96460 24454 96490 24506
rect 96490 24454 96502 24506
rect 96502 24454 96516 24506
rect 96540 24454 96554 24506
rect 96554 24454 96566 24506
rect 96566 24454 96596 24506
rect 96620 24454 96630 24506
rect 96630 24454 96676 24506
rect 96380 24452 96436 24454
rect 96460 24452 96516 24454
rect 96540 24452 96596 24454
rect 96620 24452 96676 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 81020 23962 81076 23964
rect 81100 23962 81156 23964
rect 81180 23962 81236 23964
rect 81260 23962 81316 23964
rect 81020 23910 81066 23962
rect 81066 23910 81076 23962
rect 81100 23910 81130 23962
rect 81130 23910 81142 23962
rect 81142 23910 81156 23962
rect 81180 23910 81194 23962
rect 81194 23910 81206 23962
rect 81206 23910 81236 23962
rect 81260 23910 81270 23962
rect 81270 23910 81316 23962
rect 81020 23908 81076 23910
rect 81100 23908 81156 23910
rect 81180 23908 81236 23910
rect 81260 23908 81316 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 81020 22874 81076 22876
rect 81100 22874 81156 22876
rect 81180 22874 81236 22876
rect 81260 22874 81316 22876
rect 81020 22822 81066 22874
rect 81066 22822 81076 22874
rect 81100 22822 81130 22874
rect 81130 22822 81142 22874
rect 81142 22822 81156 22874
rect 81180 22822 81194 22874
rect 81194 22822 81206 22874
rect 81206 22822 81236 22874
rect 81260 22822 81270 22874
rect 81270 22822 81316 22874
rect 81020 22820 81076 22822
rect 81100 22820 81156 22822
rect 81180 22820 81236 22822
rect 81260 22820 81316 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 81020 21786 81076 21788
rect 81100 21786 81156 21788
rect 81180 21786 81236 21788
rect 81260 21786 81316 21788
rect 81020 21734 81066 21786
rect 81066 21734 81076 21786
rect 81100 21734 81130 21786
rect 81130 21734 81142 21786
rect 81142 21734 81156 21786
rect 81180 21734 81194 21786
rect 81194 21734 81206 21786
rect 81206 21734 81236 21786
rect 81260 21734 81270 21786
rect 81270 21734 81316 21786
rect 81020 21732 81076 21734
rect 81100 21732 81156 21734
rect 81180 21732 81236 21734
rect 81260 21732 81316 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 81020 20698 81076 20700
rect 81100 20698 81156 20700
rect 81180 20698 81236 20700
rect 81260 20698 81316 20700
rect 81020 20646 81066 20698
rect 81066 20646 81076 20698
rect 81100 20646 81130 20698
rect 81130 20646 81142 20698
rect 81142 20646 81156 20698
rect 81180 20646 81194 20698
rect 81194 20646 81206 20698
rect 81206 20646 81236 20698
rect 81260 20646 81270 20698
rect 81270 20646 81316 20698
rect 81020 20644 81076 20646
rect 81100 20644 81156 20646
rect 81180 20644 81236 20646
rect 81260 20644 81316 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 81020 19610 81076 19612
rect 81100 19610 81156 19612
rect 81180 19610 81236 19612
rect 81260 19610 81316 19612
rect 81020 19558 81066 19610
rect 81066 19558 81076 19610
rect 81100 19558 81130 19610
rect 81130 19558 81142 19610
rect 81142 19558 81156 19610
rect 81180 19558 81194 19610
rect 81194 19558 81206 19610
rect 81206 19558 81236 19610
rect 81260 19558 81270 19610
rect 81270 19558 81316 19610
rect 81020 19556 81076 19558
rect 81100 19556 81156 19558
rect 81180 19556 81236 19558
rect 81260 19556 81316 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 81020 18522 81076 18524
rect 81100 18522 81156 18524
rect 81180 18522 81236 18524
rect 81260 18522 81316 18524
rect 81020 18470 81066 18522
rect 81066 18470 81076 18522
rect 81100 18470 81130 18522
rect 81130 18470 81142 18522
rect 81142 18470 81156 18522
rect 81180 18470 81194 18522
rect 81194 18470 81206 18522
rect 81206 18470 81236 18522
rect 81260 18470 81270 18522
rect 81270 18470 81316 18522
rect 81020 18468 81076 18470
rect 81100 18468 81156 18470
rect 81180 18468 81236 18470
rect 81260 18468 81316 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 81020 17434 81076 17436
rect 81100 17434 81156 17436
rect 81180 17434 81236 17436
rect 81260 17434 81316 17436
rect 81020 17382 81066 17434
rect 81066 17382 81076 17434
rect 81100 17382 81130 17434
rect 81130 17382 81142 17434
rect 81142 17382 81156 17434
rect 81180 17382 81194 17434
rect 81194 17382 81206 17434
rect 81206 17382 81236 17434
rect 81260 17382 81270 17434
rect 81270 17382 81316 17434
rect 81020 17380 81076 17382
rect 81100 17380 81156 17382
rect 81180 17380 81236 17382
rect 81260 17380 81316 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 81020 16346 81076 16348
rect 81100 16346 81156 16348
rect 81180 16346 81236 16348
rect 81260 16346 81316 16348
rect 81020 16294 81066 16346
rect 81066 16294 81076 16346
rect 81100 16294 81130 16346
rect 81130 16294 81142 16346
rect 81142 16294 81156 16346
rect 81180 16294 81194 16346
rect 81194 16294 81206 16346
rect 81206 16294 81236 16346
rect 81260 16294 81270 16346
rect 81270 16294 81316 16346
rect 81020 16292 81076 16294
rect 81100 16292 81156 16294
rect 81180 16292 81236 16294
rect 81260 16292 81316 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 81020 15258 81076 15260
rect 81100 15258 81156 15260
rect 81180 15258 81236 15260
rect 81260 15258 81316 15260
rect 81020 15206 81066 15258
rect 81066 15206 81076 15258
rect 81100 15206 81130 15258
rect 81130 15206 81142 15258
rect 81142 15206 81156 15258
rect 81180 15206 81194 15258
rect 81194 15206 81206 15258
rect 81206 15206 81236 15258
rect 81260 15206 81270 15258
rect 81270 15206 81316 15258
rect 81020 15204 81076 15206
rect 81100 15204 81156 15206
rect 81180 15204 81236 15206
rect 81260 15204 81316 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 81020 14170 81076 14172
rect 81100 14170 81156 14172
rect 81180 14170 81236 14172
rect 81260 14170 81316 14172
rect 81020 14118 81066 14170
rect 81066 14118 81076 14170
rect 81100 14118 81130 14170
rect 81130 14118 81142 14170
rect 81142 14118 81156 14170
rect 81180 14118 81194 14170
rect 81194 14118 81206 14170
rect 81206 14118 81236 14170
rect 81260 14118 81270 14170
rect 81270 14118 81316 14170
rect 81020 14116 81076 14118
rect 81100 14116 81156 14118
rect 81180 14116 81236 14118
rect 81260 14116 81316 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35898 2508 35954 2544
rect 35898 2488 35900 2508
rect 35900 2488 35952 2508
rect 35952 2488 35954 2508
rect 35714 2388 35716 2408
rect 35716 2388 35768 2408
rect 35768 2388 35770 2408
rect 35714 2352 35770 2388
rect 33414 1808 33470 1864
rect 35990 2352 36046 2408
rect 35806 1828 35862 1864
rect 35806 1808 35808 1828
rect 35808 1808 35860 1828
rect 35860 1808 35862 1828
rect 37278 2216 37334 2272
rect 40498 1672 40554 1728
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 45466 2508 45522 2544
rect 45466 2488 45468 2508
rect 45468 2488 45520 2508
rect 45520 2488 45522 2508
rect 45374 2352 45430 2408
rect 45742 2352 45798 2408
rect 45374 2252 45376 2272
rect 45376 2252 45428 2272
rect 45428 2252 45430 2272
rect 45374 2216 45430 2252
rect 45650 1672 45706 1728
rect 49054 2372 49110 2408
rect 49054 2352 49056 2372
rect 49056 2352 49108 2372
rect 49108 2352 49110 2372
rect 53378 2372 53434 2408
rect 53378 2352 53380 2372
rect 53380 2352 53432 2372
rect 53432 2352 53434 2372
rect 47674 1536 47730 1592
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 51078 1944 51134 2000
rect 51078 1808 51134 1864
rect 51170 1672 51226 1728
rect 51262 1556 51318 1592
rect 51262 1536 51264 1556
rect 51264 1536 51316 1556
rect 51316 1536 51318 1556
rect 55770 2508 55826 2544
rect 55770 2488 55772 2508
rect 55772 2488 55824 2508
rect 55824 2488 55826 2508
rect 56690 2624 56746 2680
rect 58438 2488 58494 2544
rect 55678 2252 55680 2272
rect 55680 2252 55732 2272
rect 55732 2252 55734 2272
rect 55678 2216 55734 2252
rect 59818 2760 59874 2816
rect 59634 2352 59690 2408
rect 59726 2252 59728 2272
rect 59728 2252 59780 2272
rect 59780 2252 59782 2272
rect 59726 2216 59782 2252
rect 60278 2508 60334 2544
rect 60278 2488 60280 2508
rect 60280 2488 60332 2508
rect 60332 2488 60334 2508
rect 60186 2216 60242 2272
rect 59910 1944 59966 2000
rect 60370 1944 60426 2000
rect 60186 1808 60242 1864
rect 60738 2216 60794 2272
rect 60554 1672 60610 1728
rect 60738 1420 60794 1456
rect 60738 1400 60740 1420
rect 60740 1400 60792 1420
rect 60792 1400 60794 1420
rect 60462 1264 60518 1320
rect 61290 2624 61346 2680
rect 61198 1264 61254 1320
rect 63406 1808 63462 1864
rect 64142 2488 64198 2544
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 65246 2896 65302 2952
rect 65154 2760 65210 2816
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 66902 2352 66958 2408
rect 67454 2252 67456 2272
rect 67456 2252 67508 2272
rect 67508 2252 67510 2272
rect 67454 2216 67510 2252
rect 69662 2080 69718 2136
rect 70306 1944 70362 2000
rect 70214 1692 70270 1728
rect 70214 1672 70216 1692
rect 70216 1672 70268 1692
rect 70268 1672 70270 1692
rect 69754 1400 69810 1456
rect 74814 2352 74870 2408
rect 74446 2252 74448 2272
rect 74448 2252 74500 2272
rect 74500 2252 74502 2272
rect 74446 2216 74502 2252
rect 73986 1692 74042 1728
rect 73986 1672 73988 1692
rect 73988 1672 74040 1692
rect 74040 1672 74042 1692
rect 76010 1400 76066 1456
rect 81020 13082 81076 13084
rect 81100 13082 81156 13084
rect 81180 13082 81236 13084
rect 81260 13082 81316 13084
rect 81020 13030 81066 13082
rect 81066 13030 81076 13082
rect 81100 13030 81130 13082
rect 81130 13030 81142 13082
rect 81142 13030 81156 13082
rect 81180 13030 81194 13082
rect 81194 13030 81206 13082
rect 81206 13030 81236 13082
rect 81260 13030 81270 13082
rect 81270 13030 81316 13082
rect 81020 13028 81076 13030
rect 81100 13028 81156 13030
rect 81180 13028 81236 13030
rect 81260 13028 81316 13030
rect 81020 11994 81076 11996
rect 81100 11994 81156 11996
rect 81180 11994 81236 11996
rect 81260 11994 81316 11996
rect 81020 11942 81066 11994
rect 81066 11942 81076 11994
rect 81100 11942 81130 11994
rect 81130 11942 81142 11994
rect 81142 11942 81156 11994
rect 81180 11942 81194 11994
rect 81194 11942 81206 11994
rect 81206 11942 81236 11994
rect 81260 11942 81270 11994
rect 81270 11942 81316 11994
rect 81020 11940 81076 11942
rect 81100 11940 81156 11942
rect 81180 11940 81236 11942
rect 81260 11940 81316 11942
rect 81020 10906 81076 10908
rect 81100 10906 81156 10908
rect 81180 10906 81236 10908
rect 81260 10906 81316 10908
rect 81020 10854 81066 10906
rect 81066 10854 81076 10906
rect 81100 10854 81130 10906
rect 81130 10854 81142 10906
rect 81142 10854 81156 10906
rect 81180 10854 81194 10906
rect 81194 10854 81206 10906
rect 81206 10854 81236 10906
rect 81260 10854 81270 10906
rect 81270 10854 81316 10906
rect 81020 10852 81076 10854
rect 81100 10852 81156 10854
rect 81180 10852 81236 10854
rect 81260 10852 81316 10854
rect 81020 9818 81076 9820
rect 81100 9818 81156 9820
rect 81180 9818 81236 9820
rect 81260 9818 81316 9820
rect 81020 9766 81066 9818
rect 81066 9766 81076 9818
rect 81100 9766 81130 9818
rect 81130 9766 81142 9818
rect 81142 9766 81156 9818
rect 81180 9766 81194 9818
rect 81194 9766 81206 9818
rect 81206 9766 81236 9818
rect 81260 9766 81270 9818
rect 81270 9766 81316 9818
rect 81020 9764 81076 9766
rect 81100 9764 81156 9766
rect 81180 9764 81236 9766
rect 81260 9764 81316 9766
rect 81020 8730 81076 8732
rect 81100 8730 81156 8732
rect 81180 8730 81236 8732
rect 81260 8730 81316 8732
rect 81020 8678 81066 8730
rect 81066 8678 81076 8730
rect 81100 8678 81130 8730
rect 81130 8678 81142 8730
rect 81142 8678 81156 8730
rect 81180 8678 81194 8730
rect 81194 8678 81206 8730
rect 81206 8678 81236 8730
rect 81260 8678 81270 8730
rect 81270 8678 81316 8730
rect 81020 8676 81076 8678
rect 81100 8676 81156 8678
rect 81180 8676 81236 8678
rect 81260 8676 81316 8678
rect 81020 7642 81076 7644
rect 81100 7642 81156 7644
rect 81180 7642 81236 7644
rect 81260 7642 81316 7644
rect 81020 7590 81066 7642
rect 81066 7590 81076 7642
rect 81100 7590 81130 7642
rect 81130 7590 81142 7642
rect 81142 7590 81156 7642
rect 81180 7590 81194 7642
rect 81194 7590 81206 7642
rect 81206 7590 81236 7642
rect 81260 7590 81270 7642
rect 81270 7590 81316 7642
rect 81020 7588 81076 7590
rect 81100 7588 81156 7590
rect 81180 7588 81236 7590
rect 81260 7588 81316 7590
rect 81020 6554 81076 6556
rect 81100 6554 81156 6556
rect 81180 6554 81236 6556
rect 81260 6554 81316 6556
rect 81020 6502 81066 6554
rect 81066 6502 81076 6554
rect 81100 6502 81130 6554
rect 81130 6502 81142 6554
rect 81142 6502 81156 6554
rect 81180 6502 81194 6554
rect 81194 6502 81206 6554
rect 81206 6502 81236 6554
rect 81260 6502 81270 6554
rect 81270 6502 81316 6554
rect 81020 6500 81076 6502
rect 81100 6500 81156 6502
rect 81180 6500 81236 6502
rect 81260 6500 81316 6502
rect 81020 5466 81076 5468
rect 81100 5466 81156 5468
rect 81180 5466 81236 5468
rect 81260 5466 81316 5468
rect 81020 5414 81066 5466
rect 81066 5414 81076 5466
rect 81100 5414 81130 5466
rect 81130 5414 81142 5466
rect 81142 5414 81156 5466
rect 81180 5414 81194 5466
rect 81194 5414 81206 5466
rect 81206 5414 81236 5466
rect 81260 5414 81270 5466
rect 81270 5414 81316 5466
rect 81020 5412 81076 5414
rect 81100 5412 81156 5414
rect 81180 5412 81236 5414
rect 81260 5412 81316 5414
rect 81020 4378 81076 4380
rect 81100 4378 81156 4380
rect 81180 4378 81236 4380
rect 81260 4378 81316 4380
rect 81020 4326 81066 4378
rect 81066 4326 81076 4378
rect 81100 4326 81130 4378
rect 81130 4326 81142 4378
rect 81142 4326 81156 4378
rect 81180 4326 81194 4378
rect 81194 4326 81206 4378
rect 81206 4326 81236 4378
rect 81260 4326 81270 4378
rect 81270 4326 81316 4378
rect 81020 4324 81076 4326
rect 81100 4324 81156 4326
rect 81180 4324 81236 4326
rect 81260 4324 81316 4326
rect 81020 3290 81076 3292
rect 81100 3290 81156 3292
rect 81180 3290 81236 3292
rect 81260 3290 81316 3292
rect 81020 3238 81066 3290
rect 81066 3238 81076 3290
rect 81100 3238 81130 3290
rect 81130 3238 81142 3290
rect 81142 3238 81156 3290
rect 81180 3238 81194 3290
rect 81194 3238 81206 3290
rect 81206 3238 81236 3290
rect 81260 3238 81270 3290
rect 81270 3238 81316 3290
rect 81020 3236 81076 3238
rect 81100 3236 81156 3238
rect 81180 3236 81236 3238
rect 81260 3236 81316 3238
rect 77666 1420 77722 1456
rect 77666 1400 77668 1420
rect 77668 1400 77720 1420
rect 77720 1400 77722 1420
rect 79506 2216 79562 2272
rect 81438 2388 81440 2408
rect 81440 2388 81492 2408
rect 81492 2388 81494 2408
rect 81438 2352 81494 2388
rect 81020 2202 81076 2204
rect 81100 2202 81156 2204
rect 81180 2202 81236 2204
rect 81260 2202 81316 2204
rect 81020 2150 81066 2202
rect 81066 2150 81076 2202
rect 81100 2150 81130 2202
rect 81130 2150 81142 2202
rect 81142 2150 81156 2202
rect 81180 2150 81194 2202
rect 81194 2150 81206 2202
rect 81206 2150 81236 2202
rect 81260 2150 81270 2202
rect 81270 2150 81316 2202
rect 81020 2148 81076 2150
rect 81100 2148 81156 2150
rect 81180 2148 81236 2150
rect 81260 2148 81316 2150
rect 96380 23418 96436 23420
rect 96460 23418 96516 23420
rect 96540 23418 96596 23420
rect 96620 23418 96676 23420
rect 96380 23366 96426 23418
rect 96426 23366 96436 23418
rect 96460 23366 96490 23418
rect 96490 23366 96502 23418
rect 96502 23366 96516 23418
rect 96540 23366 96554 23418
rect 96554 23366 96566 23418
rect 96566 23366 96596 23418
rect 96620 23366 96630 23418
rect 96630 23366 96676 23418
rect 96380 23364 96436 23366
rect 96460 23364 96516 23366
rect 96540 23364 96596 23366
rect 96620 23364 96676 23366
rect 96380 22330 96436 22332
rect 96460 22330 96516 22332
rect 96540 22330 96596 22332
rect 96620 22330 96676 22332
rect 96380 22278 96426 22330
rect 96426 22278 96436 22330
rect 96460 22278 96490 22330
rect 96490 22278 96502 22330
rect 96502 22278 96516 22330
rect 96540 22278 96554 22330
rect 96554 22278 96566 22330
rect 96566 22278 96596 22330
rect 96620 22278 96630 22330
rect 96630 22278 96676 22330
rect 96380 22276 96436 22278
rect 96460 22276 96516 22278
rect 96540 22276 96596 22278
rect 96620 22276 96676 22278
rect 96380 21242 96436 21244
rect 96460 21242 96516 21244
rect 96540 21242 96596 21244
rect 96620 21242 96676 21244
rect 96380 21190 96426 21242
rect 96426 21190 96436 21242
rect 96460 21190 96490 21242
rect 96490 21190 96502 21242
rect 96502 21190 96516 21242
rect 96540 21190 96554 21242
rect 96554 21190 96566 21242
rect 96566 21190 96596 21242
rect 96620 21190 96630 21242
rect 96630 21190 96676 21242
rect 96380 21188 96436 21190
rect 96460 21188 96516 21190
rect 96540 21188 96596 21190
rect 96620 21188 96676 21190
rect 96380 20154 96436 20156
rect 96460 20154 96516 20156
rect 96540 20154 96596 20156
rect 96620 20154 96676 20156
rect 96380 20102 96426 20154
rect 96426 20102 96436 20154
rect 96460 20102 96490 20154
rect 96490 20102 96502 20154
rect 96502 20102 96516 20154
rect 96540 20102 96554 20154
rect 96554 20102 96566 20154
rect 96566 20102 96596 20154
rect 96620 20102 96630 20154
rect 96630 20102 96676 20154
rect 96380 20100 96436 20102
rect 96460 20100 96516 20102
rect 96540 20100 96596 20102
rect 96620 20100 96676 20102
rect 96380 19066 96436 19068
rect 96460 19066 96516 19068
rect 96540 19066 96596 19068
rect 96620 19066 96676 19068
rect 96380 19014 96426 19066
rect 96426 19014 96436 19066
rect 96460 19014 96490 19066
rect 96490 19014 96502 19066
rect 96502 19014 96516 19066
rect 96540 19014 96554 19066
rect 96554 19014 96566 19066
rect 96566 19014 96596 19066
rect 96620 19014 96630 19066
rect 96630 19014 96676 19066
rect 96380 19012 96436 19014
rect 96460 19012 96516 19014
rect 96540 19012 96596 19014
rect 96620 19012 96676 19014
rect 96380 17978 96436 17980
rect 96460 17978 96516 17980
rect 96540 17978 96596 17980
rect 96620 17978 96676 17980
rect 96380 17926 96426 17978
rect 96426 17926 96436 17978
rect 96460 17926 96490 17978
rect 96490 17926 96502 17978
rect 96502 17926 96516 17978
rect 96540 17926 96554 17978
rect 96554 17926 96566 17978
rect 96566 17926 96596 17978
rect 96620 17926 96630 17978
rect 96630 17926 96676 17978
rect 96380 17924 96436 17926
rect 96460 17924 96516 17926
rect 96540 17924 96596 17926
rect 96620 17924 96676 17926
rect 96380 16890 96436 16892
rect 96460 16890 96516 16892
rect 96540 16890 96596 16892
rect 96620 16890 96676 16892
rect 96380 16838 96426 16890
rect 96426 16838 96436 16890
rect 96460 16838 96490 16890
rect 96490 16838 96502 16890
rect 96502 16838 96516 16890
rect 96540 16838 96554 16890
rect 96554 16838 96566 16890
rect 96566 16838 96596 16890
rect 96620 16838 96630 16890
rect 96630 16838 96676 16890
rect 96380 16836 96436 16838
rect 96460 16836 96516 16838
rect 96540 16836 96596 16838
rect 96620 16836 96676 16838
rect 96380 15802 96436 15804
rect 96460 15802 96516 15804
rect 96540 15802 96596 15804
rect 96620 15802 96676 15804
rect 96380 15750 96426 15802
rect 96426 15750 96436 15802
rect 96460 15750 96490 15802
rect 96490 15750 96502 15802
rect 96502 15750 96516 15802
rect 96540 15750 96554 15802
rect 96554 15750 96566 15802
rect 96566 15750 96596 15802
rect 96620 15750 96630 15802
rect 96630 15750 96676 15802
rect 96380 15748 96436 15750
rect 96460 15748 96516 15750
rect 96540 15748 96596 15750
rect 96620 15748 96676 15750
rect 96380 14714 96436 14716
rect 96460 14714 96516 14716
rect 96540 14714 96596 14716
rect 96620 14714 96676 14716
rect 96380 14662 96426 14714
rect 96426 14662 96436 14714
rect 96460 14662 96490 14714
rect 96490 14662 96502 14714
rect 96502 14662 96516 14714
rect 96540 14662 96554 14714
rect 96554 14662 96566 14714
rect 96566 14662 96596 14714
rect 96620 14662 96630 14714
rect 96630 14662 96676 14714
rect 96380 14660 96436 14662
rect 96460 14660 96516 14662
rect 96540 14660 96596 14662
rect 96620 14660 96676 14662
rect 96380 13626 96436 13628
rect 96460 13626 96516 13628
rect 96540 13626 96596 13628
rect 96620 13626 96676 13628
rect 96380 13574 96426 13626
rect 96426 13574 96436 13626
rect 96460 13574 96490 13626
rect 96490 13574 96502 13626
rect 96502 13574 96516 13626
rect 96540 13574 96554 13626
rect 96554 13574 96566 13626
rect 96566 13574 96596 13626
rect 96620 13574 96630 13626
rect 96630 13574 96676 13626
rect 96380 13572 96436 13574
rect 96460 13572 96516 13574
rect 96540 13572 96596 13574
rect 96620 13572 96676 13574
rect 96380 12538 96436 12540
rect 96460 12538 96516 12540
rect 96540 12538 96596 12540
rect 96620 12538 96676 12540
rect 96380 12486 96426 12538
rect 96426 12486 96436 12538
rect 96460 12486 96490 12538
rect 96490 12486 96502 12538
rect 96502 12486 96516 12538
rect 96540 12486 96554 12538
rect 96554 12486 96566 12538
rect 96566 12486 96596 12538
rect 96620 12486 96630 12538
rect 96630 12486 96676 12538
rect 96380 12484 96436 12486
rect 96460 12484 96516 12486
rect 96540 12484 96596 12486
rect 96620 12484 96676 12486
rect 96380 11450 96436 11452
rect 96460 11450 96516 11452
rect 96540 11450 96596 11452
rect 96620 11450 96676 11452
rect 96380 11398 96426 11450
rect 96426 11398 96436 11450
rect 96460 11398 96490 11450
rect 96490 11398 96502 11450
rect 96502 11398 96516 11450
rect 96540 11398 96554 11450
rect 96554 11398 96566 11450
rect 96566 11398 96596 11450
rect 96620 11398 96630 11450
rect 96630 11398 96676 11450
rect 96380 11396 96436 11398
rect 96460 11396 96516 11398
rect 96540 11396 96596 11398
rect 96620 11396 96676 11398
rect 96380 10362 96436 10364
rect 96460 10362 96516 10364
rect 96540 10362 96596 10364
rect 96620 10362 96676 10364
rect 96380 10310 96426 10362
rect 96426 10310 96436 10362
rect 96460 10310 96490 10362
rect 96490 10310 96502 10362
rect 96502 10310 96516 10362
rect 96540 10310 96554 10362
rect 96554 10310 96566 10362
rect 96566 10310 96596 10362
rect 96620 10310 96630 10362
rect 96630 10310 96676 10362
rect 96380 10308 96436 10310
rect 96460 10308 96516 10310
rect 96540 10308 96596 10310
rect 96620 10308 96676 10310
rect 96380 9274 96436 9276
rect 96460 9274 96516 9276
rect 96540 9274 96596 9276
rect 96620 9274 96676 9276
rect 96380 9222 96426 9274
rect 96426 9222 96436 9274
rect 96460 9222 96490 9274
rect 96490 9222 96502 9274
rect 96502 9222 96516 9274
rect 96540 9222 96554 9274
rect 96554 9222 96566 9274
rect 96566 9222 96596 9274
rect 96620 9222 96630 9274
rect 96630 9222 96676 9274
rect 96380 9220 96436 9222
rect 96460 9220 96516 9222
rect 96540 9220 96596 9222
rect 96620 9220 96676 9222
rect 96380 8186 96436 8188
rect 96460 8186 96516 8188
rect 96540 8186 96596 8188
rect 96620 8186 96676 8188
rect 96380 8134 96426 8186
rect 96426 8134 96436 8186
rect 96460 8134 96490 8186
rect 96490 8134 96502 8186
rect 96502 8134 96516 8186
rect 96540 8134 96554 8186
rect 96554 8134 96566 8186
rect 96566 8134 96596 8186
rect 96620 8134 96630 8186
rect 96630 8134 96676 8186
rect 96380 8132 96436 8134
rect 96460 8132 96516 8134
rect 96540 8132 96596 8134
rect 96620 8132 96676 8134
rect 96380 7098 96436 7100
rect 96460 7098 96516 7100
rect 96540 7098 96596 7100
rect 96620 7098 96676 7100
rect 96380 7046 96426 7098
rect 96426 7046 96436 7098
rect 96460 7046 96490 7098
rect 96490 7046 96502 7098
rect 96502 7046 96516 7098
rect 96540 7046 96554 7098
rect 96554 7046 96566 7098
rect 96566 7046 96596 7098
rect 96620 7046 96630 7098
rect 96630 7046 96676 7098
rect 96380 7044 96436 7046
rect 96460 7044 96516 7046
rect 96540 7044 96596 7046
rect 96620 7044 96676 7046
rect 96380 6010 96436 6012
rect 96460 6010 96516 6012
rect 96540 6010 96596 6012
rect 96620 6010 96676 6012
rect 96380 5958 96426 6010
rect 96426 5958 96436 6010
rect 96460 5958 96490 6010
rect 96490 5958 96502 6010
rect 96502 5958 96516 6010
rect 96540 5958 96554 6010
rect 96554 5958 96566 6010
rect 96566 5958 96596 6010
rect 96620 5958 96630 6010
rect 96630 5958 96676 6010
rect 96380 5956 96436 5958
rect 96460 5956 96516 5958
rect 96540 5956 96596 5958
rect 96620 5956 96676 5958
rect 96380 4922 96436 4924
rect 96460 4922 96516 4924
rect 96540 4922 96596 4924
rect 96620 4922 96676 4924
rect 96380 4870 96426 4922
rect 96426 4870 96436 4922
rect 96460 4870 96490 4922
rect 96490 4870 96502 4922
rect 96502 4870 96516 4922
rect 96540 4870 96554 4922
rect 96554 4870 96566 4922
rect 96566 4870 96596 4922
rect 96620 4870 96630 4922
rect 96630 4870 96676 4922
rect 96380 4868 96436 4870
rect 96460 4868 96516 4870
rect 96540 4868 96596 4870
rect 96620 4868 96676 4870
rect 96380 3834 96436 3836
rect 96460 3834 96516 3836
rect 96540 3834 96596 3836
rect 96620 3834 96676 3836
rect 96380 3782 96426 3834
rect 96426 3782 96436 3834
rect 96460 3782 96490 3834
rect 96490 3782 96502 3834
rect 96502 3782 96516 3834
rect 96540 3782 96554 3834
rect 96554 3782 96566 3834
rect 96566 3782 96596 3834
rect 96620 3782 96630 3834
rect 96630 3782 96676 3834
rect 96380 3780 96436 3782
rect 96460 3780 96516 3782
rect 96540 3780 96596 3782
rect 96620 3780 96676 3782
rect 96380 2746 96436 2748
rect 96460 2746 96516 2748
rect 96540 2746 96596 2748
rect 96620 2746 96676 2748
rect 96380 2694 96426 2746
rect 96426 2694 96436 2746
rect 96460 2694 96490 2746
rect 96490 2694 96502 2746
rect 96502 2694 96516 2746
rect 96540 2694 96554 2746
rect 96554 2694 96566 2746
rect 96566 2694 96596 2746
rect 96620 2694 96630 2746
rect 96630 2694 96676 2746
rect 96380 2692 96436 2694
rect 96460 2692 96516 2694
rect 96540 2692 96596 2694
rect 96620 2692 96676 2694
rect 97630 3052 97686 3088
rect 97630 3032 97632 3052
rect 97632 3032 97684 3052
rect 97684 3032 97686 3052
rect 97538 2352 97594 2408
rect 111740 35930 111796 35932
rect 111820 35930 111876 35932
rect 111900 35930 111956 35932
rect 111980 35930 112036 35932
rect 111740 35878 111786 35930
rect 111786 35878 111796 35930
rect 111820 35878 111850 35930
rect 111850 35878 111862 35930
rect 111862 35878 111876 35930
rect 111900 35878 111914 35930
rect 111914 35878 111926 35930
rect 111926 35878 111956 35930
rect 111980 35878 111990 35930
rect 111990 35878 112036 35930
rect 111740 35876 111796 35878
rect 111820 35876 111876 35878
rect 111900 35876 111956 35878
rect 111980 35876 112036 35878
rect 111740 34842 111796 34844
rect 111820 34842 111876 34844
rect 111900 34842 111956 34844
rect 111980 34842 112036 34844
rect 111740 34790 111786 34842
rect 111786 34790 111796 34842
rect 111820 34790 111850 34842
rect 111850 34790 111862 34842
rect 111862 34790 111876 34842
rect 111900 34790 111914 34842
rect 111914 34790 111926 34842
rect 111926 34790 111956 34842
rect 111980 34790 111990 34842
rect 111990 34790 112036 34842
rect 111740 34788 111796 34790
rect 111820 34788 111876 34790
rect 111900 34788 111956 34790
rect 111980 34788 112036 34790
rect 111740 33754 111796 33756
rect 111820 33754 111876 33756
rect 111900 33754 111956 33756
rect 111980 33754 112036 33756
rect 111740 33702 111786 33754
rect 111786 33702 111796 33754
rect 111820 33702 111850 33754
rect 111850 33702 111862 33754
rect 111862 33702 111876 33754
rect 111900 33702 111914 33754
rect 111914 33702 111926 33754
rect 111926 33702 111956 33754
rect 111980 33702 111990 33754
rect 111990 33702 112036 33754
rect 111740 33700 111796 33702
rect 111820 33700 111876 33702
rect 111900 33700 111956 33702
rect 111980 33700 112036 33702
rect 98458 2624 98514 2680
rect 98734 2488 98790 2544
rect 99654 3168 99710 3224
rect 99562 2624 99618 2680
rect 100574 3168 100630 3224
rect 100758 3032 100814 3088
rect 105450 2488 105506 2544
rect 105726 2388 105728 2408
rect 105728 2388 105780 2408
rect 105780 2388 105782 2408
rect 105726 2352 105782 2388
rect 111740 32666 111796 32668
rect 111820 32666 111876 32668
rect 111900 32666 111956 32668
rect 111980 32666 112036 32668
rect 111740 32614 111786 32666
rect 111786 32614 111796 32666
rect 111820 32614 111850 32666
rect 111850 32614 111862 32666
rect 111862 32614 111876 32666
rect 111900 32614 111914 32666
rect 111914 32614 111926 32666
rect 111926 32614 111956 32666
rect 111980 32614 111990 32666
rect 111990 32614 112036 32666
rect 111740 32612 111796 32614
rect 111820 32612 111876 32614
rect 111900 32612 111956 32614
rect 111980 32612 112036 32614
rect 111740 31578 111796 31580
rect 111820 31578 111876 31580
rect 111900 31578 111956 31580
rect 111980 31578 112036 31580
rect 111740 31526 111786 31578
rect 111786 31526 111796 31578
rect 111820 31526 111850 31578
rect 111850 31526 111862 31578
rect 111862 31526 111876 31578
rect 111900 31526 111914 31578
rect 111914 31526 111926 31578
rect 111926 31526 111956 31578
rect 111980 31526 111990 31578
rect 111990 31526 112036 31578
rect 111740 31524 111796 31526
rect 111820 31524 111876 31526
rect 111900 31524 111956 31526
rect 111980 31524 112036 31526
rect 111740 30490 111796 30492
rect 111820 30490 111876 30492
rect 111900 30490 111956 30492
rect 111980 30490 112036 30492
rect 111740 30438 111786 30490
rect 111786 30438 111796 30490
rect 111820 30438 111850 30490
rect 111850 30438 111862 30490
rect 111862 30438 111876 30490
rect 111900 30438 111914 30490
rect 111914 30438 111926 30490
rect 111926 30438 111956 30490
rect 111980 30438 111990 30490
rect 111990 30438 112036 30490
rect 111740 30436 111796 30438
rect 111820 30436 111876 30438
rect 111900 30436 111956 30438
rect 111980 30436 112036 30438
rect 111740 29402 111796 29404
rect 111820 29402 111876 29404
rect 111900 29402 111956 29404
rect 111980 29402 112036 29404
rect 111740 29350 111786 29402
rect 111786 29350 111796 29402
rect 111820 29350 111850 29402
rect 111850 29350 111862 29402
rect 111862 29350 111876 29402
rect 111900 29350 111914 29402
rect 111914 29350 111926 29402
rect 111926 29350 111956 29402
rect 111980 29350 111990 29402
rect 111990 29350 112036 29402
rect 111740 29348 111796 29350
rect 111820 29348 111876 29350
rect 111900 29348 111956 29350
rect 111980 29348 112036 29350
rect 111740 28314 111796 28316
rect 111820 28314 111876 28316
rect 111900 28314 111956 28316
rect 111980 28314 112036 28316
rect 111740 28262 111786 28314
rect 111786 28262 111796 28314
rect 111820 28262 111850 28314
rect 111850 28262 111862 28314
rect 111862 28262 111876 28314
rect 111900 28262 111914 28314
rect 111914 28262 111926 28314
rect 111926 28262 111956 28314
rect 111980 28262 111990 28314
rect 111990 28262 112036 28314
rect 111740 28260 111796 28262
rect 111820 28260 111876 28262
rect 111900 28260 111956 28262
rect 111980 28260 112036 28262
rect 111740 27226 111796 27228
rect 111820 27226 111876 27228
rect 111900 27226 111956 27228
rect 111980 27226 112036 27228
rect 111740 27174 111786 27226
rect 111786 27174 111796 27226
rect 111820 27174 111850 27226
rect 111850 27174 111862 27226
rect 111862 27174 111876 27226
rect 111900 27174 111914 27226
rect 111914 27174 111926 27226
rect 111926 27174 111956 27226
rect 111980 27174 111990 27226
rect 111990 27174 112036 27226
rect 111740 27172 111796 27174
rect 111820 27172 111876 27174
rect 111900 27172 111956 27174
rect 111980 27172 112036 27174
rect 111740 26138 111796 26140
rect 111820 26138 111876 26140
rect 111900 26138 111956 26140
rect 111980 26138 112036 26140
rect 111740 26086 111786 26138
rect 111786 26086 111796 26138
rect 111820 26086 111850 26138
rect 111850 26086 111862 26138
rect 111862 26086 111876 26138
rect 111900 26086 111914 26138
rect 111914 26086 111926 26138
rect 111926 26086 111956 26138
rect 111980 26086 111990 26138
rect 111990 26086 112036 26138
rect 111740 26084 111796 26086
rect 111820 26084 111876 26086
rect 111900 26084 111956 26086
rect 111980 26084 112036 26086
rect 111740 25050 111796 25052
rect 111820 25050 111876 25052
rect 111900 25050 111956 25052
rect 111980 25050 112036 25052
rect 111740 24998 111786 25050
rect 111786 24998 111796 25050
rect 111820 24998 111850 25050
rect 111850 24998 111862 25050
rect 111862 24998 111876 25050
rect 111900 24998 111914 25050
rect 111914 24998 111926 25050
rect 111926 24998 111956 25050
rect 111980 24998 111990 25050
rect 111990 24998 112036 25050
rect 111740 24996 111796 24998
rect 111820 24996 111876 24998
rect 111900 24996 111956 24998
rect 111980 24996 112036 24998
rect 111740 23962 111796 23964
rect 111820 23962 111876 23964
rect 111900 23962 111956 23964
rect 111980 23962 112036 23964
rect 111740 23910 111786 23962
rect 111786 23910 111796 23962
rect 111820 23910 111850 23962
rect 111850 23910 111862 23962
rect 111862 23910 111876 23962
rect 111900 23910 111914 23962
rect 111914 23910 111926 23962
rect 111926 23910 111956 23962
rect 111980 23910 111990 23962
rect 111990 23910 112036 23962
rect 111740 23908 111796 23910
rect 111820 23908 111876 23910
rect 111900 23908 111956 23910
rect 111980 23908 112036 23910
rect 111740 22874 111796 22876
rect 111820 22874 111876 22876
rect 111900 22874 111956 22876
rect 111980 22874 112036 22876
rect 111740 22822 111786 22874
rect 111786 22822 111796 22874
rect 111820 22822 111850 22874
rect 111850 22822 111862 22874
rect 111862 22822 111876 22874
rect 111900 22822 111914 22874
rect 111914 22822 111926 22874
rect 111926 22822 111956 22874
rect 111980 22822 111990 22874
rect 111990 22822 112036 22874
rect 111740 22820 111796 22822
rect 111820 22820 111876 22822
rect 111900 22820 111956 22822
rect 111980 22820 112036 22822
rect 111740 21786 111796 21788
rect 111820 21786 111876 21788
rect 111900 21786 111956 21788
rect 111980 21786 112036 21788
rect 111740 21734 111786 21786
rect 111786 21734 111796 21786
rect 111820 21734 111850 21786
rect 111850 21734 111862 21786
rect 111862 21734 111876 21786
rect 111900 21734 111914 21786
rect 111914 21734 111926 21786
rect 111926 21734 111956 21786
rect 111980 21734 111990 21786
rect 111990 21734 112036 21786
rect 111740 21732 111796 21734
rect 111820 21732 111876 21734
rect 111900 21732 111956 21734
rect 111980 21732 112036 21734
rect 111740 20698 111796 20700
rect 111820 20698 111876 20700
rect 111900 20698 111956 20700
rect 111980 20698 112036 20700
rect 111740 20646 111786 20698
rect 111786 20646 111796 20698
rect 111820 20646 111850 20698
rect 111850 20646 111862 20698
rect 111862 20646 111876 20698
rect 111900 20646 111914 20698
rect 111914 20646 111926 20698
rect 111926 20646 111956 20698
rect 111980 20646 111990 20698
rect 111990 20646 112036 20698
rect 111740 20644 111796 20646
rect 111820 20644 111876 20646
rect 111900 20644 111956 20646
rect 111980 20644 112036 20646
rect 111740 19610 111796 19612
rect 111820 19610 111876 19612
rect 111900 19610 111956 19612
rect 111980 19610 112036 19612
rect 111740 19558 111786 19610
rect 111786 19558 111796 19610
rect 111820 19558 111850 19610
rect 111850 19558 111862 19610
rect 111862 19558 111876 19610
rect 111900 19558 111914 19610
rect 111914 19558 111926 19610
rect 111926 19558 111956 19610
rect 111980 19558 111990 19610
rect 111990 19558 112036 19610
rect 111740 19556 111796 19558
rect 111820 19556 111876 19558
rect 111900 19556 111956 19558
rect 111980 19556 112036 19558
rect 111740 18522 111796 18524
rect 111820 18522 111876 18524
rect 111900 18522 111956 18524
rect 111980 18522 112036 18524
rect 111740 18470 111786 18522
rect 111786 18470 111796 18522
rect 111820 18470 111850 18522
rect 111850 18470 111862 18522
rect 111862 18470 111876 18522
rect 111900 18470 111914 18522
rect 111914 18470 111926 18522
rect 111926 18470 111956 18522
rect 111980 18470 111990 18522
rect 111990 18470 112036 18522
rect 111740 18468 111796 18470
rect 111820 18468 111876 18470
rect 111900 18468 111956 18470
rect 111980 18468 112036 18470
rect 111740 17434 111796 17436
rect 111820 17434 111876 17436
rect 111900 17434 111956 17436
rect 111980 17434 112036 17436
rect 111740 17382 111786 17434
rect 111786 17382 111796 17434
rect 111820 17382 111850 17434
rect 111850 17382 111862 17434
rect 111862 17382 111876 17434
rect 111900 17382 111914 17434
rect 111914 17382 111926 17434
rect 111926 17382 111956 17434
rect 111980 17382 111990 17434
rect 111990 17382 112036 17434
rect 111740 17380 111796 17382
rect 111820 17380 111876 17382
rect 111900 17380 111956 17382
rect 111980 17380 112036 17382
rect 111740 16346 111796 16348
rect 111820 16346 111876 16348
rect 111900 16346 111956 16348
rect 111980 16346 112036 16348
rect 111740 16294 111786 16346
rect 111786 16294 111796 16346
rect 111820 16294 111850 16346
rect 111850 16294 111862 16346
rect 111862 16294 111876 16346
rect 111900 16294 111914 16346
rect 111914 16294 111926 16346
rect 111926 16294 111956 16346
rect 111980 16294 111990 16346
rect 111990 16294 112036 16346
rect 111740 16292 111796 16294
rect 111820 16292 111876 16294
rect 111900 16292 111956 16294
rect 111980 16292 112036 16294
rect 111740 15258 111796 15260
rect 111820 15258 111876 15260
rect 111900 15258 111956 15260
rect 111980 15258 112036 15260
rect 111740 15206 111786 15258
rect 111786 15206 111796 15258
rect 111820 15206 111850 15258
rect 111850 15206 111862 15258
rect 111862 15206 111876 15258
rect 111900 15206 111914 15258
rect 111914 15206 111926 15258
rect 111926 15206 111956 15258
rect 111980 15206 111990 15258
rect 111990 15206 112036 15258
rect 111740 15204 111796 15206
rect 111820 15204 111876 15206
rect 111900 15204 111956 15206
rect 111980 15204 112036 15206
rect 111740 14170 111796 14172
rect 111820 14170 111876 14172
rect 111900 14170 111956 14172
rect 111980 14170 112036 14172
rect 111740 14118 111786 14170
rect 111786 14118 111796 14170
rect 111820 14118 111850 14170
rect 111850 14118 111862 14170
rect 111862 14118 111876 14170
rect 111900 14118 111914 14170
rect 111914 14118 111926 14170
rect 111926 14118 111956 14170
rect 111980 14118 111990 14170
rect 111990 14118 112036 14170
rect 111740 14116 111796 14118
rect 111820 14116 111876 14118
rect 111900 14116 111956 14118
rect 111980 14116 112036 14118
rect 111740 13082 111796 13084
rect 111820 13082 111876 13084
rect 111900 13082 111956 13084
rect 111980 13082 112036 13084
rect 111740 13030 111786 13082
rect 111786 13030 111796 13082
rect 111820 13030 111850 13082
rect 111850 13030 111862 13082
rect 111862 13030 111876 13082
rect 111900 13030 111914 13082
rect 111914 13030 111926 13082
rect 111926 13030 111956 13082
rect 111980 13030 111990 13082
rect 111990 13030 112036 13082
rect 111740 13028 111796 13030
rect 111820 13028 111876 13030
rect 111900 13028 111956 13030
rect 111980 13028 112036 13030
rect 111740 11994 111796 11996
rect 111820 11994 111876 11996
rect 111900 11994 111956 11996
rect 111980 11994 112036 11996
rect 111740 11942 111786 11994
rect 111786 11942 111796 11994
rect 111820 11942 111850 11994
rect 111850 11942 111862 11994
rect 111862 11942 111876 11994
rect 111900 11942 111914 11994
rect 111914 11942 111926 11994
rect 111926 11942 111956 11994
rect 111980 11942 111990 11994
rect 111990 11942 112036 11994
rect 111740 11940 111796 11942
rect 111820 11940 111876 11942
rect 111900 11940 111956 11942
rect 111980 11940 112036 11942
rect 111740 10906 111796 10908
rect 111820 10906 111876 10908
rect 111900 10906 111956 10908
rect 111980 10906 112036 10908
rect 111740 10854 111786 10906
rect 111786 10854 111796 10906
rect 111820 10854 111850 10906
rect 111850 10854 111862 10906
rect 111862 10854 111876 10906
rect 111900 10854 111914 10906
rect 111914 10854 111926 10906
rect 111926 10854 111956 10906
rect 111980 10854 111990 10906
rect 111990 10854 112036 10906
rect 111740 10852 111796 10854
rect 111820 10852 111876 10854
rect 111900 10852 111956 10854
rect 111980 10852 112036 10854
rect 111740 9818 111796 9820
rect 111820 9818 111876 9820
rect 111900 9818 111956 9820
rect 111980 9818 112036 9820
rect 111740 9766 111786 9818
rect 111786 9766 111796 9818
rect 111820 9766 111850 9818
rect 111850 9766 111862 9818
rect 111862 9766 111876 9818
rect 111900 9766 111914 9818
rect 111914 9766 111926 9818
rect 111926 9766 111956 9818
rect 111980 9766 111990 9818
rect 111990 9766 112036 9818
rect 111740 9764 111796 9766
rect 111820 9764 111876 9766
rect 111900 9764 111956 9766
rect 111980 9764 112036 9766
rect 111740 8730 111796 8732
rect 111820 8730 111876 8732
rect 111900 8730 111956 8732
rect 111980 8730 112036 8732
rect 111740 8678 111786 8730
rect 111786 8678 111796 8730
rect 111820 8678 111850 8730
rect 111850 8678 111862 8730
rect 111862 8678 111876 8730
rect 111900 8678 111914 8730
rect 111914 8678 111926 8730
rect 111926 8678 111956 8730
rect 111980 8678 111990 8730
rect 111990 8678 112036 8730
rect 111740 8676 111796 8678
rect 111820 8676 111876 8678
rect 111900 8676 111956 8678
rect 111980 8676 112036 8678
rect 111740 7642 111796 7644
rect 111820 7642 111876 7644
rect 111900 7642 111956 7644
rect 111980 7642 112036 7644
rect 111740 7590 111786 7642
rect 111786 7590 111796 7642
rect 111820 7590 111850 7642
rect 111850 7590 111862 7642
rect 111862 7590 111876 7642
rect 111900 7590 111914 7642
rect 111914 7590 111926 7642
rect 111926 7590 111956 7642
rect 111980 7590 111990 7642
rect 111990 7590 112036 7642
rect 111740 7588 111796 7590
rect 111820 7588 111876 7590
rect 111900 7588 111956 7590
rect 111980 7588 112036 7590
rect 111740 6554 111796 6556
rect 111820 6554 111876 6556
rect 111900 6554 111956 6556
rect 111980 6554 112036 6556
rect 111740 6502 111786 6554
rect 111786 6502 111796 6554
rect 111820 6502 111850 6554
rect 111850 6502 111862 6554
rect 111862 6502 111876 6554
rect 111900 6502 111914 6554
rect 111914 6502 111926 6554
rect 111926 6502 111956 6554
rect 111980 6502 111990 6554
rect 111990 6502 112036 6554
rect 111740 6500 111796 6502
rect 111820 6500 111876 6502
rect 111900 6500 111956 6502
rect 111980 6500 112036 6502
rect 111740 5466 111796 5468
rect 111820 5466 111876 5468
rect 111900 5466 111956 5468
rect 111980 5466 112036 5468
rect 111740 5414 111786 5466
rect 111786 5414 111796 5466
rect 111820 5414 111850 5466
rect 111850 5414 111862 5466
rect 111862 5414 111876 5466
rect 111900 5414 111914 5466
rect 111914 5414 111926 5466
rect 111926 5414 111956 5466
rect 111980 5414 111990 5466
rect 111990 5414 112036 5466
rect 111740 5412 111796 5414
rect 111820 5412 111876 5414
rect 111900 5412 111956 5414
rect 111980 5412 112036 5414
rect 111740 4378 111796 4380
rect 111820 4378 111876 4380
rect 111900 4378 111956 4380
rect 111980 4378 112036 4380
rect 111740 4326 111786 4378
rect 111786 4326 111796 4378
rect 111820 4326 111850 4378
rect 111850 4326 111862 4378
rect 111862 4326 111876 4378
rect 111900 4326 111914 4378
rect 111914 4326 111926 4378
rect 111926 4326 111956 4378
rect 111980 4326 111990 4378
rect 111990 4326 112036 4378
rect 111740 4324 111796 4326
rect 111820 4324 111876 4326
rect 111900 4324 111956 4326
rect 111980 4324 112036 4326
rect 111740 3290 111796 3292
rect 111820 3290 111876 3292
rect 111900 3290 111956 3292
rect 111980 3290 112036 3292
rect 111740 3238 111786 3290
rect 111786 3238 111796 3290
rect 111820 3238 111850 3290
rect 111850 3238 111862 3290
rect 111862 3238 111876 3290
rect 111900 3238 111914 3290
rect 111914 3238 111926 3290
rect 111926 3238 111956 3290
rect 111980 3238 111990 3290
rect 111990 3238 112036 3290
rect 111740 3236 111796 3238
rect 111820 3236 111876 3238
rect 111900 3236 111956 3238
rect 111980 3236 112036 3238
rect 111740 2202 111796 2204
rect 111820 2202 111876 2204
rect 111900 2202 111956 2204
rect 111980 2202 112036 2204
rect 111740 2150 111786 2202
rect 111786 2150 111796 2202
rect 111820 2150 111850 2202
rect 111850 2150 111862 2202
rect 111862 2150 111876 2202
rect 111900 2150 111914 2202
rect 111914 2150 111926 2202
rect 111926 2150 111956 2202
rect 111980 2150 111990 2202
rect 111990 2150 112036 2202
rect 111740 2148 111796 2150
rect 111820 2148 111876 2150
rect 111900 2148 111956 2150
rect 111980 2148 112036 2150
rect 117226 38528 117282 38584
rect 118054 37576 118110 37632
rect 117226 3168 117282 3224
rect 118054 36644 118110 36680
rect 118054 36624 118056 36644
rect 118056 36624 118108 36644
rect 118108 36624 118110 36644
rect 118054 35672 118110 35728
rect 118054 34720 118110 34776
rect 118054 33904 118110 33960
rect 118054 32952 118110 33008
rect 118054 32000 118110 32056
rect 118054 31084 118056 31104
rect 118056 31084 118108 31104
rect 118108 31084 118110 31104
rect 118054 31048 118110 31084
rect 118054 30116 118110 30152
rect 118054 30096 118056 30116
rect 118056 30096 118108 30116
rect 118108 30096 118110 30116
rect 118054 29144 118110 29200
rect 118054 28364 118056 28384
rect 118056 28364 118108 28384
rect 118108 28364 118110 28384
rect 118054 28328 118110 28364
rect 118054 27376 118110 27432
rect 118054 26424 118110 26480
rect 118054 25472 118110 25528
rect 118054 24556 118056 24576
rect 118056 24556 118108 24576
rect 118108 24556 118110 24576
rect 118054 24520 118110 24556
rect 118054 23588 118110 23624
rect 118054 23568 118056 23588
rect 118056 23568 118108 23588
rect 118108 23568 118110 23588
rect 118054 22752 118110 22808
rect 118054 21836 118056 21856
rect 118056 21836 118108 21856
rect 118108 21836 118110 21856
rect 118054 21800 118110 21836
rect 118054 20848 118110 20904
rect 118054 19896 118110 19952
rect 118054 18944 118110 19000
rect 118054 18028 118056 18048
rect 118056 18028 118108 18048
rect 118108 18028 118110 18048
rect 118054 17992 118110 18028
rect 118054 17176 118110 17232
rect 117778 9696 117834 9752
rect 117778 8744 117834 8800
rect 117778 7812 117834 7848
rect 117778 7792 117780 7812
rect 117780 7792 117832 7812
rect 117832 7792 117834 7812
rect 117778 6840 117834 6896
rect 117778 6024 117834 6080
rect 117134 2216 117190 2272
rect 117778 5072 117834 5128
rect 117778 4120 117834 4176
rect 118054 16224 118110 16280
rect 118054 15308 118056 15328
rect 118056 15308 118108 15328
rect 118108 15308 118110 15328
rect 118054 15272 118110 15308
rect 118054 14320 118110 14376
rect 118054 13368 118110 13424
rect 118054 12416 118110 12472
rect 118054 11620 118110 11656
rect 118054 11600 118056 11620
rect 118056 11600 118108 11620
rect 118108 11600 118110 11620
rect 118054 10648 118110 10704
rect 117778 1264 117834 1320
rect 116490 448 116546 504
<< metal3 >>
rect 117129 39538 117195 39541
rect 119200 39538 120000 39568
rect 117129 39536 120000 39538
rect 117129 39480 117134 39536
rect 117190 39480 120000 39536
rect 117129 39478 120000 39480
rect 117129 39475 117195 39478
rect 119200 39448 120000 39478
rect 117221 38586 117287 38589
rect 119200 38586 120000 38616
rect 117221 38584 120000 38586
rect 117221 38528 117226 38584
rect 117282 38528 120000 38584
rect 117221 38526 120000 38528
rect 117221 38523 117287 38526
rect 119200 38496 120000 38526
rect 118049 37634 118115 37637
rect 119200 37634 120000 37664
rect 118049 37632 120000 37634
rect 118049 37576 118054 37632
rect 118110 37576 120000 37632
rect 118049 37574 120000 37576
rect 118049 37571 118115 37574
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 65648 37568 65968 37569
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 37503 65968 37504
rect 96368 37568 96688 37569
rect 96368 37504 96376 37568
rect 96440 37504 96456 37568
rect 96520 37504 96536 37568
rect 96600 37504 96616 37568
rect 96680 37504 96688 37568
rect 119200 37544 120000 37574
rect 96368 37503 96688 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 81008 37024 81328 37025
rect 81008 36960 81016 37024
rect 81080 36960 81096 37024
rect 81160 36960 81176 37024
rect 81240 36960 81256 37024
rect 81320 36960 81328 37024
rect 81008 36959 81328 36960
rect 111728 37024 112048 37025
rect 111728 36960 111736 37024
rect 111800 36960 111816 37024
rect 111880 36960 111896 37024
rect 111960 36960 111976 37024
rect 112040 36960 112048 37024
rect 111728 36959 112048 36960
rect 118049 36682 118115 36685
rect 119200 36682 120000 36712
rect 118049 36680 120000 36682
rect 118049 36624 118054 36680
rect 118110 36624 120000 36680
rect 118049 36622 120000 36624
rect 118049 36619 118115 36622
rect 119200 36592 120000 36622
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 65648 36480 65968 36481
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 36415 65968 36416
rect 96368 36480 96688 36481
rect 96368 36416 96376 36480
rect 96440 36416 96456 36480
rect 96520 36416 96536 36480
rect 96600 36416 96616 36480
rect 96680 36416 96688 36480
rect 96368 36415 96688 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 81008 35936 81328 35937
rect 81008 35872 81016 35936
rect 81080 35872 81096 35936
rect 81160 35872 81176 35936
rect 81240 35872 81256 35936
rect 81320 35872 81328 35936
rect 81008 35871 81328 35872
rect 111728 35936 112048 35937
rect 111728 35872 111736 35936
rect 111800 35872 111816 35936
rect 111880 35872 111896 35936
rect 111960 35872 111976 35936
rect 112040 35872 112048 35936
rect 111728 35871 112048 35872
rect 118049 35730 118115 35733
rect 119200 35730 120000 35760
rect 118049 35728 120000 35730
rect 118049 35672 118054 35728
rect 118110 35672 120000 35728
rect 118049 35670 120000 35672
rect 118049 35667 118115 35670
rect 119200 35640 120000 35670
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 65648 35392 65968 35393
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 35327 65968 35328
rect 96368 35392 96688 35393
rect 96368 35328 96376 35392
rect 96440 35328 96456 35392
rect 96520 35328 96536 35392
rect 96600 35328 96616 35392
rect 96680 35328 96688 35392
rect 96368 35327 96688 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 81008 34848 81328 34849
rect 81008 34784 81016 34848
rect 81080 34784 81096 34848
rect 81160 34784 81176 34848
rect 81240 34784 81256 34848
rect 81320 34784 81328 34848
rect 81008 34783 81328 34784
rect 111728 34848 112048 34849
rect 111728 34784 111736 34848
rect 111800 34784 111816 34848
rect 111880 34784 111896 34848
rect 111960 34784 111976 34848
rect 112040 34784 112048 34848
rect 111728 34783 112048 34784
rect 118049 34778 118115 34781
rect 119200 34778 120000 34808
rect 118049 34776 120000 34778
rect 118049 34720 118054 34776
rect 118110 34720 120000 34776
rect 118049 34718 120000 34720
rect 118049 34715 118115 34718
rect 119200 34688 120000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 65648 34304 65968 34305
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 34239 65968 34240
rect 96368 34304 96688 34305
rect 96368 34240 96376 34304
rect 96440 34240 96456 34304
rect 96520 34240 96536 34304
rect 96600 34240 96616 34304
rect 96680 34240 96688 34304
rect 96368 34239 96688 34240
rect 118049 33962 118115 33965
rect 119200 33962 120000 33992
rect 118049 33960 120000 33962
rect 118049 33904 118054 33960
rect 118110 33904 120000 33960
rect 118049 33902 120000 33904
rect 118049 33899 118115 33902
rect 119200 33872 120000 33902
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 81008 33760 81328 33761
rect 81008 33696 81016 33760
rect 81080 33696 81096 33760
rect 81160 33696 81176 33760
rect 81240 33696 81256 33760
rect 81320 33696 81328 33760
rect 81008 33695 81328 33696
rect 111728 33760 112048 33761
rect 111728 33696 111736 33760
rect 111800 33696 111816 33760
rect 111880 33696 111896 33760
rect 111960 33696 111976 33760
rect 112040 33696 112048 33760
rect 111728 33695 112048 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 65648 33216 65968 33217
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 33151 65968 33152
rect 96368 33216 96688 33217
rect 96368 33152 96376 33216
rect 96440 33152 96456 33216
rect 96520 33152 96536 33216
rect 96600 33152 96616 33216
rect 96680 33152 96688 33216
rect 96368 33151 96688 33152
rect 118049 33010 118115 33013
rect 119200 33010 120000 33040
rect 118049 33008 120000 33010
rect 118049 32952 118054 33008
rect 118110 32952 120000 33008
rect 118049 32950 120000 32952
rect 118049 32947 118115 32950
rect 119200 32920 120000 32950
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 81008 32672 81328 32673
rect 81008 32608 81016 32672
rect 81080 32608 81096 32672
rect 81160 32608 81176 32672
rect 81240 32608 81256 32672
rect 81320 32608 81328 32672
rect 81008 32607 81328 32608
rect 111728 32672 112048 32673
rect 111728 32608 111736 32672
rect 111800 32608 111816 32672
rect 111880 32608 111896 32672
rect 111960 32608 111976 32672
rect 112040 32608 112048 32672
rect 111728 32607 112048 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 65648 32128 65968 32129
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 32063 65968 32064
rect 96368 32128 96688 32129
rect 96368 32064 96376 32128
rect 96440 32064 96456 32128
rect 96520 32064 96536 32128
rect 96600 32064 96616 32128
rect 96680 32064 96688 32128
rect 96368 32063 96688 32064
rect 118049 32058 118115 32061
rect 119200 32058 120000 32088
rect 118049 32056 120000 32058
rect 118049 32000 118054 32056
rect 118110 32000 120000 32056
rect 118049 31998 120000 32000
rect 118049 31995 118115 31998
rect 119200 31968 120000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 81008 31584 81328 31585
rect 81008 31520 81016 31584
rect 81080 31520 81096 31584
rect 81160 31520 81176 31584
rect 81240 31520 81256 31584
rect 81320 31520 81328 31584
rect 81008 31519 81328 31520
rect 111728 31584 112048 31585
rect 111728 31520 111736 31584
rect 111800 31520 111816 31584
rect 111880 31520 111896 31584
rect 111960 31520 111976 31584
rect 112040 31520 112048 31584
rect 111728 31519 112048 31520
rect 118049 31106 118115 31109
rect 119200 31106 120000 31136
rect 118049 31104 120000 31106
rect 118049 31048 118054 31104
rect 118110 31048 120000 31104
rect 118049 31046 120000 31048
rect 118049 31043 118115 31046
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 65648 31040 65968 31041
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 30975 65968 30976
rect 96368 31040 96688 31041
rect 96368 30976 96376 31040
rect 96440 30976 96456 31040
rect 96520 30976 96536 31040
rect 96600 30976 96616 31040
rect 96680 30976 96688 31040
rect 119200 31016 120000 31046
rect 96368 30975 96688 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 81008 30496 81328 30497
rect 81008 30432 81016 30496
rect 81080 30432 81096 30496
rect 81160 30432 81176 30496
rect 81240 30432 81256 30496
rect 81320 30432 81328 30496
rect 81008 30431 81328 30432
rect 111728 30496 112048 30497
rect 111728 30432 111736 30496
rect 111800 30432 111816 30496
rect 111880 30432 111896 30496
rect 111960 30432 111976 30496
rect 112040 30432 112048 30496
rect 111728 30431 112048 30432
rect 118049 30154 118115 30157
rect 119200 30154 120000 30184
rect 118049 30152 120000 30154
rect 118049 30096 118054 30152
rect 118110 30096 120000 30152
rect 118049 30094 120000 30096
rect 118049 30091 118115 30094
rect 119200 30064 120000 30094
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 65648 29952 65968 29953
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 29887 65968 29888
rect 96368 29952 96688 29953
rect 96368 29888 96376 29952
rect 96440 29888 96456 29952
rect 96520 29888 96536 29952
rect 96600 29888 96616 29952
rect 96680 29888 96688 29952
rect 96368 29887 96688 29888
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 81008 29408 81328 29409
rect 81008 29344 81016 29408
rect 81080 29344 81096 29408
rect 81160 29344 81176 29408
rect 81240 29344 81256 29408
rect 81320 29344 81328 29408
rect 81008 29343 81328 29344
rect 111728 29408 112048 29409
rect 111728 29344 111736 29408
rect 111800 29344 111816 29408
rect 111880 29344 111896 29408
rect 111960 29344 111976 29408
rect 112040 29344 112048 29408
rect 111728 29343 112048 29344
rect 118049 29202 118115 29205
rect 119200 29202 120000 29232
rect 118049 29200 120000 29202
rect 118049 29144 118054 29200
rect 118110 29144 120000 29200
rect 118049 29142 120000 29144
rect 118049 29139 118115 29142
rect 119200 29112 120000 29142
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 65648 28864 65968 28865
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 28799 65968 28800
rect 96368 28864 96688 28865
rect 96368 28800 96376 28864
rect 96440 28800 96456 28864
rect 96520 28800 96536 28864
rect 96600 28800 96616 28864
rect 96680 28800 96688 28864
rect 96368 28799 96688 28800
rect 118049 28386 118115 28389
rect 119200 28386 120000 28416
rect 118049 28384 120000 28386
rect 118049 28328 118054 28384
rect 118110 28328 120000 28384
rect 118049 28326 120000 28328
rect 118049 28323 118115 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 81008 28320 81328 28321
rect 81008 28256 81016 28320
rect 81080 28256 81096 28320
rect 81160 28256 81176 28320
rect 81240 28256 81256 28320
rect 81320 28256 81328 28320
rect 81008 28255 81328 28256
rect 111728 28320 112048 28321
rect 111728 28256 111736 28320
rect 111800 28256 111816 28320
rect 111880 28256 111896 28320
rect 111960 28256 111976 28320
rect 112040 28256 112048 28320
rect 119200 28296 120000 28326
rect 111728 28255 112048 28256
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 65648 27776 65968 27777
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 27711 65968 27712
rect 96368 27776 96688 27777
rect 96368 27712 96376 27776
rect 96440 27712 96456 27776
rect 96520 27712 96536 27776
rect 96600 27712 96616 27776
rect 96680 27712 96688 27776
rect 96368 27711 96688 27712
rect 118049 27434 118115 27437
rect 119200 27434 120000 27464
rect 118049 27432 120000 27434
rect 118049 27376 118054 27432
rect 118110 27376 120000 27432
rect 118049 27374 120000 27376
rect 118049 27371 118115 27374
rect 119200 27344 120000 27374
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 27167 50608 27168
rect 81008 27232 81328 27233
rect 81008 27168 81016 27232
rect 81080 27168 81096 27232
rect 81160 27168 81176 27232
rect 81240 27168 81256 27232
rect 81320 27168 81328 27232
rect 81008 27167 81328 27168
rect 111728 27232 112048 27233
rect 111728 27168 111736 27232
rect 111800 27168 111816 27232
rect 111880 27168 111896 27232
rect 111960 27168 111976 27232
rect 112040 27168 112048 27232
rect 111728 27167 112048 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 65648 26688 65968 26689
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 26623 65968 26624
rect 96368 26688 96688 26689
rect 96368 26624 96376 26688
rect 96440 26624 96456 26688
rect 96520 26624 96536 26688
rect 96600 26624 96616 26688
rect 96680 26624 96688 26688
rect 96368 26623 96688 26624
rect 118049 26482 118115 26485
rect 119200 26482 120000 26512
rect 118049 26480 120000 26482
rect 118049 26424 118054 26480
rect 118110 26424 120000 26480
rect 118049 26422 120000 26424
rect 118049 26419 118115 26422
rect 119200 26392 120000 26422
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 81008 26144 81328 26145
rect 81008 26080 81016 26144
rect 81080 26080 81096 26144
rect 81160 26080 81176 26144
rect 81240 26080 81256 26144
rect 81320 26080 81328 26144
rect 81008 26079 81328 26080
rect 111728 26144 112048 26145
rect 111728 26080 111736 26144
rect 111800 26080 111816 26144
rect 111880 26080 111896 26144
rect 111960 26080 111976 26144
rect 112040 26080 112048 26144
rect 111728 26079 112048 26080
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 65648 25600 65968 25601
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 25535 65968 25536
rect 96368 25600 96688 25601
rect 96368 25536 96376 25600
rect 96440 25536 96456 25600
rect 96520 25536 96536 25600
rect 96600 25536 96616 25600
rect 96680 25536 96688 25600
rect 96368 25535 96688 25536
rect 118049 25530 118115 25533
rect 119200 25530 120000 25560
rect 118049 25528 120000 25530
rect 118049 25472 118054 25528
rect 118110 25472 120000 25528
rect 118049 25470 120000 25472
rect 118049 25467 118115 25470
rect 119200 25440 120000 25470
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 81008 25056 81328 25057
rect 81008 24992 81016 25056
rect 81080 24992 81096 25056
rect 81160 24992 81176 25056
rect 81240 24992 81256 25056
rect 81320 24992 81328 25056
rect 81008 24991 81328 24992
rect 111728 25056 112048 25057
rect 111728 24992 111736 25056
rect 111800 24992 111816 25056
rect 111880 24992 111896 25056
rect 111960 24992 111976 25056
rect 112040 24992 112048 25056
rect 111728 24991 112048 24992
rect 118049 24578 118115 24581
rect 119200 24578 120000 24608
rect 118049 24576 120000 24578
rect 118049 24520 118054 24576
rect 118110 24520 120000 24576
rect 118049 24518 120000 24520
rect 118049 24515 118115 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 65648 24512 65968 24513
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 24447 65968 24448
rect 96368 24512 96688 24513
rect 96368 24448 96376 24512
rect 96440 24448 96456 24512
rect 96520 24448 96536 24512
rect 96600 24448 96616 24512
rect 96680 24448 96688 24512
rect 119200 24488 120000 24518
rect 96368 24447 96688 24448
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 81008 23968 81328 23969
rect 81008 23904 81016 23968
rect 81080 23904 81096 23968
rect 81160 23904 81176 23968
rect 81240 23904 81256 23968
rect 81320 23904 81328 23968
rect 81008 23903 81328 23904
rect 111728 23968 112048 23969
rect 111728 23904 111736 23968
rect 111800 23904 111816 23968
rect 111880 23904 111896 23968
rect 111960 23904 111976 23968
rect 112040 23904 112048 23968
rect 111728 23903 112048 23904
rect 118049 23626 118115 23629
rect 119200 23626 120000 23656
rect 118049 23624 120000 23626
rect 118049 23568 118054 23624
rect 118110 23568 120000 23624
rect 118049 23566 120000 23568
rect 118049 23563 118115 23566
rect 119200 23536 120000 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 65648 23424 65968 23425
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 23359 65968 23360
rect 96368 23424 96688 23425
rect 96368 23360 96376 23424
rect 96440 23360 96456 23424
rect 96520 23360 96536 23424
rect 96600 23360 96616 23424
rect 96680 23360 96688 23424
rect 96368 23359 96688 23360
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 81008 22880 81328 22881
rect 81008 22816 81016 22880
rect 81080 22816 81096 22880
rect 81160 22816 81176 22880
rect 81240 22816 81256 22880
rect 81320 22816 81328 22880
rect 81008 22815 81328 22816
rect 111728 22880 112048 22881
rect 111728 22816 111736 22880
rect 111800 22816 111816 22880
rect 111880 22816 111896 22880
rect 111960 22816 111976 22880
rect 112040 22816 112048 22880
rect 111728 22815 112048 22816
rect 118049 22810 118115 22813
rect 119200 22810 120000 22840
rect 118049 22808 120000 22810
rect 118049 22752 118054 22808
rect 118110 22752 120000 22808
rect 118049 22750 120000 22752
rect 118049 22747 118115 22750
rect 119200 22720 120000 22750
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 65648 22336 65968 22337
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 22271 65968 22272
rect 96368 22336 96688 22337
rect 96368 22272 96376 22336
rect 96440 22272 96456 22336
rect 96520 22272 96536 22336
rect 96600 22272 96616 22336
rect 96680 22272 96688 22336
rect 96368 22271 96688 22272
rect 118049 21858 118115 21861
rect 119200 21858 120000 21888
rect 118049 21856 120000 21858
rect 118049 21800 118054 21856
rect 118110 21800 120000 21856
rect 118049 21798 120000 21800
rect 118049 21795 118115 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 81008 21792 81328 21793
rect 81008 21728 81016 21792
rect 81080 21728 81096 21792
rect 81160 21728 81176 21792
rect 81240 21728 81256 21792
rect 81320 21728 81328 21792
rect 81008 21727 81328 21728
rect 111728 21792 112048 21793
rect 111728 21728 111736 21792
rect 111800 21728 111816 21792
rect 111880 21728 111896 21792
rect 111960 21728 111976 21792
rect 112040 21728 112048 21792
rect 119200 21768 120000 21798
rect 111728 21727 112048 21728
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 65648 21248 65968 21249
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 21183 65968 21184
rect 96368 21248 96688 21249
rect 96368 21184 96376 21248
rect 96440 21184 96456 21248
rect 96520 21184 96536 21248
rect 96600 21184 96616 21248
rect 96680 21184 96688 21248
rect 96368 21183 96688 21184
rect 118049 20906 118115 20909
rect 119200 20906 120000 20936
rect 118049 20904 120000 20906
rect 118049 20848 118054 20904
rect 118110 20848 120000 20904
rect 118049 20846 120000 20848
rect 118049 20843 118115 20846
rect 119200 20816 120000 20846
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 81008 20704 81328 20705
rect 81008 20640 81016 20704
rect 81080 20640 81096 20704
rect 81160 20640 81176 20704
rect 81240 20640 81256 20704
rect 81320 20640 81328 20704
rect 81008 20639 81328 20640
rect 111728 20704 112048 20705
rect 111728 20640 111736 20704
rect 111800 20640 111816 20704
rect 111880 20640 111896 20704
rect 111960 20640 111976 20704
rect 112040 20640 112048 20704
rect 111728 20639 112048 20640
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 65648 20160 65968 20161
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 20095 65968 20096
rect 96368 20160 96688 20161
rect 96368 20096 96376 20160
rect 96440 20096 96456 20160
rect 96520 20096 96536 20160
rect 96600 20096 96616 20160
rect 96680 20096 96688 20160
rect 96368 20095 96688 20096
rect 118049 19954 118115 19957
rect 119200 19954 120000 19984
rect 118049 19952 120000 19954
rect 118049 19896 118054 19952
rect 118110 19896 120000 19952
rect 118049 19894 120000 19896
rect 118049 19891 118115 19894
rect 119200 19864 120000 19894
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 81008 19616 81328 19617
rect 81008 19552 81016 19616
rect 81080 19552 81096 19616
rect 81160 19552 81176 19616
rect 81240 19552 81256 19616
rect 81320 19552 81328 19616
rect 81008 19551 81328 19552
rect 111728 19616 112048 19617
rect 111728 19552 111736 19616
rect 111800 19552 111816 19616
rect 111880 19552 111896 19616
rect 111960 19552 111976 19616
rect 112040 19552 112048 19616
rect 111728 19551 112048 19552
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 65648 19072 65968 19073
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 19007 65968 19008
rect 96368 19072 96688 19073
rect 96368 19008 96376 19072
rect 96440 19008 96456 19072
rect 96520 19008 96536 19072
rect 96600 19008 96616 19072
rect 96680 19008 96688 19072
rect 96368 19007 96688 19008
rect 118049 19002 118115 19005
rect 119200 19002 120000 19032
rect 118049 19000 120000 19002
rect 118049 18944 118054 19000
rect 118110 18944 120000 19000
rect 118049 18942 120000 18944
rect 118049 18939 118115 18942
rect 119200 18912 120000 18942
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 81008 18528 81328 18529
rect 81008 18464 81016 18528
rect 81080 18464 81096 18528
rect 81160 18464 81176 18528
rect 81240 18464 81256 18528
rect 81320 18464 81328 18528
rect 81008 18463 81328 18464
rect 111728 18528 112048 18529
rect 111728 18464 111736 18528
rect 111800 18464 111816 18528
rect 111880 18464 111896 18528
rect 111960 18464 111976 18528
rect 112040 18464 112048 18528
rect 111728 18463 112048 18464
rect 118049 18050 118115 18053
rect 119200 18050 120000 18080
rect 118049 18048 120000 18050
rect 118049 17992 118054 18048
rect 118110 17992 120000 18048
rect 118049 17990 120000 17992
rect 118049 17987 118115 17990
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 65648 17984 65968 17985
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 17919 65968 17920
rect 96368 17984 96688 17985
rect 96368 17920 96376 17984
rect 96440 17920 96456 17984
rect 96520 17920 96536 17984
rect 96600 17920 96616 17984
rect 96680 17920 96688 17984
rect 119200 17960 120000 17990
rect 96368 17919 96688 17920
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 81008 17440 81328 17441
rect 81008 17376 81016 17440
rect 81080 17376 81096 17440
rect 81160 17376 81176 17440
rect 81240 17376 81256 17440
rect 81320 17376 81328 17440
rect 81008 17375 81328 17376
rect 111728 17440 112048 17441
rect 111728 17376 111736 17440
rect 111800 17376 111816 17440
rect 111880 17376 111896 17440
rect 111960 17376 111976 17440
rect 112040 17376 112048 17440
rect 111728 17375 112048 17376
rect 118049 17234 118115 17237
rect 119200 17234 120000 17264
rect 118049 17232 120000 17234
rect 118049 17176 118054 17232
rect 118110 17176 120000 17232
rect 118049 17174 120000 17176
rect 118049 17171 118115 17174
rect 119200 17144 120000 17174
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 65648 16896 65968 16897
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 16831 65968 16832
rect 96368 16896 96688 16897
rect 96368 16832 96376 16896
rect 96440 16832 96456 16896
rect 96520 16832 96536 16896
rect 96600 16832 96616 16896
rect 96680 16832 96688 16896
rect 96368 16831 96688 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 16287 50608 16288
rect 81008 16352 81328 16353
rect 81008 16288 81016 16352
rect 81080 16288 81096 16352
rect 81160 16288 81176 16352
rect 81240 16288 81256 16352
rect 81320 16288 81328 16352
rect 81008 16287 81328 16288
rect 111728 16352 112048 16353
rect 111728 16288 111736 16352
rect 111800 16288 111816 16352
rect 111880 16288 111896 16352
rect 111960 16288 111976 16352
rect 112040 16288 112048 16352
rect 111728 16287 112048 16288
rect 118049 16282 118115 16285
rect 119200 16282 120000 16312
rect 118049 16280 120000 16282
rect 118049 16224 118054 16280
rect 118110 16224 120000 16280
rect 118049 16222 120000 16224
rect 118049 16219 118115 16222
rect 119200 16192 120000 16222
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 65648 15808 65968 15809
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 15743 65968 15744
rect 96368 15808 96688 15809
rect 96368 15744 96376 15808
rect 96440 15744 96456 15808
rect 96520 15744 96536 15808
rect 96600 15744 96616 15808
rect 96680 15744 96688 15808
rect 96368 15743 96688 15744
rect 118049 15330 118115 15333
rect 119200 15330 120000 15360
rect 118049 15328 120000 15330
rect 118049 15272 118054 15328
rect 118110 15272 120000 15328
rect 118049 15270 120000 15272
rect 118049 15267 118115 15270
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 81008 15264 81328 15265
rect 81008 15200 81016 15264
rect 81080 15200 81096 15264
rect 81160 15200 81176 15264
rect 81240 15200 81256 15264
rect 81320 15200 81328 15264
rect 81008 15199 81328 15200
rect 111728 15264 112048 15265
rect 111728 15200 111736 15264
rect 111800 15200 111816 15264
rect 111880 15200 111896 15264
rect 111960 15200 111976 15264
rect 112040 15200 112048 15264
rect 119200 15240 120000 15270
rect 111728 15199 112048 15200
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 65648 14720 65968 14721
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 14655 65968 14656
rect 96368 14720 96688 14721
rect 96368 14656 96376 14720
rect 96440 14656 96456 14720
rect 96520 14656 96536 14720
rect 96600 14656 96616 14720
rect 96680 14656 96688 14720
rect 96368 14655 96688 14656
rect 118049 14378 118115 14381
rect 119200 14378 120000 14408
rect 118049 14376 120000 14378
rect 118049 14320 118054 14376
rect 118110 14320 120000 14376
rect 118049 14318 120000 14320
rect 118049 14315 118115 14318
rect 119200 14288 120000 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 81008 14176 81328 14177
rect 81008 14112 81016 14176
rect 81080 14112 81096 14176
rect 81160 14112 81176 14176
rect 81240 14112 81256 14176
rect 81320 14112 81328 14176
rect 81008 14111 81328 14112
rect 111728 14176 112048 14177
rect 111728 14112 111736 14176
rect 111800 14112 111816 14176
rect 111880 14112 111896 14176
rect 111960 14112 111976 14176
rect 112040 14112 112048 14176
rect 111728 14111 112048 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 65648 13632 65968 13633
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 13567 65968 13568
rect 96368 13632 96688 13633
rect 96368 13568 96376 13632
rect 96440 13568 96456 13632
rect 96520 13568 96536 13632
rect 96600 13568 96616 13632
rect 96680 13568 96688 13632
rect 96368 13567 96688 13568
rect 118049 13426 118115 13429
rect 119200 13426 120000 13456
rect 118049 13424 120000 13426
rect 118049 13368 118054 13424
rect 118110 13368 120000 13424
rect 118049 13366 120000 13368
rect 118049 13363 118115 13366
rect 119200 13336 120000 13366
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 81008 13088 81328 13089
rect 81008 13024 81016 13088
rect 81080 13024 81096 13088
rect 81160 13024 81176 13088
rect 81240 13024 81256 13088
rect 81320 13024 81328 13088
rect 81008 13023 81328 13024
rect 111728 13088 112048 13089
rect 111728 13024 111736 13088
rect 111800 13024 111816 13088
rect 111880 13024 111896 13088
rect 111960 13024 111976 13088
rect 112040 13024 112048 13088
rect 111728 13023 112048 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 65648 12544 65968 12545
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 12479 65968 12480
rect 96368 12544 96688 12545
rect 96368 12480 96376 12544
rect 96440 12480 96456 12544
rect 96520 12480 96536 12544
rect 96600 12480 96616 12544
rect 96680 12480 96688 12544
rect 96368 12479 96688 12480
rect 118049 12474 118115 12477
rect 119200 12474 120000 12504
rect 118049 12472 120000 12474
rect 118049 12416 118054 12472
rect 118110 12416 120000 12472
rect 118049 12414 120000 12416
rect 118049 12411 118115 12414
rect 119200 12384 120000 12414
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 81008 12000 81328 12001
rect 81008 11936 81016 12000
rect 81080 11936 81096 12000
rect 81160 11936 81176 12000
rect 81240 11936 81256 12000
rect 81320 11936 81328 12000
rect 81008 11935 81328 11936
rect 111728 12000 112048 12001
rect 111728 11936 111736 12000
rect 111800 11936 111816 12000
rect 111880 11936 111896 12000
rect 111960 11936 111976 12000
rect 112040 11936 112048 12000
rect 111728 11935 112048 11936
rect 118049 11658 118115 11661
rect 119200 11658 120000 11688
rect 118049 11656 120000 11658
rect 118049 11600 118054 11656
rect 118110 11600 120000 11656
rect 118049 11598 120000 11600
rect 118049 11595 118115 11598
rect 119200 11568 120000 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 65648 11456 65968 11457
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 11391 65968 11392
rect 96368 11456 96688 11457
rect 96368 11392 96376 11456
rect 96440 11392 96456 11456
rect 96520 11392 96536 11456
rect 96600 11392 96616 11456
rect 96680 11392 96688 11456
rect 96368 11391 96688 11392
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 81008 10912 81328 10913
rect 81008 10848 81016 10912
rect 81080 10848 81096 10912
rect 81160 10848 81176 10912
rect 81240 10848 81256 10912
rect 81320 10848 81328 10912
rect 81008 10847 81328 10848
rect 111728 10912 112048 10913
rect 111728 10848 111736 10912
rect 111800 10848 111816 10912
rect 111880 10848 111896 10912
rect 111960 10848 111976 10912
rect 112040 10848 112048 10912
rect 111728 10847 112048 10848
rect 118049 10706 118115 10709
rect 119200 10706 120000 10736
rect 118049 10704 120000 10706
rect 118049 10648 118054 10704
rect 118110 10648 120000 10704
rect 118049 10646 120000 10648
rect 118049 10643 118115 10646
rect 119200 10616 120000 10646
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 65648 10368 65968 10369
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 10303 65968 10304
rect 96368 10368 96688 10369
rect 96368 10304 96376 10368
rect 96440 10304 96456 10368
rect 96520 10304 96536 10368
rect 96600 10304 96616 10368
rect 96680 10304 96688 10368
rect 96368 10303 96688 10304
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 81008 9824 81328 9825
rect 81008 9760 81016 9824
rect 81080 9760 81096 9824
rect 81160 9760 81176 9824
rect 81240 9760 81256 9824
rect 81320 9760 81328 9824
rect 81008 9759 81328 9760
rect 111728 9824 112048 9825
rect 111728 9760 111736 9824
rect 111800 9760 111816 9824
rect 111880 9760 111896 9824
rect 111960 9760 111976 9824
rect 112040 9760 112048 9824
rect 111728 9759 112048 9760
rect 117773 9754 117839 9757
rect 119200 9754 120000 9784
rect 117773 9752 120000 9754
rect 117773 9696 117778 9752
rect 117834 9696 120000 9752
rect 117773 9694 120000 9696
rect 117773 9691 117839 9694
rect 119200 9664 120000 9694
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 65648 9280 65968 9281
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 9215 65968 9216
rect 96368 9280 96688 9281
rect 96368 9216 96376 9280
rect 96440 9216 96456 9280
rect 96520 9216 96536 9280
rect 96600 9216 96616 9280
rect 96680 9216 96688 9280
rect 96368 9215 96688 9216
rect 117773 8802 117839 8805
rect 119200 8802 120000 8832
rect 117773 8800 120000 8802
rect 117773 8744 117778 8800
rect 117834 8744 120000 8800
rect 117773 8742 120000 8744
rect 117773 8739 117839 8742
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 81008 8736 81328 8737
rect 81008 8672 81016 8736
rect 81080 8672 81096 8736
rect 81160 8672 81176 8736
rect 81240 8672 81256 8736
rect 81320 8672 81328 8736
rect 81008 8671 81328 8672
rect 111728 8736 112048 8737
rect 111728 8672 111736 8736
rect 111800 8672 111816 8736
rect 111880 8672 111896 8736
rect 111960 8672 111976 8736
rect 112040 8672 112048 8736
rect 119200 8712 120000 8742
rect 111728 8671 112048 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 65648 8192 65968 8193
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 8127 65968 8128
rect 96368 8192 96688 8193
rect 96368 8128 96376 8192
rect 96440 8128 96456 8192
rect 96520 8128 96536 8192
rect 96600 8128 96616 8192
rect 96680 8128 96688 8192
rect 96368 8127 96688 8128
rect 117773 7850 117839 7853
rect 119200 7850 120000 7880
rect 117773 7848 120000 7850
rect 117773 7792 117778 7848
rect 117834 7792 120000 7848
rect 117773 7790 120000 7792
rect 117773 7787 117839 7790
rect 119200 7760 120000 7790
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 81008 7648 81328 7649
rect 81008 7584 81016 7648
rect 81080 7584 81096 7648
rect 81160 7584 81176 7648
rect 81240 7584 81256 7648
rect 81320 7584 81328 7648
rect 81008 7583 81328 7584
rect 111728 7648 112048 7649
rect 111728 7584 111736 7648
rect 111800 7584 111816 7648
rect 111880 7584 111896 7648
rect 111960 7584 111976 7648
rect 112040 7584 112048 7648
rect 111728 7583 112048 7584
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 65648 7104 65968 7105
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 7039 65968 7040
rect 96368 7104 96688 7105
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 7039 96688 7040
rect 117773 6898 117839 6901
rect 119200 6898 120000 6928
rect 117773 6896 120000 6898
rect 117773 6840 117778 6896
rect 117834 6840 120000 6896
rect 117773 6838 120000 6840
rect 117773 6835 117839 6838
rect 119200 6808 120000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 81008 6560 81328 6561
rect 81008 6496 81016 6560
rect 81080 6496 81096 6560
rect 81160 6496 81176 6560
rect 81240 6496 81256 6560
rect 81320 6496 81328 6560
rect 81008 6495 81328 6496
rect 111728 6560 112048 6561
rect 111728 6496 111736 6560
rect 111800 6496 111816 6560
rect 111880 6496 111896 6560
rect 111960 6496 111976 6560
rect 112040 6496 112048 6560
rect 111728 6495 112048 6496
rect 117773 6082 117839 6085
rect 119200 6082 120000 6112
rect 117773 6080 120000 6082
rect 117773 6024 117778 6080
rect 117834 6024 120000 6080
rect 117773 6022 120000 6024
rect 117773 6019 117839 6022
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 65648 6016 65968 6017
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 5951 65968 5952
rect 96368 6016 96688 6017
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 119200 5992 120000 6022
rect 96368 5951 96688 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 81008 5472 81328 5473
rect 81008 5408 81016 5472
rect 81080 5408 81096 5472
rect 81160 5408 81176 5472
rect 81240 5408 81256 5472
rect 81320 5408 81328 5472
rect 81008 5407 81328 5408
rect 111728 5472 112048 5473
rect 111728 5408 111736 5472
rect 111800 5408 111816 5472
rect 111880 5408 111896 5472
rect 111960 5408 111976 5472
rect 112040 5408 112048 5472
rect 111728 5407 112048 5408
rect 117773 5130 117839 5133
rect 119200 5130 120000 5160
rect 117773 5128 120000 5130
rect 117773 5072 117778 5128
rect 117834 5072 120000 5128
rect 117773 5070 120000 5072
rect 117773 5067 117839 5070
rect 119200 5040 120000 5070
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 65648 4928 65968 4929
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 4863 65968 4864
rect 96368 4928 96688 4929
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 4863 96688 4864
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 81008 4384 81328 4385
rect 81008 4320 81016 4384
rect 81080 4320 81096 4384
rect 81160 4320 81176 4384
rect 81240 4320 81256 4384
rect 81320 4320 81328 4384
rect 81008 4319 81328 4320
rect 111728 4384 112048 4385
rect 111728 4320 111736 4384
rect 111800 4320 111816 4384
rect 111880 4320 111896 4384
rect 111960 4320 111976 4384
rect 112040 4320 112048 4384
rect 111728 4319 112048 4320
rect 117773 4178 117839 4181
rect 119200 4178 120000 4208
rect 117773 4176 120000 4178
rect 117773 4120 117778 4176
rect 117834 4120 120000 4176
rect 117773 4118 120000 4120
rect 117773 4115 117839 4118
rect 119200 4088 120000 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 65648 3840 65968 3841
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 3775 65968 3776
rect 96368 3840 96688 3841
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 3775 96688 3776
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 81008 3296 81328 3297
rect 81008 3232 81016 3296
rect 81080 3232 81096 3296
rect 81160 3232 81176 3296
rect 81240 3232 81256 3296
rect 81320 3232 81328 3296
rect 81008 3231 81328 3232
rect 111728 3296 112048 3297
rect 111728 3232 111736 3296
rect 111800 3232 111816 3296
rect 111880 3232 111896 3296
rect 111960 3232 111976 3296
rect 112040 3232 112048 3296
rect 111728 3231 112048 3232
rect 99649 3226 99715 3229
rect 100569 3226 100635 3229
rect 99649 3224 100635 3226
rect 99649 3168 99654 3224
rect 99710 3168 100574 3224
rect 100630 3168 100635 3224
rect 99649 3166 100635 3168
rect 99649 3163 99715 3166
rect 100569 3163 100635 3166
rect 117221 3226 117287 3229
rect 119200 3226 120000 3256
rect 117221 3224 120000 3226
rect 117221 3168 117226 3224
rect 117282 3168 120000 3224
rect 117221 3166 120000 3168
rect 117221 3163 117287 3166
rect 119200 3136 120000 3166
rect 97625 3090 97691 3093
rect 100753 3090 100819 3093
rect 97625 3088 100819 3090
rect 97625 3032 97630 3088
rect 97686 3032 100758 3088
rect 100814 3032 100819 3088
rect 97625 3030 100819 3032
rect 97625 3027 97691 3030
rect 100753 3027 100819 3030
rect 65241 2954 65307 2957
rect 57930 2952 65307 2954
rect 57930 2896 65246 2952
rect 65302 2896 65307 2952
rect 57930 2894 65307 2896
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 56685 2682 56751 2685
rect 57930 2682 57990 2894
rect 65241 2891 65307 2894
rect 59813 2818 59879 2821
rect 65149 2818 65215 2821
rect 59813 2816 65215 2818
rect 59813 2760 59818 2816
rect 59874 2760 65154 2816
rect 65210 2760 65215 2816
rect 59813 2758 65215 2760
rect 59813 2755 59879 2758
rect 65149 2755 65215 2758
rect 65648 2752 65968 2753
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2687 65968 2688
rect 96368 2752 96688 2753
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 2687 96688 2688
rect 61285 2682 61351 2685
rect 56685 2680 57990 2682
rect 56685 2624 56690 2680
rect 56746 2624 57990 2680
rect 56685 2622 57990 2624
rect 59862 2680 61351 2682
rect 59862 2624 61290 2680
rect 61346 2624 61351 2680
rect 59862 2622 61351 2624
rect 56685 2619 56751 2622
rect 35893 2546 35959 2549
rect 45461 2546 45527 2549
rect 35893 2544 45527 2546
rect 35893 2488 35898 2544
rect 35954 2488 45466 2544
rect 45522 2488 45527 2544
rect 35893 2486 45527 2488
rect 35893 2483 35959 2486
rect 45461 2483 45527 2486
rect 55765 2546 55831 2549
rect 58433 2546 58499 2549
rect 59862 2546 59922 2622
rect 61285 2619 61351 2622
rect 98453 2682 98519 2685
rect 99557 2682 99623 2685
rect 98453 2680 99623 2682
rect 98453 2624 98458 2680
rect 98514 2624 99562 2680
rect 99618 2624 99623 2680
rect 98453 2622 99623 2624
rect 98453 2619 98519 2622
rect 99557 2619 99623 2622
rect 55765 2544 58499 2546
rect 55765 2488 55770 2544
rect 55826 2488 58438 2544
rect 58494 2488 58499 2544
rect 55765 2486 58499 2488
rect 55765 2483 55831 2486
rect 58433 2483 58499 2486
rect 58574 2486 59922 2546
rect 60273 2546 60339 2549
rect 64137 2546 64203 2549
rect 60273 2544 64203 2546
rect 60273 2488 60278 2544
rect 60334 2488 64142 2544
rect 64198 2488 64203 2544
rect 60273 2486 64203 2488
rect 35709 2410 35775 2413
rect 35985 2410 36051 2413
rect 35709 2408 36051 2410
rect 35709 2352 35714 2408
rect 35770 2352 35990 2408
rect 36046 2352 36051 2408
rect 35709 2350 36051 2352
rect 35709 2347 35775 2350
rect 35985 2347 36051 2350
rect 45369 2410 45435 2413
rect 45737 2410 45803 2413
rect 45369 2408 45803 2410
rect 45369 2352 45374 2408
rect 45430 2352 45742 2408
rect 45798 2352 45803 2408
rect 45369 2350 45803 2352
rect 45369 2347 45435 2350
rect 45737 2347 45803 2350
rect 49049 2410 49115 2413
rect 53373 2410 53439 2413
rect 58574 2410 58634 2486
rect 60273 2483 60339 2486
rect 64137 2483 64203 2486
rect 98729 2546 98795 2549
rect 105445 2546 105511 2549
rect 98729 2544 105511 2546
rect 98729 2488 98734 2544
rect 98790 2488 105450 2544
rect 105506 2488 105511 2544
rect 98729 2486 105511 2488
rect 98729 2483 98795 2486
rect 105445 2483 105511 2486
rect 49049 2408 51090 2410
rect 49049 2352 49054 2408
rect 49110 2352 51090 2408
rect 49049 2350 51090 2352
rect 49049 2347 49115 2350
rect 37273 2274 37339 2277
rect 45369 2274 45435 2277
rect 37273 2272 45435 2274
rect 37273 2216 37278 2272
rect 37334 2216 45374 2272
rect 45430 2216 45435 2272
rect 37273 2214 45435 2216
rect 37273 2211 37339 2214
rect 45369 2211 45435 2214
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 51030 2138 51090 2350
rect 53373 2408 58634 2410
rect 53373 2352 53378 2408
rect 53434 2352 58634 2408
rect 53373 2350 58634 2352
rect 59629 2410 59695 2413
rect 66897 2410 66963 2413
rect 59629 2408 66963 2410
rect 59629 2352 59634 2408
rect 59690 2352 66902 2408
rect 66958 2352 66963 2408
rect 59629 2350 66963 2352
rect 53373 2347 53439 2350
rect 59629 2347 59695 2350
rect 66897 2347 66963 2350
rect 74809 2410 74875 2413
rect 81433 2410 81499 2413
rect 74809 2408 81499 2410
rect 74809 2352 74814 2408
rect 74870 2352 81438 2408
rect 81494 2352 81499 2408
rect 74809 2350 81499 2352
rect 74809 2347 74875 2350
rect 81433 2347 81499 2350
rect 97533 2410 97599 2413
rect 105721 2410 105787 2413
rect 97533 2408 105787 2410
rect 97533 2352 97538 2408
rect 97594 2352 105726 2408
rect 105782 2352 105787 2408
rect 97533 2350 105787 2352
rect 97533 2347 97599 2350
rect 105721 2347 105787 2350
rect 55673 2274 55739 2277
rect 59721 2274 59787 2277
rect 55673 2272 59787 2274
rect 55673 2216 55678 2272
rect 55734 2216 59726 2272
rect 59782 2216 59787 2272
rect 55673 2214 59787 2216
rect 55673 2211 55739 2214
rect 59721 2211 59787 2214
rect 60181 2274 60247 2277
rect 60590 2274 60596 2276
rect 60181 2272 60596 2274
rect 60181 2216 60186 2272
rect 60242 2216 60596 2272
rect 60181 2214 60596 2216
rect 60181 2211 60247 2214
rect 60590 2212 60596 2214
rect 60660 2212 60666 2276
rect 60733 2274 60799 2277
rect 67449 2274 67515 2277
rect 60733 2272 67515 2274
rect 60733 2216 60738 2272
rect 60794 2216 67454 2272
rect 67510 2216 67515 2272
rect 60733 2214 67515 2216
rect 60733 2211 60799 2214
rect 67449 2211 67515 2214
rect 74441 2274 74507 2277
rect 79501 2274 79567 2277
rect 74441 2272 79567 2274
rect 74441 2216 74446 2272
rect 74502 2216 79506 2272
rect 79562 2216 79567 2272
rect 74441 2214 79567 2216
rect 74441 2211 74507 2214
rect 79501 2211 79567 2214
rect 117129 2274 117195 2277
rect 119200 2274 120000 2304
rect 117129 2272 120000 2274
rect 117129 2216 117134 2272
rect 117190 2216 120000 2272
rect 117129 2214 120000 2216
rect 117129 2211 117195 2214
rect 81008 2208 81328 2209
rect 81008 2144 81016 2208
rect 81080 2144 81096 2208
rect 81160 2144 81176 2208
rect 81240 2144 81256 2208
rect 81320 2144 81328 2208
rect 81008 2143 81328 2144
rect 111728 2208 112048 2209
rect 111728 2144 111736 2208
rect 111800 2144 111816 2208
rect 111880 2144 111896 2208
rect 111960 2144 111976 2208
rect 112040 2144 112048 2208
rect 119200 2184 120000 2214
rect 111728 2143 112048 2144
rect 69657 2138 69723 2141
rect 51030 2136 69723 2138
rect 51030 2080 69662 2136
rect 69718 2080 69723 2136
rect 51030 2078 69723 2080
rect 69657 2075 69723 2078
rect 51073 2002 51139 2005
rect 59905 2002 59971 2005
rect 60365 2002 60431 2005
rect 51073 2000 59971 2002
rect 51073 1944 51078 2000
rect 51134 1944 59910 2000
rect 59966 1944 59971 2000
rect 51073 1942 59971 1944
rect 51073 1939 51139 1942
rect 59905 1939 59971 1942
rect 60046 2000 60431 2002
rect 60046 1944 60370 2000
rect 60426 1944 60431 2000
rect 60046 1942 60431 1944
rect 33409 1866 33475 1869
rect 35801 1866 35867 1869
rect 33409 1864 35867 1866
rect 33409 1808 33414 1864
rect 33470 1808 35806 1864
rect 35862 1808 35867 1864
rect 33409 1806 35867 1808
rect 33409 1803 33475 1806
rect 35801 1803 35867 1806
rect 51073 1866 51139 1869
rect 60046 1866 60106 1942
rect 60365 1939 60431 1942
rect 60590 1940 60596 2004
rect 60660 2002 60666 2004
rect 70301 2002 70367 2005
rect 60660 2000 70367 2002
rect 60660 1944 70306 2000
rect 70362 1944 70367 2000
rect 60660 1942 70367 1944
rect 60660 1940 60666 1942
rect 70301 1939 70367 1942
rect 51073 1864 60106 1866
rect 51073 1808 51078 1864
rect 51134 1808 60106 1864
rect 51073 1806 60106 1808
rect 60181 1866 60247 1869
rect 63401 1866 63467 1869
rect 60181 1864 63467 1866
rect 60181 1808 60186 1864
rect 60242 1808 63406 1864
rect 63462 1808 63467 1864
rect 60181 1806 63467 1808
rect 51073 1803 51139 1806
rect 60181 1803 60247 1806
rect 63401 1803 63467 1806
rect 40493 1730 40559 1733
rect 45645 1730 45711 1733
rect 40493 1728 45711 1730
rect 40493 1672 40498 1728
rect 40554 1672 45650 1728
rect 45706 1672 45711 1728
rect 40493 1670 45711 1672
rect 40493 1667 40559 1670
rect 45645 1667 45711 1670
rect 51165 1730 51231 1733
rect 60549 1730 60615 1733
rect 51165 1728 60615 1730
rect 51165 1672 51170 1728
rect 51226 1672 60554 1728
rect 60610 1672 60615 1728
rect 51165 1670 60615 1672
rect 51165 1667 51231 1670
rect 60549 1667 60615 1670
rect 70209 1730 70275 1733
rect 73981 1730 74047 1733
rect 70209 1728 74047 1730
rect 70209 1672 70214 1728
rect 70270 1672 73986 1728
rect 74042 1672 74047 1728
rect 70209 1670 74047 1672
rect 70209 1667 70275 1670
rect 73981 1667 74047 1670
rect 47669 1594 47735 1597
rect 51257 1594 51323 1597
rect 47669 1592 51323 1594
rect 47669 1536 47674 1592
rect 47730 1536 51262 1592
rect 51318 1536 51323 1592
rect 47669 1534 51323 1536
rect 47669 1531 47735 1534
rect 51257 1531 51323 1534
rect 60733 1458 60799 1461
rect 69749 1458 69815 1461
rect 60733 1456 69815 1458
rect 60733 1400 60738 1456
rect 60794 1400 69754 1456
rect 69810 1400 69815 1456
rect 60733 1398 69815 1400
rect 60733 1395 60799 1398
rect 69749 1395 69815 1398
rect 76005 1458 76071 1461
rect 77661 1458 77727 1461
rect 76005 1456 77727 1458
rect 76005 1400 76010 1456
rect 76066 1400 77666 1456
rect 77722 1400 77727 1456
rect 76005 1398 77727 1400
rect 76005 1395 76071 1398
rect 77661 1395 77727 1398
rect 60457 1322 60523 1325
rect 61193 1322 61259 1325
rect 60457 1320 61259 1322
rect 60457 1264 60462 1320
rect 60518 1264 61198 1320
rect 61254 1264 61259 1320
rect 60457 1262 61259 1264
rect 60457 1259 60523 1262
rect 61193 1259 61259 1262
rect 117773 1322 117839 1325
rect 119200 1322 120000 1352
rect 117773 1320 120000 1322
rect 117773 1264 117778 1320
rect 117834 1264 120000 1320
rect 117773 1262 120000 1264
rect 117773 1259 117839 1262
rect 119200 1232 120000 1262
rect 116485 506 116551 509
rect 119200 506 120000 536
rect 116485 504 120000 506
rect 116485 448 116490 504
rect 116546 448 120000 504
rect 116485 446 120000 448
rect 116485 443 116551 446
rect 119200 416 120000 446
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 96376 37564 96440 37568
rect 96376 37508 96380 37564
rect 96380 37508 96436 37564
rect 96436 37508 96440 37564
rect 96376 37504 96440 37508
rect 96456 37564 96520 37568
rect 96456 37508 96460 37564
rect 96460 37508 96516 37564
rect 96516 37508 96520 37564
rect 96456 37504 96520 37508
rect 96536 37564 96600 37568
rect 96536 37508 96540 37564
rect 96540 37508 96596 37564
rect 96596 37508 96600 37564
rect 96536 37504 96600 37508
rect 96616 37564 96680 37568
rect 96616 37508 96620 37564
rect 96620 37508 96676 37564
rect 96676 37508 96680 37564
rect 96616 37504 96680 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 81016 37020 81080 37024
rect 81016 36964 81020 37020
rect 81020 36964 81076 37020
rect 81076 36964 81080 37020
rect 81016 36960 81080 36964
rect 81096 37020 81160 37024
rect 81096 36964 81100 37020
rect 81100 36964 81156 37020
rect 81156 36964 81160 37020
rect 81096 36960 81160 36964
rect 81176 37020 81240 37024
rect 81176 36964 81180 37020
rect 81180 36964 81236 37020
rect 81236 36964 81240 37020
rect 81176 36960 81240 36964
rect 81256 37020 81320 37024
rect 81256 36964 81260 37020
rect 81260 36964 81316 37020
rect 81316 36964 81320 37020
rect 81256 36960 81320 36964
rect 111736 37020 111800 37024
rect 111736 36964 111740 37020
rect 111740 36964 111796 37020
rect 111796 36964 111800 37020
rect 111736 36960 111800 36964
rect 111816 37020 111880 37024
rect 111816 36964 111820 37020
rect 111820 36964 111876 37020
rect 111876 36964 111880 37020
rect 111816 36960 111880 36964
rect 111896 37020 111960 37024
rect 111896 36964 111900 37020
rect 111900 36964 111956 37020
rect 111956 36964 111960 37020
rect 111896 36960 111960 36964
rect 111976 37020 112040 37024
rect 111976 36964 111980 37020
rect 111980 36964 112036 37020
rect 112036 36964 112040 37020
rect 111976 36960 112040 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 96376 36476 96440 36480
rect 96376 36420 96380 36476
rect 96380 36420 96436 36476
rect 96436 36420 96440 36476
rect 96376 36416 96440 36420
rect 96456 36476 96520 36480
rect 96456 36420 96460 36476
rect 96460 36420 96516 36476
rect 96516 36420 96520 36476
rect 96456 36416 96520 36420
rect 96536 36476 96600 36480
rect 96536 36420 96540 36476
rect 96540 36420 96596 36476
rect 96596 36420 96600 36476
rect 96536 36416 96600 36420
rect 96616 36476 96680 36480
rect 96616 36420 96620 36476
rect 96620 36420 96676 36476
rect 96676 36420 96680 36476
rect 96616 36416 96680 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 81016 35932 81080 35936
rect 81016 35876 81020 35932
rect 81020 35876 81076 35932
rect 81076 35876 81080 35932
rect 81016 35872 81080 35876
rect 81096 35932 81160 35936
rect 81096 35876 81100 35932
rect 81100 35876 81156 35932
rect 81156 35876 81160 35932
rect 81096 35872 81160 35876
rect 81176 35932 81240 35936
rect 81176 35876 81180 35932
rect 81180 35876 81236 35932
rect 81236 35876 81240 35932
rect 81176 35872 81240 35876
rect 81256 35932 81320 35936
rect 81256 35876 81260 35932
rect 81260 35876 81316 35932
rect 81316 35876 81320 35932
rect 81256 35872 81320 35876
rect 111736 35932 111800 35936
rect 111736 35876 111740 35932
rect 111740 35876 111796 35932
rect 111796 35876 111800 35932
rect 111736 35872 111800 35876
rect 111816 35932 111880 35936
rect 111816 35876 111820 35932
rect 111820 35876 111876 35932
rect 111876 35876 111880 35932
rect 111816 35872 111880 35876
rect 111896 35932 111960 35936
rect 111896 35876 111900 35932
rect 111900 35876 111956 35932
rect 111956 35876 111960 35932
rect 111896 35872 111960 35876
rect 111976 35932 112040 35936
rect 111976 35876 111980 35932
rect 111980 35876 112036 35932
rect 112036 35876 112040 35932
rect 111976 35872 112040 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 96376 35388 96440 35392
rect 96376 35332 96380 35388
rect 96380 35332 96436 35388
rect 96436 35332 96440 35388
rect 96376 35328 96440 35332
rect 96456 35388 96520 35392
rect 96456 35332 96460 35388
rect 96460 35332 96516 35388
rect 96516 35332 96520 35388
rect 96456 35328 96520 35332
rect 96536 35388 96600 35392
rect 96536 35332 96540 35388
rect 96540 35332 96596 35388
rect 96596 35332 96600 35388
rect 96536 35328 96600 35332
rect 96616 35388 96680 35392
rect 96616 35332 96620 35388
rect 96620 35332 96676 35388
rect 96676 35332 96680 35388
rect 96616 35328 96680 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 81016 34844 81080 34848
rect 81016 34788 81020 34844
rect 81020 34788 81076 34844
rect 81076 34788 81080 34844
rect 81016 34784 81080 34788
rect 81096 34844 81160 34848
rect 81096 34788 81100 34844
rect 81100 34788 81156 34844
rect 81156 34788 81160 34844
rect 81096 34784 81160 34788
rect 81176 34844 81240 34848
rect 81176 34788 81180 34844
rect 81180 34788 81236 34844
rect 81236 34788 81240 34844
rect 81176 34784 81240 34788
rect 81256 34844 81320 34848
rect 81256 34788 81260 34844
rect 81260 34788 81316 34844
rect 81316 34788 81320 34844
rect 81256 34784 81320 34788
rect 111736 34844 111800 34848
rect 111736 34788 111740 34844
rect 111740 34788 111796 34844
rect 111796 34788 111800 34844
rect 111736 34784 111800 34788
rect 111816 34844 111880 34848
rect 111816 34788 111820 34844
rect 111820 34788 111876 34844
rect 111876 34788 111880 34844
rect 111816 34784 111880 34788
rect 111896 34844 111960 34848
rect 111896 34788 111900 34844
rect 111900 34788 111956 34844
rect 111956 34788 111960 34844
rect 111896 34784 111960 34788
rect 111976 34844 112040 34848
rect 111976 34788 111980 34844
rect 111980 34788 112036 34844
rect 112036 34788 112040 34844
rect 111976 34784 112040 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 96376 34300 96440 34304
rect 96376 34244 96380 34300
rect 96380 34244 96436 34300
rect 96436 34244 96440 34300
rect 96376 34240 96440 34244
rect 96456 34300 96520 34304
rect 96456 34244 96460 34300
rect 96460 34244 96516 34300
rect 96516 34244 96520 34300
rect 96456 34240 96520 34244
rect 96536 34300 96600 34304
rect 96536 34244 96540 34300
rect 96540 34244 96596 34300
rect 96596 34244 96600 34300
rect 96536 34240 96600 34244
rect 96616 34300 96680 34304
rect 96616 34244 96620 34300
rect 96620 34244 96676 34300
rect 96676 34244 96680 34300
rect 96616 34240 96680 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 81016 33756 81080 33760
rect 81016 33700 81020 33756
rect 81020 33700 81076 33756
rect 81076 33700 81080 33756
rect 81016 33696 81080 33700
rect 81096 33756 81160 33760
rect 81096 33700 81100 33756
rect 81100 33700 81156 33756
rect 81156 33700 81160 33756
rect 81096 33696 81160 33700
rect 81176 33756 81240 33760
rect 81176 33700 81180 33756
rect 81180 33700 81236 33756
rect 81236 33700 81240 33756
rect 81176 33696 81240 33700
rect 81256 33756 81320 33760
rect 81256 33700 81260 33756
rect 81260 33700 81316 33756
rect 81316 33700 81320 33756
rect 81256 33696 81320 33700
rect 111736 33756 111800 33760
rect 111736 33700 111740 33756
rect 111740 33700 111796 33756
rect 111796 33700 111800 33756
rect 111736 33696 111800 33700
rect 111816 33756 111880 33760
rect 111816 33700 111820 33756
rect 111820 33700 111876 33756
rect 111876 33700 111880 33756
rect 111816 33696 111880 33700
rect 111896 33756 111960 33760
rect 111896 33700 111900 33756
rect 111900 33700 111956 33756
rect 111956 33700 111960 33756
rect 111896 33696 111960 33700
rect 111976 33756 112040 33760
rect 111976 33700 111980 33756
rect 111980 33700 112036 33756
rect 112036 33700 112040 33756
rect 111976 33696 112040 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 96376 33212 96440 33216
rect 96376 33156 96380 33212
rect 96380 33156 96436 33212
rect 96436 33156 96440 33212
rect 96376 33152 96440 33156
rect 96456 33212 96520 33216
rect 96456 33156 96460 33212
rect 96460 33156 96516 33212
rect 96516 33156 96520 33212
rect 96456 33152 96520 33156
rect 96536 33212 96600 33216
rect 96536 33156 96540 33212
rect 96540 33156 96596 33212
rect 96596 33156 96600 33212
rect 96536 33152 96600 33156
rect 96616 33212 96680 33216
rect 96616 33156 96620 33212
rect 96620 33156 96676 33212
rect 96676 33156 96680 33212
rect 96616 33152 96680 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 81016 32668 81080 32672
rect 81016 32612 81020 32668
rect 81020 32612 81076 32668
rect 81076 32612 81080 32668
rect 81016 32608 81080 32612
rect 81096 32668 81160 32672
rect 81096 32612 81100 32668
rect 81100 32612 81156 32668
rect 81156 32612 81160 32668
rect 81096 32608 81160 32612
rect 81176 32668 81240 32672
rect 81176 32612 81180 32668
rect 81180 32612 81236 32668
rect 81236 32612 81240 32668
rect 81176 32608 81240 32612
rect 81256 32668 81320 32672
rect 81256 32612 81260 32668
rect 81260 32612 81316 32668
rect 81316 32612 81320 32668
rect 81256 32608 81320 32612
rect 111736 32668 111800 32672
rect 111736 32612 111740 32668
rect 111740 32612 111796 32668
rect 111796 32612 111800 32668
rect 111736 32608 111800 32612
rect 111816 32668 111880 32672
rect 111816 32612 111820 32668
rect 111820 32612 111876 32668
rect 111876 32612 111880 32668
rect 111816 32608 111880 32612
rect 111896 32668 111960 32672
rect 111896 32612 111900 32668
rect 111900 32612 111956 32668
rect 111956 32612 111960 32668
rect 111896 32608 111960 32612
rect 111976 32668 112040 32672
rect 111976 32612 111980 32668
rect 111980 32612 112036 32668
rect 112036 32612 112040 32668
rect 111976 32608 112040 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 96376 32124 96440 32128
rect 96376 32068 96380 32124
rect 96380 32068 96436 32124
rect 96436 32068 96440 32124
rect 96376 32064 96440 32068
rect 96456 32124 96520 32128
rect 96456 32068 96460 32124
rect 96460 32068 96516 32124
rect 96516 32068 96520 32124
rect 96456 32064 96520 32068
rect 96536 32124 96600 32128
rect 96536 32068 96540 32124
rect 96540 32068 96596 32124
rect 96596 32068 96600 32124
rect 96536 32064 96600 32068
rect 96616 32124 96680 32128
rect 96616 32068 96620 32124
rect 96620 32068 96676 32124
rect 96676 32068 96680 32124
rect 96616 32064 96680 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 81016 31580 81080 31584
rect 81016 31524 81020 31580
rect 81020 31524 81076 31580
rect 81076 31524 81080 31580
rect 81016 31520 81080 31524
rect 81096 31580 81160 31584
rect 81096 31524 81100 31580
rect 81100 31524 81156 31580
rect 81156 31524 81160 31580
rect 81096 31520 81160 31524
rect 81176 31580 81240 31584
rect 81176 31524 81180 31580
rect 81180 31524 81236 31580
rect 81236 31524 81240 31580
rect 81176 31520 81240 31524
rect 81256 31580 81320 31584
rect 81256 31524 81260 31580
rect 81260 31524 81316 31580
rect 81316 31524 81320 31580
rect 81256 31520 81320 31524
rect 111736 31580 111800 31584
rect 111736 31524 111740 31580
rect 111740 31524 111796 31580
rect 111796 31524 111800 31580
rect 111736 31520 111800 31524
rect 111816 31580 111880 31584
rect 111816 31524 111820 31580
rect 111820 31524 111876 31580
rect 111876 31524 111880 31580
rect 111816 31520 111880 31524
rect 111896 31580 111960 31584
rect 111896 31524 111900 31580
rect 111900 31524 111956 31580
rect 111956 31524 111960 31580
rect 111896 31520 111960 31524
rect 111976 31580 112040 31584
rect 111976 31524 111980 31580
rect 111980 31524 112036 31580
rect 112036 31524 112040 31580
rect 111976 31520 112040 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 96376 31036 96440 31040
rect 96376 30980 96380 31036
rect 96380 30980 96436 31036
rect 96436 30980 96440 31036
rect 96376 30976 96440 30980
rect 96456 31036 96520 31040
rect 96456 30980 96460 31036
rect 96460 30980 96516 31036
rect 96516 30980 96520 31036
rect 96456 30976 96520 30980
rect 96536 31036 96600 31040
rect 96536 30980 96540 31036
rect 96540 30980 96596 31036
rect 96596 30980 96600 31036
rect 96536 30976 96600 30980
rect 96616 31036 96680 31040
rect 96616 30980 96620 31036
rect 96620 30980 96676 31036
rect 96676 30980 96680 31036
rect 96616 30976 96680 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 81016 30492 81080 30496
rect 81016 30436 81020 30492
rect 81020 30436 81076 30492
rect 81076 30436 81080 30492
rect 81016 30432 81080 30436
rect 81096 30492 81160 30496
rect 81096 30436 81100 30492
rect 81100 30436 81156 30492
rect 81156 30436 81160 30492
rect 81096 30432 81160 30436
rect 81176 30492 81240 30496
rect 81176 30436 81180 30492
rect 81180 30436 81236 30492
rect 81236 30436 81240 30492
rect 81176 30432 81240 30436
rect 81256 30492 81320 30496
rect 81256 30436 81260 30492
rect 81260 30436 81316 30492
rect 81316 30436 81320 30492
rect 81256 30432 81320 30436
rect 111736 30492 111800 30496
rect 111736 30436 111740 30492
rect 111740 30436 111796 30492
rect 111796 30436 111800 30492
rect 111736 30432 111800 30436
rect 111816 30492 111880 30496
rect 111816 30436 111820 30492
rect 111820 30436 111876 30492
rect 111876 30436 111880 30492
rect 111816 30432 111880 30436
rect 111896 30492 111960 30496
rect 111896 30436 111900 30492
rect 111900 30436 111956 30492
rect 111956 30436 111960 30492
rect 111896 30432 111960 30436
rect 111976 30492 112040 30496
rect 111976 30436 111980 30492
rect 111980 30436 112036 30492
rect 112036 30436 112040 30492
rect 111976 30432 112040 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 96376 29948 96440 29952
rect 96376 29892 96380 29948
rect 96380 29892 96436 29948
rect 96436 29892 96440 29948
rect 96376 29888 96440 29892
rect 96456 29948 96520 29952
rect 96456 29892 96460 29948
rect 96460 29892 96516 29948
rect 96516 29892 96520 29948
rect 96456 29888 96520 29892
rect 96536 29948 96600 29952
rect 96536 29892 96540 29948
rect 96540 29892 96596 29948
rect 96596 29892 96600 29948
rect 96536 29888 96600 29892
rect 96616 29948 96680 29952
rect 96616 29892 96620 29948
rect 96620 29892 96676 29948
rect 96676 29892 96680 29948
rect 96616 29888 96680 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 81016 29404 81080 29408
rect 81016 29348 81020 29404
rect 81020 29348 81076 29404
rect 81076 29348 81080 29404
rect 81016 29344 81080 29348
rect 81096 29404 81160 29408
rect 81096 29348 81100 29404
rect 81100 29348 81156 29404
rect 81156 29348 81160 29404
rect 81096 29344 81160 29348
rect 81176 29404 81240 29408
rect 81176 29348 81180 29404
rect 81180 29348 81236 29404
rect 81236 29348 81240 29404
rect 81176 29344 81240 29348
rect 81256 29404 81320 29408
rect 81256 29348 81260 29404
rect 81260 29348 81316 29404
rect 81316 29348 81320 29404
rect 81256 29344 81320 29348
rect 111736 29404 111800 29408
rect 111736 29348 111740 29404
rect 111740 29348 111796 29404
rect 111796 29348 111800 29404
rect 111736 29344 111800 29348
rect 111816 29404 111880 29408
rect 111816 29348 111820 29404
rect 111820 29348 111876 29404
rect 111876 29348 111880 29404
rect 111816 29344 111880 29348
rect 111896 29404 111960 29408
rect 111896 29348 111900 29404
rect 111900 29348 111956 29404
rect 111956 29348 111960 29404
rect 111896 29344 111960 29348
rect 111976 29404 112040 29408
rect 111976 29348 111980 29404
rect 111980 29348 112036 29404
rect 112036 29348 112040 29404
rect 111976 29344 112040 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 96376 28860 96440 28864
rect 96376 28804 96380 28860
rect 96380 28804 96436 28860
rect 96436 28804 96440 28860
rect 96376 28800 96440 28804
rect 96456 28860 96520 28864
rect 96456 28804 96460 28860
rect 96460 28804 96516 28860
rect 96516 28804 96520 28860
rect 96456 28800 96520 28804
rect 96536 28860 96600 28864
rect 96536 28804 96540 28860
rect 96540 28804 96596 28860
rect 96596 28804 96600 28860
rect 96536 28800 96600 28804
rect 96616 28860 96680 28864
rect 96616 28804 96620 28860
rect 96620 28804 96676 28860
rect 96676 28804 96680 28860
rect 96616 28800 96680 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 81016 28316 81080 28320
rect 81016 28260 81020 28316
rect 81020 28260 81076 28316
rect 81076 28260 81080 28316
rect 81016 28256 81080 28260
rect 81096 28316 81160 28320
rect 81096 28260 81100 28316
rect 81100 28260 81156 28316
rect 81156 28260 81160 28316
rect 81096 28256 81160 28260
rect 81176 28316 81240 28320
rect 81176 28260 81180 28316
rect 81180 28260 81236 28316
rect 81236 28260 81240 28316
rect 81176 28256 81240 28260
rect 81256 28316 81320 28320
rect 81256 28260 81260 28316
rect 81260 28260 81316 28316
rect 81316 28260 81320 28316
rect 81256 28256 81320 28260
rect 111736 28316 111800 28320
rect 111736 28260 111740 28316
rect 111740 28260 111796 28316
rect 111796 28260 111800 28316
rect 111736 28256 111800 28260
rect 111816 28316 111880 28320
rect 111816 28260 111820 28316
rect 111820 28260 111876 28316
rect 111876 28260 111880 28316
rect 111816 28256 111880 28260
rect 111896 28316 111960 28320
rect 111896 28260 111900 28316
rect 111900 28260 111956 28316
rect 111956 28260 111960 28316
rect 111896 28256 111960 28260
rect 111976 28316 112040 28320
rect 111976 28260 111980 28316
rect 111980 28260 112036 28316
rect 112036 28260 112040 28316
rect 111976 28256 112040 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 96376 27772 96440 27776
rect 96376 27716 96380 27772
rect 96380 27716 96436 27772
rect 96436 27716 96440 27772
rect 96376 27712 96440 27716
rect 96456 27772 96520 27776
rect 96456 27716 96460 27772
rect 96460 27716 96516 27772
rect 96516 27716 96520 27772
rect 96456 27712 96520 27716
rect 96536 27772 96600 27776
rect 96536 27716 96540 27772
rect 96540 27716 96596 27772
rect 96596 27716 96600 27772
rect 96536 27712 96600 27716
rect 96616 27772 96680 27776
rect 96616 27716 96620 27772
rect 96620 27716 96676 27772
rect 96676 27716 96680 27772
rect 96616 27712 96680 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 81016 27228 81080 27232
rect 81016 27172 81020 27228
rect 81020 27172 81076 27228
rect 81076 27172 81080 27228
rect 81016 27168 81080 27172
rect 81096 27228 81160 27232
rect 81096 27172 81100 27228
rect 81100 27172 81156 27228
rect 81156 27172 81160 27228
rect 81096 27168 81160 27172
rect 81176 27228 81240 27232
rect 81176 27172 81180 27228
rect 81180 27172 81236 27228
rect 81236 27172 81240 27228
rect 81176 27168 81240 27172
rect 81256 27228 81320 27232
rect 81256 27172 81260 27228
rect 81260 27172 81316 27228
rect 81316 27172 81320 27228
rect 81256 27168 81320 27172
rect 111736 27228 111800 27232
rect 111736 27172 111740 27228
rect 111740 27172 111796 27228
rect 111796 27172 111800 27228
rect 111736 27168 111800 27172
rect 111816 27228 111880 27232
rect 111816 27172 111820 27228
rect 111820 27172 111876 27228
rect 111876 27172 111880 27228
rect 111816 27168 111880 27172
rect 111896 27228 111960 27232
rect 111896 27172 111900 27228
rect 111900 27172 111956 27228
rect 111956 27172 111960 27228
rect 111896 27168 111960 27172
rect 111976 27228 112040 27232
rect 111976 27172 111980 27228
rect 111980 27172 112036 27228
rect 112036 27172 112040 27228
rect 111976 27168 112040 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 96376 26684 96440 26688
rect 96376 26628 96380 26684
rect 96380 26628 96436 26684
rect 96436 26628 96440 26684
rect 96376 26624 96440 26628
rect 96456 26684 96520 26688
rect 96456 26628 96460 26684
rect 96460 26628 96516 26684
rect 96516 26628 96520 26684
rect 96456 26624 96520 26628
rect 96536 26684 96600 26688
rect 96536 26628 96540 26684
rect 96540 26628 96596 26684
rect 96596 26628 96600 26684
rect 96536 26624 96600 26628
rect 96616 26684 96680 26688
rect 96616 26628 96620 26684
rect 96620 26628 96676 26684
rect 96676 26628 96680 26684
rect 96616 26624 96680 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 81016 26140 81080 26144
rect 81016 26084 81020 26140
rect 81020 26084 81076 26140
rect 81076 26084 81080 26140
rect 81016 26080 81080 26084
rect 81096 26140 81160 26144
rect 81096 26084 81100 26140
rect 81100 26084 81156 26140
rect 81156 26084 81160 26140
rect 81096 26080 81160 26084
rect 81176 26140 81240 26144
rect 81176 26084 81180 26140
rect 81180 26084 81236 26140
rect 81236 26084 81240 26140
rect 81176 26080 81240 26084
rect 81256 26140 81320 26144
rect 81256 26084 81260 26140
rect 81260 26084 81316 26140
rect 81316 26084 81320 26140
rect 81256 26080 81320 26084
rect 111736 26140 111800 26144
rect 111736 26084 111740 26140
rect 111740 26084 111796 26140
rect 111796 26084 111800 26140
rect 111736 26080 111800 26084
rect 111816 26140 111880 26144
rect 111816 26084 111820 26140
rect 111820 26084 111876 26140
rect 111876 26084 111880 26140
rect 111816 26080 111880 26084
rect 111896 26140 111960 26144
rect 111896 26084 111900 26140
rect 111900 26084 111956 26140
rect 111956 26084 111960 26140
rect 111896 26080 111960 26084
rect 111976 26140 112040 26144
rect 111976 26084 111980 26140
rect 111980 26084 112036 26140
rect 112036 26084 112040 26140
rect 111976 26080 112040 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 96376 25596 96440 25600
rect 96376 25540 96380 25596
rect 96380 25540 96436 25596
rect 96436 25540 96440 25596
rect 96376 25536 96440 25540
rect 96456 25596 96520 25600
rect 96456 25540 96460 25596
rect 96460 25540 96516 25596
rect 96516 25540 96520 25596
rect 96456 25536 96520 25540
rect 96536 25596 96600 25600
rect 96536 25540 96540 25596
rect 96540 25540 96596 25596
rect 96596 25540 96600 25596
rect 96536 25536 96600 25540
rect 96616 25596 96680 25600
rect 96616 25540 96620 25596
rect 96620 25540 96676 25596
rect 96676 25540 96680 25596
rect 96616 25536 96680 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 81016 25052 81080 25056
rect 81016 24996 81020 25052
rect 81020 24996 81076 25052
rect 81076 24996 81080 25052
rect 81016 24992 81080 24996
rect 81096 25052 81160 25056
rect 81096 24996 81100 25052
rect 81100 24996 81156 25052
rect 81156 24996 81160 25052
rect 81096 24992 81160 24996
rect 81176 25052 81240 25056
rect 81176 24996 81180 25052
rect 81180 24996 81236 25052
rect 81236 24996 81240 25052
rect 81176 24992 81240 24996
rect 81256 25052 81320 25056
rect 81256 24996 81260 25052
rect 81260 24996 81316 25052
rect 81316 24996 81320 25052
rect 81256 24992 81320 24996
rect 111736 25052 111800 25056
rect 111736 24996 111740 25052
rect 111740 24996 111796 25052
rect 111796 24996 111800 25052
rect 111736 24992 111800 24996
rect 111816 25052 111880 25056
rect 111816 24996 111820 25052
rect 111820 24996 111876 25052
rect 111876 24996 111880 25052
rect 111816 24992 111880 24996
rect 111896 25052 111960 25056
rect 111896 24996 111900 25052
rect 111900 24996 111956 25052
rect 111956 24996 111960 25052
rect 111896 24992 111960 24996
rect 111976 25052 112040 25056
rect 111976 24996 111980 25052
rect 111980 24996 112036 25052
rect 112036 24996 112040 25052
rect 111976 24992 112040 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 96376 24508 96440 24512
rect 96376 24452 96380 24508
rect 96380 24452 96436 24508
rect 96436 24452 96440 24508
rect 96376 24448 96440 24452
rect 96456 24508 96520 24512
rect 96456 24452 96460 24508
rect 96460 24452 96516 24508
rect 96516 24452 96520 24508
rect 96456 24448 96520 24452
rect 96536 24508 96600 24512
rect 96536 24452 96540 24508
rect 96540 24452 96596 24508
rect 96596 24452 96600 24508
rect 96536 24448 96600 24452
rect 96616 24508 96680 24512
rect 96616 24452 96620 24508
rect 96620 24452 96676 24508
rect 96676 24452 96680 24508
rect 96616 24448 96680 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 81016 23964 81080 23968
rect 81016 23908 81020 23964
rect 81020 23908 81076 23964
rect 81076 23908 81080 23964
rect 81016 23904 81080 23908
rect 81096 23964 81160 23968
rect 81096 23908 81100 23964
rect 81100 23908 81156 23964
rect 81156 23908 81160 23964
rect 81096 23904 81160 23908
rect 81176 23964 81240 23968
rect 81176 23908 81180 23964
rect 81180 23908 81236 23964
rect 81236 23908 81240 23964
rect 81176 23904 81240 23908
rect 81256 23964 81320 23968
rect 81256 23908 81260 23964
rect 81260 23908 81316 23964
rect 81316 23908 81320 23964
rect 81256 23904 81320 23908
rect 111736 23964 111800 23968
rect 111736 23908 111740 23964
rect 111740 23908 111796 23964
rect 111796 23908 111800 23964
rect 111736 23904 111800 23908
rect 111816 23964 111880 23968
rect 111816 23908 111820 23964
rect 111820 23908 111876 23964
rect 111876 23908 111880 23964
rect 111816 23904 111880 23908
rect 111896 23964 111960 23968
rect 111896 23908 111900 23964
rect 111900 23908 111956 23964
rect 111956 23908 111960 23964
rect 111896 23904 111960 23908
rect 111976 23964 112040 23968
rect 111976 23908 111980 23964
rect 111980 23908 112036 23964
rect 112036 23908 112040 23964
rect 111976 23904 112040 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 96376 23420 96440 23424
rect 96376 23364 96380 23420
rect 96380 23364 96436 23420
rect 96436 23364 96440 23420
rect 96376 23360 96440 23364
rect 96456 23420 96520 23424
rect 96456 23364 96460 23420
rect 96460 23364 96516 23420
rect 96516 23364 96520 23420
rect 96456 23360 96520 23364
rect 96536 23420 96600 23424
rect 96536 23364 96540 23420
rect 96540 23364 96596 23420
rect 96596 23364 96600 23420
rect 96536 23360 96600 23364
rect 96616 23420 96680 23424
rect 96616 23364 96620 23420
rect 96620 23364 96676 23420
rect 96676 23364 96680 23420
rect 96616 23360 96680 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 81016 22876 81080 22880
rect 81016 22820 81020 22876
rect 81020 22820 81076 22876
rect 81076 22820 81080 22876
rect 81016 22816 81080 22820
rect 81096 22876 81160 22880
rect 81096 22820 81100 22876
rect 81100 22820 81156 22876
rect 81156 22820 81160 22876
rect 81096 22816 81160 22820
rect 81176 22876 81240 22880
rect 81176 22820 81180 22876
rect 81180 22820 81236 22876
rect 81236 22820 81240 22876
rect 81176 22816 81240 22820
rect 81256 22876 81320 22880
rect 81256 22820 81260 22876
rect 81260 22820 81316 22876
rect 81316 22820 81320 22876
rect 81256 22816 81320 22820
rect 111736 22876 111800 22880
rect 111736 22820 111740 22876
rect 111740 22820 111796 22876
rect 111796 22820 111800 22876
rect 111736 22816 111800 22820
rect 111816 22876 111880 22880
rect 111816 22820 111820 22876
rect 111820 22820 111876 22876
rect 111876 22820 111880 22876
rect 111816 22816 111880 22820
rect 111896 22876 111960 22880
rect 111896 22820 111900 22876
rect 111900 22820 111956 22876
rect 111956 22820 111960 22876
rect 111896 22816 111960 22820
rect 111976 22876 112040 22880
rect 111976 22820 111980 22876
rect 111980 22820 112036 22876
rect 112036 22820 112040 22876
rect 111976 22816 112040 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 96376 22332 96440 22336
rect 96376 22276 96380 22332
rect 96380 22276 96436 22332
rect 96436 22276 96440 22332
rect 96376 22272 96440 22276
rect 96456 22332 96520 22336
rect 96456 22276 96460 22332
rect 96460 22276 96516 22332
rect 96516 22276 96520 22332
rect 96456 22272 96520 22276
rect 96536 22332 96600 22336
rect 96536 22276 96540 22332
rect 96540 22276 96596 22332
rect 96596 22276 96600 22332
rect 96536 22272 96600 22276
rect 96616 22332 96680 22336
rect 96616 22276 96620 22332
rect 96620 22276 96676 22332
rect 96676 22276 96680 22332
rect 96616 22272 96680 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 81016 21788 81080 21792
rect 81016 21732 81020 21788
rect 81020 21732 81076 21788
rect 81076 21732 81080 21788
rect 81016 21728 81080 21732
rect 81096 21788 81160 21792
rect 81096 21732 81100 21788
rect 81100 21732 81156 21788
rect 81156 21732 81160 21788
rect 81096 21728 81160 21732
rect 81176 21788 81240 21792
rect 81176 21732 81180 21788
rect 81180 21732 81236 21788
rect 81236 21732 81240 21788
rect 81176 21728 81240 21732
rect 81256 21788 81320 21792
rect 81256 21732 81260 21788
rect 81260 21732 81316 21788
rect 81316 21732 81320 21788
rect 81256 21728 81320 21732
rect 111736 21788 111800 21792
rect 111736 21732 111740 21788
rect 111740 21732 111796 21788
rect 111796 21732 111800 21788
rect 111736 21728 111800 21732
rect 111816 21788 111880 21792
rect 111816 21732 111820 21788
rect 111820 21732 111876 21788
rect 111876 21732 111880 21788
rect 111816 21728 111880 21732
rect 111896 21788 111960 21792
rect 111896 21732 111900 21788
rect 111900 21732 111956 21788
rect 111956 21732 111960 21788
rect 111896 21728 111960 21732
rect 111976 21788 112040 21792
rect 111976 21732 111980 21788
rect 111980 21732 112036 21788
rect 112036 21732 112040 21788
rect 111976 21728 112040 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 96376 21244 96440 21248
rect 96376 21188 96380 21244
rect 96380 21188 96436 21244
rect 96436 21188 96440 21244
rect 96376 21184 96440 21188
rect 96456 21244 96520 21248
rect 96456 21188 96460 21244
rect 96460 21188 96516 21244
rect 96516 21188 96520 21244
rect 96456 21184 96520 21188
rect 96536 21244 96600 21248
rect 96536 21188 96540 21244
rect 96540 21188 96596 21244
rect 96596 21188 96600 21244
rect 96536 21184 96600 21188
rect 96616 21244 96680 21248
rect 96616 21188 96620 21244
rect 96620 21188 96676 21244
rect 96676 21188 96680 21244
rect 96616 21184 96680 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 81016 20700 81080 20704
rect 81016 20644 81020 20700
rect 81020 20644 81076 20700
rect 81076 20644 81080 20700
rect 81016 20640 81080 20644
rect 81096 20700 81160 20704
rect 81096 20644 81100 20700
rect 81100 20644 81156 20700
rect 81156 20644 81160 20700
rect 81096 20640 81160 20644
rect 81176 20700 81240 20704
rect 81176 20644 81180 20700
rect 81180 20644 81236 20700
rect 81236 20644 81240 20700
rect 81176 20640 81240 20644
rect 81256 20700 81320 20704
rect 81256 20644 81260 20700
rect 81260 20644 81316 20700
rect 81316 20644 81320 20700
rect 81256 20640 81320 20644
rect 111736 20700 111800 20704
rect 111736 20644 111740 20700
rect 111740 20644 111796 20700
rect 111796 20644 111800 20700
rect 111736 20640 111800 20644
rect 111816 20700 111880 20704
rect 111816 20644 111820 20700
rect 111820 20644 111876 20700
rect 111876 20644 111880 20700
rect 111816 20640 111880 20644
rect 111896 20700 111960 20704
rect 111896 20644 111900 20700
rect 111900 20644 111956 20700
rect 111956 20644 111960 20700
rect 111896 20640 111960 20644
rect 111976 20700 112040 20704
rect 111976 20644 111980 20700
rect 111980 20644 112036 20700
rect 112036 20644 112040 20700
rect 111976 20640 112040 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 96376 20156 96440 20160
rect 96376 20100 96380 20156
rect 96380 20100 96436 20156
rect 96436 20100 96440 20156
rect 96376 20096 96440 20100
rect 96456 20156 96520 20160
rect 96456 20100 96460 20156
rect 96460 20100 96516 20156
rect 96516 20100 96520 20156
rect 96456 20096 96520 20100
rect 96536 20156 96600 20160
rect 96536 20100 96540 20156
rect 96540 20100 96596 20156
rect 96596 20100 96600 20156
rect 96536 20096 96600 20100
rect 96616 20156 96680 20160
rect 96616 20100 96620 20156
rect 96620 20100 96676 20156
rect 96676 20100 96680 20156
rect 96616 20096 96680 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 81016 19612 81080 19616
rect 81016 19556 81020 19612
rect 81020 19556 81076 19612
rect 81076 19556 81080 19612
rect 81016 19552 81080 19556
rect 81096 19612 81160 19616
rect 81096 19556 81100 19612
rect 81100 19556 81156 19612
rect 81156 19556 81160 19612
rect 81096 19552 81160 19556
rect 81176 19612 81240 19616
rect 81176 19556 81180 19612
rect 81180 19556 81236 19612
rect 81236 19556 81240 19612
rect 81176 19552 81240 19556
rect 81256 19612 81320 19616
rect 81256 19556 81260 19612
rect 81260 19556 81316 19612
rect 81316 19556 81320 19612
rect 81256 19552 81320 19556
rect 111736 19612 111800 19616
rect 111736 19556 111740 19612
rect 111740 19556 111796 19612
rect 111796 19556 111800 19612
rect 111736 19552 111800 19556
rect 111816 19612 111880 19616
rect 111816 19556 111820 19612
rect 111820 19556 111876 19612
rect 111876 19556 111880 19612
rect 111816 19552 111880 19556
rect 111896 19612 111960 19616
rect 111896 19556 111900 19612
rect 111900 19556 111956 19612
rect 111956 19556 111960 19612
rect 111896 19552 111960 19556
rect 111976 19612 112040 19616
rect 111976 19556 111980 19612
rect 111980 19556 112036 19612
rect 112036 19556 112040 19612
rect 111976 19552 112040 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 96376 19068 96440 19072
rect 96376 19012 96380 19068
rect 96380 19012 96436 19068
rect 96436 19012 96440 19068
rect 96376 19008 96440 19012
rect 96456 19068 96520 19072
rect 96456 19012 96460 19068
rect 96460 19012 96516 19068
rect 96516 19012 96520 19068
rect 96456 19008 96520 19012
rect 96536 19068 96600 19072
rect 96536 19012 96540 19068
rect 96540 19012 96596 19068
rect 96596 19012 96600 19068
rect 96536 19008 96600 19012
rect 96616 19068 96680 19072
rect 96616 19012 96620 19068
rect 96620 19012 96676 19068
rect 96676 19012 96680 19068
rect 96616 19008 96680 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 81016 18524 81080 18528
rect 81016 18468 81020 18524
rect 81020 18468 81076 18524
rect 81076 18468 81080 18524
rect 81016 18464 81080 18468
rect 81096 18524 81160 18528
rect 81096 18468 81100 18524
rect 81100 18468 81156 18524
rect 81156 18468 81160 18524
rect 81096 18464 81160 18468
rect 81176 18524 81240 18528
rect 81176 18468 81180 18524
rect 81180 18468 81236 18524
rect 81236 18468 81240 18524
rect 81176 18464 81240 18468
rect 81256 18524 81320 18528
rect 81256 18468 81260 18524
rect 81260 18468 81316 18524
rect 81316 18468 81320 18524
rect 81256 18464 81320 18468
rect 111736 18524 111800 18528
rect 111736 18468 111740 18524
rect 111740 18468 111796 18524
rect 111796 18468 111800 18524
rect 111736 18464 111800 18468
rect 111816 18524 111880 18528
rect 111816 18468 111820 18524
rect 111820 18468 111876 18524
rect 111876 18468 111880 18524
rect 111816 18464 111880 18468
rect 111896 18524 111960 18528
rect 111896 18468 111900 18524
rect 111900 18468 111956 18524
rect 111956 18468 111960 18524
rect 111896 18464 111960 18468
rect 111976 18524 112040 18528
rect 111976 18468 111980 18524
rect 111980 18468 112036 18524
rect 112036 18468 112040 18524
rect 111976 18464 112040 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 96376 17980 96440 17984
rect 96376 17924 96380 17980
rect 96380 17924 96436 17980
rect 96436 17924 96440 17980
rect 96376 17920 96440 17924
rect 96456 17980 96520 17984
rect 96456 17924 96460 17980
rect 96460 17924 96516 17980
rect 96516 17924 96520 17980
rect 96456 17920 96520 17924
rect 96536 17980 96600 17984
rect 96536 17924 96540 17980
rect 96540 17924 96596 17980
rect 96596 17924 96600 17980
rect 96536 17920 96600 17924
rect 96616 17980 96680 17984
rect 96616 17924 96620 17980
rect 96620 17924 96676 17980
rect 96676 17924 96680 17980
rect 96616 17920 96680 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 81016 17436 81080 17440
rect 81016 17380 81020 17436
rect 81020 17380 81076 17436
rect 81076 17380 81080 17436
rect 81016 17376 81080 17380
rect 81096 17436 81160 17440
rect 81096 17380 81100 17436
rect 81100 17380 81156 17436
rect 81156 17380 81160 17436
rect 81096 17376 81160 17380
rect 81176 17436 81240 17440
rect 81176 17380 81180 17436
rect 81180 17380 81236 17436
rect 81236 17380 81240 17436
rect 81176 17376 81240 17380
rect 81256 17436 81320 17440
rect 81256 17380 81260 17436
rect 81260 17380 81316 17436
rect 81316 17380 81320 17436
rect 81256 17376 81320 17380
rect 111736 17436 111800 17440
rect 111736 17380 111740 17436
rect 111740 17380 111796 17436
rect 111796 17380 111800 17436
rect 111736 17376 111800 17380
rect 111816 17436 111880 17440
rect 111816 17380 111820 17436
rect 111820 17380 111876 17436
rect 111876 17380 111880 17436
rect 111816 17376 111880 17380
rect 111896 17436 111960 17440
rect 111896 17380 111900 17436
rect 111900 17380 111956 17436
rect 111956 17380 111960 17436
rect 111896 17376 111960 17380
rect 111976 17436 112040 17440
rect 111976 17380 111980 17436
rect 111980 17380 112036 17436
rect 112036 17380 112040 17436
rect 111976 17376 112040 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 96376 16892 96440 16896
rect 96376 16836 96380 16892
rect 96380 16836 96436 16892
rect 96436 16836 96440 16892
rect 96376 16832 96440 16836
rect 96456 16892 96520 16896
rect 96456 16836 96460 16892
rect 96460 16836 96516 16892
rect 96516 16836 96520 16892
rect 96456 16832 96520 16836
rect 96536 16892 96600 16896
rect 96536 16836 96540 16892
rect 96540 16836 96596 16892
rect 96596 16836 96600 16892
rect 96536 16832 96600 16836
rect 96616 16892 96680 16896
rect 96616 16836 96620 16892
rect 96620 16836 96676 16892
rect 96676 16836 96680 16892
rect 96616 16832 96680 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 81016 16348 81080 16352
rect 81016 16292 81020 16348
rect 81020 16292 81076 16348
rect 81076 16292 81080 16348
rect 81016 16288 81080 16292
rect 81096 16348 81160 16352
rect 81096 16292 81100 16348
rect 81100 16292 81156 16348
rect 81156 16292 81160 16348
rect 81096 16288 81160 16292
rect 81176 16348 81240 16352
rect 81176 16292 81180 16348
rect 81180 16292 81236 16348
rect 81236 16292 81240 16348
rect 81176 16288 81240 16292
rect 81256 16348 81320 16352
rect 81256 16292 81260 16348
rect 81260 16292 81316 16348
rect 81316 16292 81320 16348
rect 81256 16288 81320 16292
rect 111736 16348 111800 16352
rect 111736 16292 111740 16348
rect 111740 16292 111796 16348
rect 111796 16292 111800 16348
rect 111736 16288 111800 16292
rect 111816 16348 111880 16352
rect 111816 16292 111820 16348
rect 111820 16292 111876 16348
rect 111876 16292 111880 16348
rect 111816 16288 111880 16292
rect 111896 16348 111960 16352
rect 111896 16292 111900 16348
rect 111900 16292 111956 16348
rect 111956 16292 111960 16348
rect 111896 16288 111960 16292
rect 111976 16348 112040 16352
rect 111976 16292 111980 16348
rect 111980 16292 112036 16348
rect 112036 16292 112040 16348
rect 111976 16288 112040 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 96376 15804 96440 15808
rect 96376 15748 96380 15804
rect 96380 15748 96436 15804
rect 96436 15748 96440 15804
rect 96376 15744 96440 15748
rect 96456 15804 96520 15808
rect 96456 15748 96460 15804
rect 96460 15748 96516 15804
rect 96516 15748 96520 15804
rect 96456 15744 96520 15748
rect 96536 15804 96600 15808
rect 96536 15748 96540 15804
rect 96540 15748 96596 15804
rect 96596 15748 96600 15804
rect 96536 15744 96600 15748
rect 96616 15804 96680 15808
rect 96616 15748 96620 15804
rect 96620 15748 96676 15804
rect 96676 15748 96680 15804
rect 96616 15744 96680 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 81016 15260 81080 15264
rect 81016 15204 81020 15260
rect 81020 15204 81076 15260
rect 81076 15204 81080 15260
rect 81016 15200 81080 15204
rect 81096 15260 81160 15264
rect 81096 15204 81100 15260
rect 81100 15204 81156 15260
rect 81156 15204 81160 15260
rect 81096 15200 81160 15204
rect 81176 15260 81240 15264
rect 81176 15204 81180 15260
rect 81180 15204 81236 15260
rect 81236 15204 81240 15260
rect 81176 15200 81240 15204
rect 81256 15260 81320 15264
rect 81256 15204 81260 15260
rect 81260 15204 81316 15260
rect 81316 15204 81320 15260
rect 81256 15200 81320 15204
rect 111736 15260 111800 15264
rect 111736 15204 111740 15260
rect 111740 15204 111796 15260
rect 111796 15204 111800 15260
rect 111736 15200 111800 15204
rect 111816 15260 111880 15264
rect 111816 15204 111820 15260
rect 111820 15204 111876 15260
rect 111876 15204 111880 15260
rect 111816 15200 111880 15204
rect 111896 15260 111960 15264
rect 111896 15204 111900 15260
rect 111900 15204 111956 15260
rect 111956 15204 111960 15260
rect 111896 15200 111960 15204
rect 111976 15260 112040 15264
rect 111976 15204 111980 15260
rect 111980 15204 112036 15260
rect 112036 15204 112040 15260
rect 111976 15200 112040 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 96376 14716 96440 14720
rect 96376 14660 96380 14716
rect 96380 14660 96436 14716
rect 96436 14660 96440 14716
rect 96376 14656 96440 14660
rect 96456 14716 96520 14720
rect 96456 14660 96460 14716
rect 96460 14660 96516 14716
rect 96516 14660 96520 14716
rect 96456 14656 96520 14660
rect 96536 14716 96600 14720
rect 96536 14660 96540 14716
rect 96540 14660 96596 14716
rect 96596 14660 96600 14716
rect 96536 14656 96600 14660
rect 96616 14716 96680 14720
rect 96616 14660 96620 14716
rect 96620 14660 96676 14716
rect 96676 14660 96680 14716
rect 96616 14656 96680 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 81016 14172 81080 14176
rect 81016 14116 81020 14172
rect 81020 14116 81076 14172
rect 81076 14116 81080 14172
rect 81016 14112 81080 14116
rect 81096 14172 81160 14176
rect 81096 14116 81100 14172
rect 81100 14116 81156 14172
rect 81156 14116 81160 14172
rect 81096 14112 81160 14116
rect 81176 14172 81240 14176
rect 81176 14116 81180 14172
rect 81180 14116 81236 14172
rect 81236 14116 81240 14172
rect 81176 14112 81240 14116
rect 81256 14172 81320 14176
rect 81256 14116 81260 14172
rect 81260 14116 81316 14172
rect 81316 14116 81320 14172
rect 81256 14112 81320 14116
rect 111736 14172 111800 14176
rect 111736 14116 111740 14172
rect 111740 14116 111796 14172
rect 111796 14116 111800 14172
rect 111736 14112 111800 14116
rect 111816 14172 111880 14176
rect 111816 14116 111820 14172
rect 111820 14116 111876 14172
rect 111876 14116 111880 14172
rect 111816 14112 111880 14116
rect 111896 14172 111960 14176
rect 111896 14116 111900 14172
rect 111900 14116 111956 14172
rect 111956 14116 111960 14172
rect 111896 14112 111960 14116
rect 111976 14172 112040 14176
rect 111976 14116 111980 14172
rect 111980 14116 112036 14172
rect 112036 14116 112040 14172
rect 111976 14112 112040 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 96376 13628 96440 13632
rect 96376 13572 96380 13628
rect 96380 13572 96436 13628
rect 96436 13572 96440 13628
rect 96376 13568 96440 13572
rect 96456 13628 96520 13632
rect 96456 13572 96460 13628
rect 96460 13572 96516 13628
rect 96516 13572 96520 13628
rect 96456 13568 96520 13572
rect 96536 13628 96600 13632
rect 96536 13572 96540 13628
rect 96540 13572 96596 13628
rect 96596 13572 96600 13628
rect 96536 13568 96600 13572
rect 96616 13628 96680 13632
rect 96616 13572 96620 13628
rect 96620 13572 96676 13628
rect 96676 13572 96680 13628
rect 96616 13568 96680 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 81016 13084 81080 13088
rect 81016 13028 81020 13084
rect 81020 13028 81076 13084
rect 81076 13028 81080 13084
rect 81016 13024 81080 13028
rect 81096 13084 81160 13088
rect 81096 13028 81100 13084
rect 81100 13028 81156 13084
rect 81156 13028 81160 13084
rect 81096 13024 81160 13028
rect 81176 13084 81240 13088
rect 81176 13028 81180 13084
rect 81180 13028 81236 13084
rect 81236 13028 81240 13084
rect 81176 13024 81240 13028
rect 81256 13084 81320 13088
rect 81256 13028 81260 13084
rect 81260 13028 81316 13084
rect 81316 13028 81320 13084
rect 81256 13024 81320 13028
rect 111736 13084 111800 13088
rect 111736 13028 111740 13084
rect 111740 13028 111796 13084
rect 111796 13028 111800 13084
rect 111736 13024 111800 13028
rect 111816 13084 111880 13088
rect 111816 13028 111820 13084
rect 111820 13028 111876 13084
rect 111876 13028 111880 13084
rect 111816 13024 111880 13028
rect 111896 13084 111960 13088
rect 111896 13028 111900 13084
rect 111900 13028 111956 13084
rect 111956 13028 111960 13084
rect 111896 13024 111960 13028
rect 111976 13084 112040 13088
rect 111976 13028 111980 13084
rect 111980 13028 112036 13084
rect 112036 13028 112040 13084
rect 111976 13024 112040 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 96376 12540 96440 12544
rect 96376 12484 96380 12540
rect 96380 12484 96436 12540
rect 96436 12484 96440 12540
rect 96376 12480 96440 12484
rect 96456 12540 96520 12544
rect 96456 12484 96460 12540
rect 96460 12484 96516 12540
rect 96516 12484 96520 12540
rect 96456 12480 96520 12484
rect 96536 12540 96600 12544
rect 96536 12484 96540 12540
rect 96540 12484 96596 12540
rect 96596 12484 96600 12540
rect 96536 12480 96600 12484
rect 96616 12540 96680 12544
rect 96616 12484 96620 12540
rect 96620 12484 96676 12540
rect 96676 12484 96680 12540
rect 96616 12480 96680 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 81016 11996 81080 12000
rect 81016 11940 81020 11996
rect 81020 11940 81076 11996
rect 81076 11940 81080 11996
rect 81016 11936 81080 11940
rect 81096 11996 81160 12000
rect 81096 11940 81100 11996
rect 81100 11940 81156 11996
rect 81156 11940 81160 11996
rect 81096 11936 81160 11940
rect 81176 11996 81240 12000
rect 81176 11940 81180 11996
rect 81180 11940 81236 11996
rect 81236 11940 81240 11996
rect 81176 11936 81240 11940
rect 81256 11996 81320 12000
rect 81256 11940 81260 11996
rect 81260 11940 81316 11996
rect 81316 11940 81320 11996
rect 81256 11936 81320 11940
rect 111736 11996 111800 12000
rect 111736 11940 111740 11996
rect 111740 11940 111796 11996
rect 111796 11940 111800 11996
rect 111736 11936 111800 11940
rect 111816 11996 111880 12000
rect 111816 11940 111820 11996
rect 111820 11940 111876 11996
rect 111876 11940 111880 11996
rect 111816 11936 111880 11940
rect 111896 11996 111960 12000
rect 111896 11940 111900 11996
rect 111900 11940 111956 11996
rect 111956 11940 111960 11996
rect 111896 11936 111960 11940
rect 111976 11996 112040 12000
rect 111976 11940 111980 11996
rect 111980 11940 112036 11996
rect 112036 11940 112040 11996
rect 111976 11936 112040 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 96376 11452 96440 11456
rect 96376 11396 96380 11452
rect 96380 11396 96436 11452
rect 96436 11396 96440 11452
rect 96376 11392 96440 11396
rect 96456 11452 96520 11456
rect 96456 11396 96460 11452
rect 96460 11396 96516 11452
rect 96516 11396 96520 11452
rect 96456 11392 96520 11396
rect 96536 11452 96600 11456
rect 96536 11396 96540 11452
rect 96540 11396 96596 11452
rect 96596 11396 96600 11452
rect 96536 11392 96600 11396
rect 96616 11452 96680 11456
rect 96616 11396 96620 11452
rect 96620 11396 96676 11452
rect 96676 11396 96680 11452
rect 96616 11392 96680 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 81016 10908 81080 10912
rect 81016 10852 81020 10908
rect 81020 10852 81076 10908
rect 81076 10852 81080 10908
rect 81016 10848 81080 10852
rect 81096 10908 81160 10912
rect 81096 10852 81100 10908
rect 81100 10852 81156 10908
rect 81156 10852 81160 10908
rect 81096 10848 81160 10852
rect 81176 10908 81240 10912
rect 81176 10852 81180 10908
rect 81180 10852 81236 10908
rect 81236 10852 81240 10908
rect 81176 10848 81240 10852
rect 81256 10908 81320 10912
rect 81256 10852 81260 10908
rect 81260 10852 81316 10908
rect 81316 10852 81320 10908
rect 81256 10848 81320 10852
rect 111736 10908 111800 10912
rect 111736 10852 111740 10908
rect 111740 10852 111796 10908
rect 111796 10852 111800 10908
rect 111736 10848 111800 10852
rect 111816 10908 111880 10912
rect 111816 10852 111820 10908
rect 111820 10852 111876 10908
rect 111876 10852 111880 10908
rect 111816 10848 111880 10852
rect 111896 10908 111960 10912
rect 111896 10852 111900 10908
rect 111900 10852 111956 10908
rect 111956 10852 111960 10908
rect 111896 10848 111960 10852
rect 111976 10908 112040 10912
rect 111976 10852 111980 10908
rect 111980 10852 112036 10908
rect 112036 10852 112040 10908
rect 111976 10848 112040 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 96376 10364 96440 10368
rect 96376 10308 96380 10364
rect 96380 10308 96436 10364
rect 96436 10308 96440 10364
rect 96376 10304 96440 10308
rect 96456 10364 96520 10368
rect 96456 10308 96460 10364
rect 96460 10308 96516 10364
rect 96516 10308 96520 10364
rect 96456 10304 96520 10308
rect 96536 10364 96600 10368
rect 96536 10308 96540 10364
rect 96540 10308 96596 10364
rect 96596 10308 96600 10364
rect 96536 10304 96600 10308
rect 96616 10364 96680 10368
rect 96616 10308 96620 10364
rect 96620 10308 96676 10364
rect 96676 10308 96680 10364
rect 96616 10304 96680 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 81016 9820 81080 9824
rect 81016 9764 81020 9820
rect 81020 9764 81076 9820
rect 81076 9764 81080 9820
rect 81016 9760 81080 9764
rect 81096 9820 81160 9824
rect 81096 9764 81100 9820
rect 81100 9764 81156 9820
rect 81156 9764 81160 9820
rect 81096 9760 81160 9764
rect 81176 9820 81240 9824
rect 81176 9764 81180 9820
rect 81180 9764 81236 9820
rect 81236 9764 81240 9820
rect 81176 9760 81240 9764
rect 81256 9820 81320 9824
rect 81256 9764 81260 9820
rect 81260 9764 81316 9820
rect 81316 9764 81320 9820
rect 81256 9760 81320 9764
rect 111736 9820 111800 9824
rect 111736 9764 111740 9820
rect 111740 9764 111796 9820
rect 111796 9764 111800 9820
rect 111736 9760 111800 9764
rect 111816 9820 111880 9824
rect 111816 9764 111820 9820
rect 111820 9764 111876 9820
rect 111876 9764 111880 9820
rect 111816 9760 111880 9764
rect 111896 9820 111960 9824
rect 111896 9764 111900 9820
rect 111900 9764 111956 9820
rect 111956 9764 111960 9820
rect 111896 9760 111960 9764
rect 111976 9820 112040 9824
rect 111976 9764 111980 9820
rect 111980 9764 112036 9820
rect 112036 9764 112040 9820
rect 111976 9760 112040 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 96376 9276 96440 9280
rect 96376 9220 96380 9276
rect 96380 9220 96436 9276
rect 96436 9220 96440 9276
rect 96376 9216 96440 9220
rect 96456 9276 96520 9280
rect 96456 9220 96460 9276
rect 96460 9220 96516 9276
rect 96516 9220 96520 9276
rect 96456 9216 96520 9220
rect 96536 9276 96600 9280
rect 96536 9220 96540 9276
rect 96540 9220 96596 9276
rect 96596 9220 96600 9276
rect 96536 9216 96600 9220
rect 96616 9276 96680 9280
rect 96616 9220 96620 9276
rect 96620 9220 96676 9276
rect 96676 9220 96680 9276
rect 96616 9216 96680 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 81016 8732 81080 8736
rect 81016 8676 81020 8732
rect 81020 8676 81076 8732
rect 81076 8676 81080 8732
rect 81016 8672 81080 8676
rect 81096 8732 81160 8736
rect 81096 8676 81100 8732
rect 81100 8676 81156 8732
rect 81156 8676 81160 8732
rect 81096 8672 81160 8676
rect 81176 8732 81240 8736
rect 81176 8676 81180 8732
rect 81180 8676 81236 8732
rect 81236 8676 81240 8732
rect 81176 8672 81240 8676
rect 81256 8732 81320 8736
rect 81256 8676 81260 8732
rect 81260 8676 81316 8732
rect 81316 8676 81320 8732
rect 81256 8672 81320 8676
rect 111736 8732 111800 8736
rect 111736 8676 111740 8732
rect 111740 8676 111796 8732
rect 111796 8676 111800 8732
rect 111736 8672 111800 8676
rect 111816 8732 111880 8736
rect 111816 8676 111820 8732
rect 111820 8676 111876 8732
rect 111876 8676 111880 8732
rect 111816 8672 111880 8676
rect 111896 8732 111960 8736
rect 111896 8676 111900 8732
rect 111900 8676 111956 8732
rect 111956 8676 111960 8732
rect 111896 8672 111960 8676
rect 111976 8732 112040 8736
rect 111976 8676 111980 8732
rect 111980 8676 112036 8732
rect 112036 8676 112040 8732
rect 111976 8672 112040 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 96376 8188 96440 8192
rect 96376 8132 96380 8188
rect 96380 8132 96436 8188
rect 96436 8132 96440 8188
rect 96376 8128 96440 8132
rect 96456 8188 96520 8192
rect 96456 8132 96460 8188
rect 96460 8132 96516 8188
rect 96516 8132 96520 8188
rect 96456 8128 96520 8132
rect 96536 8188 96600 8192
rect 96536 8132 96540 8188
rect 96540 8132 96596 8188
rect 96596 8132 96600 8188
rect 96536 8128 96600 8132
rect 96616 8188 96680 8192
rect 96616 8132 96620 8188
rect 96620 8132 96676 8188
rect 96676 8132 96680 8188
rect 96616 8128 96680 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 81016 7644 81080 7648
rect 81016 7588 81020 7644
rect 81020 7588 81076 7644
rect 81076 7588 81080 7644
rect 81016 7584 81080 7588
rect 81096 7644 81160 7648
rect 81096 7588 81100 7644
rect 81100 7588 81156 7644
rect 81156 7588 81160 7644
rect 81096 7584 81160 7588
rect 81176 7644 81240 7648
rect 81176 7588 81180 7644
rect 81180 7588 81236 7644
rect 81236 7588 81240 7644
rect 81176 7584 81240 7588
rect 81256 7644 81320 7648
rect 81256 7588 81260 7644
rect 81260 7588 81316 7644
rect 81316 7588 81320 7644
rect 81256 7584 81320 7588
rect 111736 7644 111800 7648
rect 111736 7588 111740 7644
rect 111740 7588 111796 7644
rect 111796 7588 111800 7644
rect 111736 7584 111800 7588
rect 111816 7644 111880 7648
rect 111816 7588 111820 7644
rect 111820 7588 111876 7644
rect 111876 7588 111880 7644
rect 111816 7584 111880 7588
rect 111896 7644 111960 7648
rect 111896 7588 111900 7644
rect 111900 7588 111956 7644
rect 111956 7588 111960 7644
rect 111896 7584 111960 7588
rect 111976 7644 112040 7648
rect 111976 7588 111980 7644
rect 111980 7588 112036 7644
rect 112036 7588 112040 7644
rect 111976 7584 112040 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 96376 7100 96440 7104
rect 96376 7044 96380 7100
rect 96380 7044 96436 7100
rect 96436 7044 96440 7100
rect 96376 7040 96440 7044
rect 96456 7100 96520 7104
rect 96456 7044 96460 7100
rect 96460 7044 96516 7100
rect 96516 7044 96520 7100
rect 96456 7040 96520 7044
rect 96536 7100 96600 7104
rect 96536 7044 96540 7100
rect 96540 7044 96596 7100
rect 96596 7044 96600 7100
rect 96536 7040 96600 7044
rect 96616 7100 96680 7104
rect 96616 7044 96620 7100
rect 96620 7044 96676 7100
rect 96676 7044 96680 7100
rect 96616 7040 96680 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 81016 6556 81080 6560
rect 81016 6500 81020 6556
rect 81020 6500 81076 6556
rect 81076 6500 81080 6556
rect 81016 6496 81080 6500
rect 81096 6556 81160 6560
rect 81096 6500 81100 6556
rect 81100 6500 81156 6556
rect 81156 6500 81160 6556
rect 81096 6496 81160 6500
rect 81176 6556 81240 6560
rect 81176 6500 81180 6556
rect 81180 6500 81236 6556
rect 81236 6500 81240 6556
rect 81176 6496 81240 6500
rect 81256 6556 81320 6560
rect 81256 6500 81260 6556
rect 81260 6500 81316 6556
rect 81316 6500 81320 6556
rect 81256 6496 81320 6500
rect 111736 6556 111800 6560
rect 111736 6500 111740 6556
rect 111740 6500 111796 6556
rect 111796 6500 111800 6556
rect 111736 6496 111800 6500
rect 111816 6556 111880 6560
rect 111816 6500 111820 6556
rect 111820 6500 111876 6556
rect 111876 6500 111880 6556
rect 111816 6496 111880 6500
rect 111896 6556 111960 6560
rect 111896 6500 111900 6556
rect 111900 6500 111956 6556
rect 111956 6500 111960 6556
rect 111896 6496 111960 6500
rect 111976 6556 112040 6560
rect 111976 6500 111980 6556
rect 111980 6500 112036 6556
rect 112036 6500 112040 6556
rect 111976 6496 112040 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 96376 6012 96440 6016
rect 96376 5956 96380 6012
rect 96380 5956 96436 6012
rect 96436 5956 96440 6012
rect 96376 5952 96440 5956
rect 96456 6012 96520 6016
rect 96456 5956 96460 6012
rect 96460 5956 96516 6012
rect 96516 5956 96520 6012
rect 96456 5952 96520 5956
rect 96536 6012 96600 6016
rect 96536 5956 96540 6012
rect 96540 5956 96596 6012
rect 96596 5956 96600 6012
rect 96536 5952 96600 5956
rect 96616 6012 96680 6016
rect 96616 5956 96620 6012
rect 96620 5956 96676 6012
rect 96676 5956 96680 6012
rect 96616 5952 96680 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 81016 5468 81080 5472
rect 81016 5412 81020 5468
rect 81020 5412 81076 5468
rect 81076 5412 81080 5468
rect 81016 5408 81080 5412
rect 81096 5468 81160 5472
rect 81096 5412 81100 5468
rect 81100 5412 81156 5468
rect 81156 5412 81160 5468
rect 81096 5408 81160 5412
rect 81176 5468 81240 5472
rect 81176 5412 81180 5468
rect 81180 5412 81236 5468
rect 81236 5412 81240 5468
rect 81176 5408 81240 5412
rect 81256 5468 81320 5472
rect 81256 5412 81260 5468
rect 81260 5412 81316 5468
rect 81316 5412 81320 5468
rect 81256 5408 81320 5412
rect 111736 5468 111800 5472
rect 111736 5412 111740 5468
rect 111740 5412 111796 5468
rect 111796 5412 111800 5468
rect 111736 5408 111800 5412
rect 111816 5468 111880 5472
rect 111816 5412 111820 5468
rect 111820 5412 111876 5468
rect 111876 5412 111880 5468
rect 111816 5408 111880 5412
rect 111896 5468 111960 5472
rect 111896 5412 111900 5468
rect 111900 5412 111956 5468
rect 111956 5412 111960 5468
rect 111896 5408 111960 5412
rect 111976 5468 112040 5472
rect 111976 5412 111980 5468
rect 111980 5412 112036 5468
rect 112036 5412 112040 5468
rect 111976 5408 112040 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 96376 4924 96440 4928
rect 96376 4868 96380 4924
rect 96380 4868 96436 4924
rect 96436 4868 96440 4924
rect 96376 4864 96440 4868
rect 96456 4924 96520 4928
rect 96456 4868 96460 4924
rect 96460 4868 96516 4924
rect 96516 4868 96520 4924
rect 96456 4864 96520 4868
rect 96536 4924 96600 4928
rect 96536 4868 96540 4924
rect 96540 4868 96596 4924
rect 96596 4868 96600 4924
rect 96536 4864 96600 4868
rect 96616 4924 96680 4928
rect 96616 4868 96620 4924
rect 96620 4868 96676 4924
rect 96676 4868 96680 4924
rect 96616 4864 96680 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 81016 4380 81080 4384
rect 81016 4324 81020 4380
rect 81020 4324 81076 4380
rect 81076 4324 81080 4380
rect 81016 4320 81080 4324
rect 81096 4380 81160 4384
rect 81096 4324 81100 4380
rect 81100 4324 81156 4380
rect 81156 4324 81160 4380
rect 81096 4320 81160 4324
rect 81176 4380 81240 4384
rect 81176 4324 81180 4380
rect 81180 4324 81236 4380
rect 81236 4324 81240 4380
rect 81176 4320 81240 4324
rect 81256 4380 81320 4384
rect 81256 4324 81260 4380
rect 81260 4324 81316 4380
rect 81316 4324 81320 4380
rect 81256 4320 81320 4324
rect 111736 4380 111800 4384
rect 111736 4324 111740 4380
rect 111740 4324 111796 4380
rect 111796 4324 111800 4380
rect 111736 4320 111800 4324
rect 111816 4380 111880 4384
rect 111816 4324 111820 4380
rect 111820 4324 111876 4380
rect 111876 4324 111880 4380
rect 111816 4320 111880 4324
rect 111896 4380 111960 4384
rect 111896 4324 111900 4380
rect 111900 4324 111956 4380
rect 111956 4324 111960 4380
rect 111896 4320 111960 4324
rect 111976 4380 112040 4384
rect 111976 4324 111980 4380
rect 111980 4324 112036 4380
rect 112036 4324 112040 4380
rect 111976 4320 112040 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 96376 3836 96440 3840
rect 96376 3780 96380 3836
rect 96380 3780 96436 3836
rect 96436 3780 96440 3836
rect 96376 3776 96440 3780
rect 96456 3836 96520 3840
rect 96456 3780 96460 3836
rect 96460 3780 96516 3836
rect 96516 3780 96520 3836
rect 96456 3776 96520 3780
rect 96536 3836 96600 3840
rect 96536 3780 96540 3836
rect 96540 3780 96596 3836
rect 96596 3780 96600 3836
rect 96536 3776 96600 3780
rect 96616 3836 96680 3840
rect 96616 3780 96620 3836
rect 96620 3780 96676 3836
rect 96676 3780 96680 3836
rect 96616 3776 96680 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 81016 3292 81080 3296
rect 81016 3236 81020 3292
rect 81020 3236 81076 3292
rect 81076 3236 81080 3292
rect 81016 3232 81080 3236
rect 81096 3292 81160 3296
rect 81096 3236 81100 3292
rect 81100 3236 81156 3292
rect 81156 3236 81160 3292
rect 81096 3232 81160 3236
rect 81176 3292 81240 3296
rect 81176 3236 81180 3292
rect 81180 3236 81236 3292
rect 81236 3236 81240 3292
rect 81176 3232 81240 3236
rect 81256 3292 81320 3296
rect 81256 3236 81260 3292
rect 81260 3236 81316 3292
rect 81316 3236 81320 3292
rect 81256 3232 81320 3236
rect 111736 3292 111800 3296
rect 111736 3236 111740 3292
rect 111740 3236 111796 3292
rect 111796 3236 111800 3292
rect 111736 3232 111800 3236
rect 111816 3292 111880 3296
rect 111816 3236 111820 3292
rect 111820 3236 111876 3292
rect 111876 3236 111880 3292
rect 111816 3232 111880 3236
rect 111896 3292 111960 3296
rect 111896 3236 111900 3292
rect 111900 3236 111956 3292
rect 111956 3236 111960 3292
rect 111896 3232 111960 3236
rect 111976 3292 112040 3296
rect 111976 3236 111980 3292
rect 111980 3236 112036 3292
rect 112036 3236 112040 3292
rect 111976 3232 112040 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 96376 2748 96440 2752
rect 96376 2692 96380 2748
rect 96380 2692 96436 2748
rect 96436 2692 96440 2748
rect 96376 2688 96440 2692
rect 96456 2748 96520 2752
rect 96456 2692 96460 2748
rect 96460 2692 96516 2748
rect 96516 2692 96520 2748
rect 96456 2688 96520 2692
rect 96536 2748 96600 2752
rect 96536 2692 96540 2748
rect 96540 2692 96596 2748
rect 96596 2692 96600 2748
rect 96536 2688 96600 2692
rect 96616 2748 96680 2752
rect 96616 2692 96620 2748
rect 96620 2692 96676 2748
rect 96676 2692 96680 2748
rect 96616 2688 96680 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
rect 60596 2212 60660 2276
rect 81016 2204 81080 2208
rect 81016 2148 81020 2204
rect 81020 2148 81076 2204
rect 81076 2148 81080 2204
rect 81016 2144 81080 2148
rect 81096 2204 81160 2208
rect 81096 2148 81100 2204
rect 81100 2148 81156 2204
rect 81156 2148 81160 2204
rect 81096 2144 81160 2148
rect 81176 2204 81240 2208
rect 81176 2148 81180 2204
rect 81180 2148 81236 2204
rect 81236 2148 81240 2204
rect 81176 2144 81240 2148
rect 81256 2204 81320 2208
rect 81256 2148 81260 2204
rect 81260 2148 81316 2204
rect 81316 2148 81320 2204
rect 81256 2144 81320 2148
rect 111736 2204 111800 2208
rect 111736 2148 111740 2204
rect 111740 2148 111796 2204
rect 111796 2148 111800 2204
rect 111736 2144 111800 2148
rect 111816 2204 111880 2208
rect 111816 2148 111820 2204
rect 111820 2148 111876 2204
rect 111876 2148 111880 2204
rect 111816 2144 111880 2148
rect 111896 2204 111960 2208
rect 111896 2148 111900 2204
rect 111900 2148 111956 2204
rect 111956 2148 111960 2204
rect 111896 2144 111960 2148
rect 111976 2204 112040 2208
rect 111976 2148 111980 2204
rect 111980 2148 112036 2204
rect 112036 2148 112040 2204
rect 111976 2144 112040 2148
rect 60596 1940 60660 2004
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 37024 50608 37584
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 65648 37568 65968 37584
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 60595 2276 60661 2277
rect 60595 2212 60596 2276
rect 60660 2212 60661 2276
rect 60595 2211 60661 2212
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 60598 2005 60658 2211
rect 65648 2128 65968 2688
rect 81008 37024 81328 37584
rect 81008 36960 81016 37024
rect 81080 36960 81096 37024
rect 81160 36960 81176 37024
rect 81240 36960 81256 37024
rect 81320 36960 81328 37024
rect 81008 35936 81328 36960
rect 81008 35872 81016 35936
rect 81080 35872 81096 35936
rect 81160 35872 81176 35936
rect 81240 35872 81256 35936
rect 81320 35872 81328 35936
rect 81008 34848 81328 35872
rect 81008 34784 81016 34848
rect 81080 34784 81096 34848
rect 81160 34784 81176 34848
rect 81240 34784 81256 34848
rect 81320 34784 81328 34848
rect 81008 33760 81328 34784
rect 81008 33696 81016 33760
rect 81080 33696 81096 33760
rect 81160 33696 81176 33760
rect 81240 33696 81256 33760
rect 81320 33696 81328 33760
rect 81008 32672 81328 33696
rect 81008 32608 81016 32672
rect 81080 32608 81096 32672
rect 81160 32608 81176 32672
rect 81240 32608 81256 32672
rect 81320 32608 81328 32672
rect 81008 31584 81328 32608
rect 81008 31520 81016 31584
rect 81080 31520 81096 31584
rect 81160 31520 81176 31584
rect 81240 31520 81256 31584
rect 81320 31520 81328 31584
rect 81008 30496 81328 31520
rect 81008 30432 81016 30496
rect 81080 30432 81096 30496
rect 81160 30432 81176 30496
rect 81240 30432 81256 30496
rect 81320 30432 81328 30496
rect 81008 29408 81328 30432
rect 81008 29344 81016 29408
rect 81080 29344 81096 29408
rect 81160 29344 81176 29408
rect 81240 29344 81256 29408
rect 81320 29344 81328 29408
rect 81008 28320 81328 29344
rect 81008 28256 81016 28320
rect 81080 28256 81096 28320
rect 81160 28256 81176 28320
rect 81240 28256 81256 28320
rect 81320 28256 81328 28320
rect 81008 27232 81328 28256
rect 81008 27168 81016 27232
rect 81080 27168 81096 27232
rect 81160 27168 81176 27232
rect 81240 27168 81256 27232
rect 81320 27168 81328 27232
rect 81008 26144 81328 27168
rect 81008 26080 81016 26144
rect 81080 26080 81096 26144
rect 81160 26080 81176 26144
rect 81240 26080 81256 26144
rect 81320 26080 81328 26144
rect 81008 25056 81328 26080
rect 81008 24992 81016 25056
rect 81080 24992 81096 25056
rect 81160 24992 81176 25056
rect 81240 24992 81256 25056
rect 81320 24992 81328 25056
rect 81008 23968 81328 24992
rect 81008 23904 81016 23968
rect 81080 23904 81096 23968
rect 81160 23904 81176 23968
rect 81240 23904 81256 23968
rect 81320 23904 81328 23968
rect 81008 22880 81328 23904
rect 81008 22816 81016 22880
rect 81080 22816 81096 22880
rect 81160 22816 81176 22880
rect 81240 22816 81256 22880
rect 81320 22816 81328 22880
rect 81008 21792 81328 22816
rect 81008 21728 81016 21792
rect 81080 21728 81096 21792
rect 81160 21728 81176 21792
rect 81240 21728 81256 21792
rect 81320 21728 81328 21792
rect 81008 20704 81328 21728
rect 81008 20640 81016 20704
rect 81080 20640 81096 20704
rect 81160 20640 81176 20704
rect 81240 20640 81256 20704
rect 81320 20640 81328 20704
rect 81008 19616 81328 20640
rect 81008 19552 81016 19616
rect 81080 19552 81096 19616
rect 81160 19552 81176 19616
rect 81240 19552 81256 19616
rect 81320 19552 81328 19616
rect 81008 18528 81328 19552
rect 81008 18464 81016 18528
rect 81080 18464 81096 18528
rect 81160 18464 81176 18528
rect 81240 18464 81256 18528
rect 81320 18464 81328 18528
rect 81008 17440 81328 18464
rect 81008 17376 81016 17440
rect 81080 17376 81096 17440
rect 81160 17376 81176 17440
rect 81240 17376 81256 17440
rect 81320 17376 81328 17440
rect 81008 16352 81328 17376
rect 81008 16288 81016 16352
rect 81080 16288 81096 16352
rect 81160 16288 81176 16352
rect 81240 16288 81256 16352
rect 81320 16288 81328 16352
rect 81008 15264 81328 16288
rect 81008 15200 81016 15264
rect 81080 15200 81096 15264
rect 81160 15200 81176 15264
rect 81240 15200 81256 15264
rect 81320 15200 81328 15264
rect 81008 14176 81328 15200
rect 81008 14112 81016 14176
rect 81080 14112 81096 14176
rect 81160 14112 81176 14176
rect 81240 14112 81256 14176
rect 81320 14112 81328 14176
rect 81008 13088 81328 14112
rect 81008 13024 81016 13088
rect 81080 13024 81096 13088
rect 81160 13024 81176 13088
rect 81240 13024 81256 13088
rect 81320 13024 81328 13088
rect 81008 12000 81328 13024
rect 81008 11936 81016 12000
rect 81080 11936 81096 12000
rect 81160 11936 81176 12000
rect 81240 11936 81256 12000
rect 81320 11936 81328 12000
rect 81008 10912 81328 11936
rect 81008 10848 81016 10912
rect 81080 10848 81096 10912
rect 81160 10848 81176 10912
rect 81240 10848 81256 10912
rect 81320 10848 81328 10912
rect 81008 9824 81328 10848
rect 81008 9760 81016 9824
rect 81080 9760 81096 9824
rect 81160 9760 81176 9824
rect 81240 9760 81256 9824
rect 81320 9760 81328 9824
rect 81008 8736 81328 9760
rect 81008 8672 81016 8736
rect 81080 8672 81096 8736
rect 81160 8672 81176 8736
rect 81240 8672 81256 8736
rect 81320 8672 81328 8736
rect 81008 7648 81328 8672
rect 81008 7584 81016 7648
rect 81080 7584 81096 7648
rect 81160 7584 81176 7648
rect 81240 7584 81256 7648
rect 81320 7584 81328 7648
rect 81008 6560 81328 7584
rect 81008 6496 81016 6560
rect 81080 6496 81096 6560
rect 81160 6496 81176 6560
rect 81240 6496 81256 6560
rect 81320 6496 81328 6560
rect 81008 5472 81328 6496
rect 81008 5408 81016 5472
rect 81080 5408 81096 5472
rect 81160 5408 81176 5472
rect 81240 5408 81256 5472
rect 81320 5408 81328 5472
rect 81008 4384 81328 5408
rect 81008 4320 81016 4384
rect 81080 4320 81096 4384
rect 81160 4320 81176 4384
rect 81240 4320 81256 4384
rect 81320 4320 81328 4384
rect 81008 3296 81328 4320
rect 81008 3232 81016 3296
rect 81080 3232 81096 3296
rect 81160 3232 81176 3296
rect 81240 3232 81256 3296
rect 81320 3232 81328 3296
rect 81008 2208 81328 3232
rect 81008 2144 81016 2208
rect 81080 2144 81096 2208
rect 81160 2144 81176 2208
rect 81240 2144 81256 2208
rect 81320 2144 81328 2208
rect 81008 2128 81328 2144
rect 96368 37568 96688 37584
rect 96368 37504 96376 37568
rect 96440 37504 96456 37568
rect 96520 37504 96536 37568
rect 96600 37504 96616 37568
rect 96680 37504 96688 37568
rect 96368 36480 96688 37504
rect 96368 36416 96376 36480
rect 96440 36416 96456 36480
rect 96520 36416 96536 36480
rect 96600 36416 96616 36480
rect 96680 36416 96688 36480
rect 96368 35392 96688 36416
rect 96368 35328 96376 35392
rect 96440 35328 96456 35392
rect 96520 35328 96536 35392
rect 96600 35328 96616 35392
rect 96680 35328 96688 35392
rect 96368 34304 96688 35328
rect 96368 34240 96376 34304
rect 96440 34240 96456 34304
rect 96520 34240 96536 34304
rect 96600 34240 96616 34304
rect 96680 34240 96688 34304
rect 96368 33216 96688 34240
rect 96368 33152 96376 33216
rect 96440 33152 96456 33216
rect 96520 33152 96536 33216
rect 96600 33152 96616 33216
rect 96680 33152 96688 33216
rect 96368 32128 96688 33152
rect 96368 32064 96376 32128
rect 96440 32064 96456 32128
rect 96520 32064 96536 32128
rect 96600 32064 96616 32128
rect 96680 32064 96688 32128
rect 96368 31040 96688 32064
rect 96368 30976 96376 31040
rect 96440 30976 96456 31040
rect 96520 30976 96536 31040
rect 96600 30976 96616 31040
rect 96680 30976 96688 31040
rect 96368 29952 96688 30976
rect 96368 29888 96376 29952
rect 96440 29888 96456 29952
rect 96520 29888 96536 29952
rect 96600 29888 96616 29952
rect 96680 29888 96688 29952
rect 96368 28864 96688 29888
rect 96368 28800 96376 28864
rect 96440 28800 96456 28864
rect 96520 28800 96536 28864
rect 96600 28800 96616 28864
rect 96680 28800 96688 28864
rect 96368 27776 96688 28800
rect 96368 27712 96376 27776
rect 96440 27712 96456 27776
rect 96520 27712 96536 27776
rect 96600 27712 96616 27776
rect 96680 27712 96688 27776
rect 96368 26688 96688 27712
rect 96368 26624 96376 26688
rect 96440 26624 96456 26688
rect 96520 26624 96536 26688
rect 96600 26624 96616 26688
rect 96680 26624 96688 26688
rect 96368 25600 96688 26624
rect 96368 25536 96376 25600
rect 96440 25536 96456 25600
rect 96520 25536 96536 25600
rect 96600 25536 96616 25600
rect 96680 25536 96688 25600
rect 96368 24512 96688 25536
rect 96368 24448 96376 24512
rect 96440 24448 96456 24512
rect 96520 24448 96536 24512
rect 96600 24448 96616 24512
rect 96680 24448 96688 24512
rect 96368 23424 96688 24448
rect 96368 23360 96376 23424
rect 96440 23360 96456 23424
rect 96520 23360 96536 23424
rect 96600 23360 96616 23424
rect 96680 23360 96688 23424
rect 96368 22336 96688 23360
rect 96368 22272 96376 22336
rect 96440 22272 96456 22336
rect 96520 22272 96536 22336
rect 96600 22272 96616 22336
rect 96680 22272 96688 22336
rect 96368 21248 96688 22272
rect 96368 21184 96376 21248
rect 96440 21184 96456 21248
rect 96520 21184 96536 21248
rect 96600 21184 96616 21248
rect 96680 21184 96688 21248
rect 96368 20160 96688 21184
rect 96368 20096 96376 20160
rect 96440 20096 96456 20160
rect 96520 20096 96536 20160
rect 96600 20096 96616 20160
rect 96680 20096 96688 20160
rect 96368 19072 96688 20096
rect 96368 19008 96376 19072
rect 96440 19008 96456 19072
rect 96520 19008 96536 19072
rect 96600 19008 96616 19072
rect 96680 19008 96688 19072
rect 96368 17984 96688 19008
rect 96368 17920 96376 17984
rect 96440 17920 96456 17984
rect 96520 17920 96536 17984
rect 96600 17920 96616 17984
rect 96680 17920 96688 17984
rect 96368 16896 96688 17920
rect 96368 16832 96376 16896
rect 96440 16832 96456 16896
rect 96520 16832 96536 16896
rect 96600 16832 96616 16896
rect 96680 16832 96688 16896
rect 96368 15808 96688 16832
rect 96368 15744 96376 15808
rect 96440 15744 96456 15808
rect 96520 15744 96536 15808
rect 96600 15744 96616 15808
rect 96680 15744 96688 15808
rect 96368 14720 96688 15744
rect 96368 14656 96376 14720
rect 96440 14656 96456 14720
rect 96520 14656 96536 14720
rect 96600 14656 96616 14720
rect 96680 14656 96688 14720
rect 96368 13632 96688 14656
rect 96368 13568 96376 13632
rect 96440 13568 96456 13632
rect 96520 13568 96536 13632
rect 96600 13568 96616 13632
rect 96680 13568 96688 13632
rect 96368 12544 96688 13568
rect 96368 12480 96376 12544
rect 96440 12480 96456 12544
rect 96520 12480 96536 12544
rect 96600 12480 96616 12544
rect 96680 12480 96688 12544
rect 96368 11456 96688 12480
rect 96368 11392 96376 11456
rect 96440 11392 96456 11456
rect 96520 11392 96536 11456
rect 96600 11392 96616 11456
rect 96680 11392 96688 11456
rect 96368 10368 96688 11392
rect 96368 10304 96376 10368
rect 96440 10304 96456 10368
rect 96520 10304 96536 10368
rect 96600 10304 96616 10368
rect 96680 10304 96688 10368
rect 96368 9280 96688 10304
rect 96368 9216 96376 9280
rect 96440 9216 96456 9280
rect 96520 9216 96536 9280
rect 96600 9216 96616 9280
rect 96680 9216 96688 9280
rect 96368 8192 96688 9216
rect 96368 8128 96376 8192
rect 96440 8128 96456 8192
rect 96520 8128 96536 8192
rect 96600 8128 96616 8192
rect 96680 8128 96688 8192
rect 96368 7104 96688 8128
rect 96368 7040 96376 7104
rect 96440 7040 96456 7104
rect 96520 7040 96536 7104
rect 96600 7040 96616 7104
rect 96680 7040 96688 7104
rect 96368 6016 96688 7040
rect 96368 5952 96376 6016
rect 96440 5952 96456 6016
rect 96520 5952 96536 6016
rect 96600 5952 96616 6016
rect 96680 5952 96688 6016
rect 96368 4928 96688 5952
rect 96368 4864 96376 4928
rect 96440 4864 96456 4928
rect 96520 4864 96536 4928
rect 96600 4864 96616 4928
rect 96680 4864 96688 4928
rect 96368 3840 96688 4864
rect 96368 3776 96376 3840
rect 96440 3776 96456 3840
rect 96520 3776 96536 3840
rect 96600 3776 96616 3840
rect 96680 3776 96688 3840
rect 96368 2752 96688 3776
rect 96368 2688 96376 2752
rect 96440 2688 96456 2752
rect 96520 2688 96536 2752
rect 96600 2688 96616 2752
rect 96680 2688 96688 2752
rect 96368 2128 96688 2688
rect 111728 37024 112048 37584
rect 111728 36960 111736 37024
rect 111800 36960 111816 37024
rect 111880 36960 111896 37024
rect 111960 36960 111976 37024
rect 112040 36960 112048 37024
rect 111728 35936 112048 36960
rect 111728 35872 111736 35936
rect 111800 35872 111816 35936
rect 111880 35872 111896 35936
rect 111960 35872 111976 35936
rect 112040 35872 112048 35936
rect 111728 34848 112048 35872
rect 111728 34784 111736 34848
rect 111800 34784 111816 34848
rect 111880 34784 111896 34848
rect 111960 34784 111976 34848
rect 112040 34784 112048 34848
rect 111728 33760 112048 34784
rect 111728 33696 111736 33760
rect 111800 33696 111816 33760
rect 111880 33696 111896 33760
rect 111960 33696 111976 33760
rect 112040 33696 112048 33760
rect 111728 32672 112048 33696
rect 111728 32608 111736 32672
rect 111800 32608 111816 32672
rect 111880 32608 111896 32672
rect 111960 32608 111976 32672
rect 112040 32608 112048 32672
rect 111728 31584 112048 32608
rect 111728 31520 111736 31584
rect 111800 31520 111816 31584
rect 111880 31520 111896 31584
rect 111960 31520 111976 31584
rect 112040 31520 112048 31584
rect 111728 30496 112048 31520
rect 111728 30432 111736 30496
rect 111800 30432 111816 30496
rect 111880 30432 111896 30496
rect 111960 30432 111976 30496
rect 112040 30432 112048 30496
rect 111728 29408 112048 30432
rect 111728 29344 111736 29408
rect 111800 29344 111816 29408
rect 111880 29344 111896 29408
rect 111960 29344 111976 29408
rect 112040 29344 112048 29408
rect 111728 28320 112048 29344
rect 111728 28256 111736 28320
rect 111800 28256 111816 28320
rect 111880 28256 111896 28320
rect 111960 28256 111976 28320
rect 112040 28256 112048 28320
rect 111728 27232 112048 28256
rect 111728 27168 111736 27232
rect 111800 27168 111816 27232
rect 111880 27168 111896 27232
rect 111960 27168 111976 27232
rect 112040 27168 112048 27232
rect 111728 26144 112048 27168
rect 111728 26080 111736 26144
rect 111800 26080 111816 26144
rect 111880 26080 111896 26144
rect 111960 26080 111976 26144
rect 112040 26080 112048 26144
rect 111728 25056 112048 26080
rect 111728 24992 111736 25056
rect 111800 24992 111816 25056
rect 111880 24992 111896 25056
rect 111960 24992 111976 25056
rect 112040 24992 112048 25056
rect 111728 23968 112048 24992
rect 111728 23904 111736 23968
rect 111800 23904 111816 23968
rect 111880 23904 111896 23968
rect 111960 23904 111976 23968
rect 112040 23904 112048 23968
rect 111728 22880 112048 23904
rect 111728 22816 111736 22880
rect 111800 22816 111816 22880
rect 111880 22816 111896 22880
rect 111960 22816 111976 22880
rect 112040 22816 112048 22880
rect 111728 21792 112048 22816
rect 111728 21728 111736 21792
rect 111800 21728 111816 21792
rect 111880 21728 111896 21792
rect 111960 21728 111976 21792
rect 112040 21728 112048 21792
rect 111728 20704 112048 21728
rect 111728 20640 111736 20704
rect 111800 20640 111816 20704
rect 111880 20640 111896 20704
rect 111960 20640 111976 20704
rect 112040 20640 112048 20704
rect 111728 19616 112048 20640
rect 111728 19552 111736 19616
rect 111800 19552 111816 19616
rect 111880 19552 111896 19616
rect 111960 19552 111976 19616
rect 112040 19552 112048 19616
rect 111728 18528 112048 19552
rect 111728 18464 111736 18528
rect 111800 18464 111816 18528
rect 111880 18464 111896 18528
rect 111960 18464 111976 18528
rect 112040 18464 112048 18528
rect 111728 17440 112048 18464
rect 111728 17376 111736 17440
rect 111800 17376 111816 17440
rect 111880 17376 111896 17440
rect 111960 17376 111976 17440
rect 112040 17376 112048 17440
rect 111728 16352 112048 17376
rect 111728 16288 111736 16352
rect 111800 16288 111816 16352
rect 111880 16288 111896 16352
rect 111960 16288 111976 16352
rect 112040 16288 112048 16352
rect 111728 15264 112048 16288
rect 111728 15200 111736 15264
rect 111800 15200 111816 15264
rect 111880 15200 111896 15264
rect 111960 15200 111976 15264
rect 112040 15200 112048 15264
rect 111728 14176 112048 15200
rect 111728 14112 111736 14176
rect 111800 14112 111816 14176
rect 111880 14112 111896 14176
rect 111960 14112 111976 14176
rect 112040 14112 112048 14176
rect 111728 13088 112048 14112
rect 111728 13024 111736 13088
rect 111800 13024 111816 13088
rect 111880 13024 111896 13088
rect 111960 13024 111976 13088
rect 112040 13024 112048 13088
rect 111728 12000 112048 13024
rect 111728 11936 111736 12000
rect 111800 11936 111816 12000
rect 111880 11936 111896 12000
rect 111960 11936 111976 12000
rect 112040 11936 112048 12000
rect 111728 10912 112048 11936
rect 111728 10848 111736 10912
rect 111800 10848 111816 10912
rect 111880 10848 111896 10912
rect 111960 10848 111976 10912
rect 112040 10848 112048 10912
rect 111728 9824 112048 10848
rect 111728 9760 111736 9824
rect 111800 9760 111816 9824
rect 111880 9760 111896 9824
rect 111960 9760 111976 9824
rect 112040 9760 112048 9824
rect 111728 8736 112048 9760
rect 111728 8672 111736 8736
rect 111800 8672 111816 8736
rect 111880 8672 111896 8736
rect 111960 8672 111976 8736
rect 112040 8672 112048 8736
rect 111728 7648 112048 8672
rect 111728 7584 111736 7648
rect 111800 7584 111816 7648
rect 111880 7584 111896 7648
rect 111960 7584 111976 7648
rect 112040 7584 112048 7648
rect 111728 6560 112048 7584
rect 111728 6496 111736 6560
rect 111800 6496 111816 6560
rect 111880 6496 111896 6560
rect 111960 6496 111976 6560
rect 112040 6496 112048 6560
rect 111728 5472 112048 6496
rect 111728 5408 111736 5472
rect 111800 5408 111816 5472
rect 111880 5408 111896 5472
rect 111960 5408 111976 5472
rect 112040 5408 112048 5472
rect 111728 4384 112048 5408
rect 111728 4320 111736 4384
rect 111800 4320 111816 4384
rect 111880 4320 111896 4384
rect 111960 4320 111976 4384
rect 112040 4320 112048 4384
rect 111728 3296 112048 4320
rect 111728 3232 111736 3296
rect 111800 3232 111816 3296
rect 111880 3232 111896 3296
rect 111960 3232 111976 3296
rect 112040 3232 112048 3296
rect 111728 2208 112048 3232
rect 111728 2144 111736 2208
rect 111800 2144 111816 2208
rect 111880 2144 111896 2208
rect 111960 2144 111976 2208
rect 112040 2144 112048 2208
rect 111728 2128 112048 2144
rect 60595 2004 60661 2005
rect 60595 1940 60596 2004
rect 60660 1940 60661 2004
rect 60595 1939 60661 1940
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 117484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 117484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 117484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 117484 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 117484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 117484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 117484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 117484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1644511149
transform 1 0 117484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1644511149
transform 1 0 117484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1644511149
transform 1 0 117484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1644511149
transform 1 0 117484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1644511149
transform 1 0 117484 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1644511149
transform -1 0 92000 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1644511149
transform -1 0 93380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1644511149
transform -1 0 91632 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1644511149
transform 1 0 34868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1644511149
transform -1 0 100280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1644511149
transform -1 0 105432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1644511149
transform -1 0 108468 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1644511149
transform -1 0 111688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1644511149
transform -1 0 116104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1644511149
transform -1 0 116472 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1644511149
transform 1 0 115460 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1644511149
transform 1 0 116840 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1644511149
transform 1 0 115092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1644511149
transform 1 0 56028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1644511149
transform 1 0 57132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1644511149
transform 1 0 55660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1644511149
transform 1 0 100096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1644511149
transform -1 0 82248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1644511149
transform -1 0 80776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1644511149
transform -1 0 82616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1644511149
transform 1 0 21988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1644511149
transform -1 0 65320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1644511149
transform -1 0 7176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1644511149
transform -1 0 67528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1644511149
transform -1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1644511149
transform -1 0 69092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1644511149
transform -1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1644511149
transform -1 0 70380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1644511149
transform -1 0 10488 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1644511149
transform 1 0 117484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1644511149
transform 1 0 117484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1644511149
transform 1 0 117484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1644511149
transform 1 0 117484 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1644511149
transform 1 0 110400 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1644511149
transform 1 0 79672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1644511149
transform 1 0 65412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1644511149
transform 1 0 66792 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1644511149
transform 1 0 68264 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1644511149
transform 1 0 69644 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46
timestamp 1644511149
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62
timestamp 1644511149
transform 1 0 6808 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71
timestamp 1644511149
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1644511149
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_93
timestamp 1644511149
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_97
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_102
timestamp 1644511149
transform 1 0 10488 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1644511149
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1644511149
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_124
timestamp 1644511149
transform 1 0 12512 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_157
timestamp 1644511149
transform 1 0 15548 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_175
timestamp 1644511149
transform 1 0 17204 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1644511149
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1644511149
transform 1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1644511149
transform 1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_211
timestamp 1644511149
transform 1 0 20516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1644511149
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_235
timestamp 1644511149
transform 1 0 22724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1644511149
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_259
timestamp 1644511149
transform 1 0 24932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_269
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_287
timestamp 1644511149
transform 1 0 27508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_297
timestamp 1644511149
transform 1 0 28428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_315
timestamp 1644511149
transform 1 0 30084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1644511149
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_343
timestamp 1644511149
transform 1 0 32660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_347
timestamp 1644511149
transform 1 0 33028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_351
timestamp 1644511149
transform 1 0 33396 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1644511149
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1644511149
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_375
timestamp 1644511149
transform 1 0 35604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_387
timestamp 1644511149
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_399
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_409
timestamp 1644511149
transform 1 0 38732 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 1644511149
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_427
timestamp 1644511149
transform 1 0 40388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_437
timestamp 1644511149
transform 1 0 41308 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_455
timestamp 1644511149
transform 1 0 42964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_467
timestamp 1644511149
transform 1 0 44068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1644511149
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_483
timestamp 1644511149
transform 1 0 45540 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_491
timestamp 1644511149
transform 1 0 46276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_498
timestamp 1644511149
transform 1 0 46920 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_514
timestamp 1644511149
transform 1 0 48392 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_528
timestamp 1644511149
transform 1 0 49680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_545
timestamp 1644511149
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1644511149
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_567
timestamp 1644511149
transform 1 0 53268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_577
timestamp 1644511149
transform 1 0 54188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 1644511149
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_589
timestamp 1644511149
transform 1 0 55292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_595
timestamp 1644511149
transform 1 0 55844 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_599
timestamp 1644511149
transform 1 0 56212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_607
timestamp 1644511149
transform 1 0 56948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_611
timestamp 1644511149
transform 1 0 57316 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1644511149
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_623
timestamp 1644511149
transform 1 0 58420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_631
timestamp 1644511149
transform 1 0 59156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_640
timestamp 1644511149
transform 1 0 59984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_645
timestamp 1644511149
transform 1 0 60444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_649
timestamp 1644511149
transform 1 0 60812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_656
timestamp 1644511149
transform 1 0 61456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_662
timestamp 1644511149
transform 1 0 62008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_667
timestamp 1644511149
transform 1 0 62468 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_671
timestamp 1644511149
transform 1 0 62836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_679
timestamp 1644511149
transform 1 0 63572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_689
timestamp 1644511149
transform 1 0 64492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_694
timestamp 1644511149
transform 1 0 64952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_698
timestamp 1644511149
transform 1 0 65320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_707
timestamp 1644511149
transform 1 0 66148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_711
timestamp 1644511149
transform 1 0 66516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_718
timestamp 1644511149
transform 1 0 67160 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_722
timestamp 1644511149
transform 1 0 67528 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_735
timestamp 1644511149
transform 1 0 68724 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_739
timestamp 1644511149
transform 1 0 69092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_749
timestamp 1644511149
transform 1 0 70012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_753
timestamp 1644511149
transform 1 0 70380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_757
timestamp 1644511149
transform 1 0 70748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_765
timestamp 1644511149
transform 1 0 71484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_773
timestamp 1644511149
transform 1 0 72220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_780
timestamp 1644511149
transform 1 0 72864 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_785
timestamp 1644511149
transform 1 0 73324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_791
timestamp 1644511149
transform 1 0 73876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_808
timestamp 1644511149
transform 1 0 75440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_822
timestamp 1644511149
transform 1 0 76728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_826
timestamp 1644511149
transform 1 0 77096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_836
timestamp 1644511149
transform 1 0 78016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_841
timestamp 1644511149
transform 1 0 78476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_852
timestamp 1644511149
transform 1 0 79488 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_859
timestamp 1644511149
transform 1 0 80132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_863
timestamp 1644511149
transform 1 0 80500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_866
timestamp 1644511149
transform 1 0 80776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_878
timestamp 1644511149
transform 1 0 81880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_882
timestamp 1644511149
transform 1 0 82248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_895
timestamp 1644511149
transform 1 0 83444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_906
timestamp 1644511149
transform 1 0 84456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_919
timestamp 1644511149
transform 1 0 85652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_923
timestamp 1644511149
transform 1 0 86020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_934
timestamp 1644511149
transform 1 0 87032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_938
timestamp 1644511149
transform 1 0 87400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_948
timestamp 1644511149
transform 1 0 88320 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_962
timestamp 1644511149
transform 1 0 89608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_966
timestamp 1644511149
transform 1 0 89976 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_976
timestamp 1644511149
transform 1 0 90896 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_981
timestamp 1644511149
transform 1 0 91356 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_992
timestamp 1644511149
transform 1 0 92368 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1002
timestamp 1644511149
transform 1 0 93288 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1012
timestamp 1644511149
transform 1 0 94208 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1020
timestamp 1644511149
transform 1 0 94944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1030
timestamp 1644511149
transform 1 0 95864 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1046
timestamp 1644511149
transform 1 0 97336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1059
timestamp 1644511149
transform 1 0 98532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1063
timestamp 1644511149
transform 1 0 98900 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1074
timestamp 1644511149
transform 1 0 99912 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1087
timestamp 1644511149
transform 1 0 101108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1091
timestamp 1644511149
transform 1 0 101476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1102
timestamp 1644511149
transform 1 0 102488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1115
timestamp 1644511149
transform 1 0 103684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1119
timestamp 1644511149
transform 1 0 104052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1124
timestamp 1644511149
transform 1 0 104512 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1139
timestamp 1644511149
transform 1 0 105892 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1147
timestamp 1644511149
transform 1 0 106628 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1149
timestamp 1644511149
transform 1 0 106812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1153
timestamp 1644511149
transform 1 0 107180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1163
timestamp 1644511149
transform 1 0 108100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1167
timestamp 1644511149
transform 1 0 108468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1172
timestamp 1644511149
transform 1 0 108928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1186
timestamp 1644511149
transform 1 0 110216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1193
timestamp 1644511149
transform 1 0 110860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1198
timestamp 1644511149
transform 1 0 111320 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1202
timestamp 1644511149
transform 1 0 111688 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1214
timestamp 1644511149
transform 1 0 112792 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1218
timestamp 1644511149
transform 1 0 113160 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1228
timestamp 1644511149
transform 1 0 114080 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1233
timestamp 1644511149
transform 1 0 114540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1246
timestamp 1644511149
transform 1 0 115736 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1250
timestamp 1644511149
transform 1 0 116104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1261
timestamp 1644511149
transform 1 0 117116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1273
timestamp 1644511149
transform 1 0 118220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_417
timestamp 1644511149
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_429
timestamp 1644511149
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1644511149
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1644511149
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_449
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_461
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_473
timestamp 1644511149
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1644511149
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1644511149
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_541
timestamp 1644511149
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1644511149
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1644511149
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_573
timestamp 1644511149
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1644511149
transform 1 0 54924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_595
timestamp 1644511149
transform 1 0 55844 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_607
timestamp 1644511149
transform 1 0 56948 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1644511149
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_617
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_629
timestamp 1644511149
transform 1 0 58972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_636
timestamp 1644511149
transform 1 0 59616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_640
timestamp 1644511149
transform 1 0 59984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_644
timestamp 1644511149
transform 1 0 60352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_652
timestamp 1644511149
transform 1 0 61088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_659
timestamp 1644511149
transform 1 0 61732 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1644511149
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_673
timestamp 1644511149
transform 1 0 63020 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_683
timestamp 1644511149
transform 1 0 63940 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_691
timestamp 1644511149
transform 1 0 64676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_697
timestamp 1644511149
transform 1 0 65228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_701
timestamp 1644511149
transform 1 0 65596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_706
timestamp 1644511149
transform 1 0 66056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_712
timestamp 1644511149
transform 1 0 66608 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_716
timestamp 1644511149
transform 1 0 66976 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1644511149
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1644511149
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_733
timestamp 1644511149
transform 1 0 68540 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_743
timestamp 1644511149
transform 1 0 69460 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_747
timestamp 1644511149
transform 1 0 69828 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_752
timestamp 1644511149
transform 1 0 70288 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_760
timestamp 1644511149
transform 1 0 71024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_764
timestamp 1644511149
transform 1 0 71392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_768
timestamp 1644511149
transform 1 0 71760 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_776
timestamp 1644511149
transform 1 0 72496 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_788
timestamp 1644511149
transform 1 0 73600 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_800
timestamp 1644511149
transform 1 0 74704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_806
timestamp 1644511149
transform 1 0 75256 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_818
timestamp 1644511149
transform 1 0 76360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_825
timestamp 1644511149
transform 1 0 77004 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_836
timestamp 1644511149
transform 1 0 78016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_847
timestamp 1644511149
transform 1 0 79028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_857
timestamp 1644511149
transform 1 0 79948 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_868
timestamp 1644511149
transform 1 0 80960 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_880
timestamp 1644511149
transform 1 0 82064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_890
timestamp 1644511149
transform 1 0 82984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_903
timestamp 1644511149
transform 1 0 84180 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_911
timestamp 1644511149
transform 1 0 84916 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_918
timestamp 1644511149
transform 1 0 85560 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_926
timestamp 1644511149
transform 1 0 86296 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_934
timestamp 1644511149
transform 1 0 87032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_942
timestamp 1644511149
transform 1 0 87768 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_950
timestamp 1644511149
transform 1 0 88504 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_957
timestamp 1644511149
transform 1 0 89148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_964
timestamp 1644511149
transform 1 0 89792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_972
timestamp 1644511149
transform 1 0 90528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_977
timestamp 1644511149
transform 1 0 90988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_981
timestamp 1644511149
transform 1 0 91356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_984
timestamp 1644511149
transform 1 0 91632 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_988
timestamp 1644511149
transform 1 0 92000 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_999
timestamp 1644511149
transform 1 0 93012 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1003
timestamp 1644511149
transform 1 0 93380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1007
timestamp 1644511149
transform 1 0 93748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1009
timestamp 1644511149
transform 1 0 93932 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_1017
timestamp 1644511149
transform 1 0 94668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1023
timestamp 1644511149
transform 1 0 95220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1033
timestamp 1644511149
transform 1 0 96140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1041
timestamp 1644511149
transform 1 0 96876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1047
timestamp 1644511149
transform 1 0 97428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1052
timestamp 1644511149
transform 1 0 97888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1060
timestamp 1644511149
transform 1 0 98624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1074
timestamp 1644511149
transform 1 0 99912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1082
timestamp 1644511149
transform 1 0 100648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1089
timestamp 1644511149
transform 1 0 101292 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1097
timestamp 1644511149
transform 1 0 102028 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1103
timestamp 1644511149
transform 1 0 102580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1110
timestamp 1644511149
transform 1 0 103224 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1118
timestamp 1644511149
transform 1 0 103960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1125
timestamp 1644511149
transform 1 0 104604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1130
timestamp 1644511149
transform 1 0 105064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1134
timestamp 1644511149
transform 1 0 105432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1145
timestamp 1644511149
transform 1 0 106444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1153
timestamp 1644511149
transform 1 0 107180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1157
timestamp 1644511149
transform 1 0 107548 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1161
timestamp 1644511149
transform 1 0 107916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1169
timestamp 1644511149
transform 1 0 108652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1175
timestamp 1644511149
transform 1 0 109204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1186
timestamp 1644511149
transform 1 0 110216 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1194
timestamp 1644511149
transform 1 0 110952 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1206
timestamp 1644511149
transform 1 0 112056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_1214
timestamp 1644511149
transform 1 0 112792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1225
timestamp 1644511149
transform 1 0 113804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1231
timestamp 1644511149
transform 1 0 114356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_1233
timestamp 1644511149
transform 1 0 114540 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1241
timestamp 1644511149
transform 1 0 115276 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1245
timestamp 1644511149
transform 1 0 115644 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_1256
timestamp 1644511149
transform 1 0 116656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1263
timestamp 1644511149
transform 1 0 117300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_1273
timestamp 1644511149
transform 1 0 118220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1644511149
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1644511149
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_433
timestamp 1644511149
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_445
timestamp 1644511149
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1644511149
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_489
timestamp 1644511149
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_501
timestamp 1644511149
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_513
timestamp 1644511149
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1644511149
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1644511149
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_613
timestamp 1644511149
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_625
timestamp 1644511149
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1644511149
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1644511149
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_645
timestamp 1644511149
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_657
timestamp 1644511149
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_669
timestamp 1644511149
transform 1 0 62652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_675
timestamp 1644511149
transform 1 0 63204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_687
timestamp 1644511149
transform 1 0 64308 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1644511149
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_701
timestamp 1644511149
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_713
timestamp 1644511149
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_725
timestamp 1644511149
transform 1 0 67804 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_729
timestamp 1644511149
transform 1 0 68172 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_732
timestamp 1644511149
transform 1 0 68448 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_737
timestamp 1644511149
transform 1 0 68908 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 1644511149
transform 1 0 70012 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 1644511149
transform 1 0 70564 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_757
timestamp 1644511149
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_769
timestamp 1644511149
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_781
timestamp 1644511149
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_793
timestamp 1644511149
transform 1 0 74060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 1644511149
transform 1 0 75164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 1644511149
transform 1 0 75716 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_813
timestamp 1644511149
transform 1 0 75900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_817
timestamp 1644511149
transform 1 0 76268 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_821
timestamp 1644511149
transform 1 0 76636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_833
timestamp 1644511149
transform 1 0 77740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_845
timestamp 1644511149
transform 1 0 78844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_857
timestamp 1644511149
transform 1 0 79948 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_865
timestamp 1644511149
transform 1 0 80684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_869
timestamp 1644511149
transform 1 0 81052 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_877
timestamp 1644511149
transform 1 0 81788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_883
timestamp 1644511149
transform 1 0 82340 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_895
timestamp 1644511149
transform 1 0 83444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_899
timestamp 1644511149
transform 1 0 83812 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_914
timestamp 1644511149
transform 1 0 85192 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_922
timestamp 1644511149
transform 1 0 85928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_925
timestamp 1644511149
transform 1 0 86204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_930
timestamp 1644511149
transform 1 0 86664 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_945
timestamp 1644511149
transform 1 0 88044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_957
timestamp 1644511149
transform 1 0 89148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_969
timestamp 1644511149
transform 1 0 90252 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_977
timestamp 1644511149
transform 1 0 90988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_981
timestamp 1644511149
transform 1 0 91356 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_986
timestamp 1644511149
transform 1 0 91816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_994
timestamp 1644511149
transform 1 0 92552 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1006
timestamp 1644511149
transform 1 0 93656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1018
timestamp 1644511149
transform 1 0 94760 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1030
timestamp 1644511149
transform 1 0 95864 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1040
timestamp 1644511149
transform 1 0 96784 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1056
timestamp 1644511149
transform 1 0 98256 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1060
timestamp 1644511149
transform 1 0 98624 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1067
timestamp 1644511149
transform 1 0 99268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1075
timestamp 1644511149
transform 1 0 100004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1083
timestamp 1644511149
transform 1 0 100740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1091
timestamp 1644511149
transform 1 0 101476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1093
timestamp 1644511149
transform 1 0 101660 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1105
timestamp 1644511149
transform 1 0 102764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1117
timestamp 1644511149
transform 1 0 103868 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_1129
timestamp 1644511149
transform 1 0 104972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1137
timestamp 1644511149
transform 1 0 105708 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1142
timestamp 1644511149
transform 1 0 106168 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1152
timestamp 1644511149
transform 1 0 107088 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1164
timestamp 1644511149
transform 1 0 108192 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1176
timestamp 1644511149
transform 1 0 109296 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1188
timestamp 1644511149
transform 1 0 110400 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1200
timestamp 1644511149
transform 1 0 111504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1205
timestamp 1644511149
transform 1 0 111964 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1209
timestamp 1644511149
transform 1 0 112332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_1221
timestamp 1644511149
transform 1 0 113436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_1233
timestamp 1644511149
transform 1 0 114540 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_1243
timestamp 1644511149
transform 1 0 115460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1255
timestamp 1644511149
transform 1 0 116564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1259
timestamp 1644511149
transform 1 0 116932 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_1261
timestamp 1644511149
transform 1 0 117116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_1273
timestamp 1644511149
transform 1 0 118220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_417
timestamp 1644511149
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_429
timestamp 1644511149
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1644511149
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_485
timestamp 1644511149
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1644511149
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_629
timestamp 1644511149
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_641
timestamp 1644511149
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_653
timestamp 1644511149
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1644511149
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1644511149
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_673
timestamp 1644511149
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_685
timestamp 1644511149
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_697
timestamp 1644511149
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_709
timestamp 1644511149
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1644511149
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1644511149
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_729
timestamp 1644511149
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_741
timestamp 1644511149
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_753
timestamp 1644511149
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_765
timestamp 1644511149
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1644511149
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1644511149
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_785
timestamp 1644511149
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_797
timestamp 1644511149
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_809
timestamp 1644511149
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_821
timestamp 1644511149
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1644511149
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1644511149
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_841
timestamp 1644511149
transform 1 0 78476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_853
timestamp 1644511149
transform 1 0 79580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_865
timestamp 1644511149
transform 1 0 80684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_877
timestamp 1644511149
transform 1 0 81788 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 1644511149
transform 1 0 82892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 1644511149
transform 1 0 83444 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_897
timestamp 1644511149
transform 1 0 83628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_909
timestamp 1644511149
transform 1 0 84732 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_921
timestamp 1644511149
transform 1 0 85836 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_933
timestamp 1644511149
transform 1 0 86940 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_945
timestamp 1644511149
transform 1 0 88044 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_951
timestamp 1644511149
transform 1 0 88596 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_953
timestamp 1644511149
transform 1 0 88780 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_965
timestamp 1644511149
transform 1 0 89884 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_977
timestamp 1644511149
transform 1 0 90988 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_989
timestamp 1644511149
transform 1 0 92092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1001
timestamp 1644511149
transform 1 0 93196 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1007
timestamp 1644511149
transform 1 0 93748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1009
timestamp 1644511149
transform 1 0 93932 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1021
timestamp 1644511149
transform 1 0 95036 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1033
timestamp 1644511149
transform 1 0 96140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1045
timestamp 1644511149
transform 1 0 97244 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1054
timestamp 1644511149
transform 1 0 98072 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_1062
timestamp 1644511149
transform 1 0 98808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1065
timestamp 1644511149
transform 1 0 99084 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1077
timestamp 1644511149
transform 1 0 100188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1081
timestamp 1644511149
transform 1 0 100556 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1085
timestamp 1644511149
transform 1 0 100924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1097
timestamp 1644511149
transform 1 0 102028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1109
timestamp 1644511149
transform 1 0 103132 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_1117
timestamp 1644511149
transform 1 0 103868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1121
timestamp 1644511149
transform 1 0 104236 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1133
timestamp 1644511149
transform 1 0 105340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1145
timestamp 1644511149
transform 1 0 106444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1157
timestamp 1644511149
transform 1 0 107548 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1169
timestamp 1644511149
transform 1 0 108652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1175
timestamp 1644511149
transform 1 0 109204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1177
timestamp 1644511149
transform 1 0 109388 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1189
timestamp 1644511149
transform 1 0 110492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1201
timestamp 1644511149
transform 1 0 111596 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_1213
timestamp 1644511149
transform 1 0 112700 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1225
timestamp 1644511149
transform 1 0 113804 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1231
timestamp 1644511149
transform 1 0 114356 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1233
timestamp 1644511149
transform 1 0 114540 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_1240
timestamp 1644511149
transform 1 0 115184 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1246
timestamp 1644511149
transform 1 0 115736 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1251
timestamp 1644511149
transform 1 0 116196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_1259
timestamp 1644511149
transform 1 0 116932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_1273
timestamp 1644511149
transform 1 0 118220 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_445
timestamp 1644511149
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_457
timestamp 1644511149
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1644511149
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1644511149
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_477
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_489
timestamp 1644511149
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_501
timestamp 1644511149
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_513
timestamp 1644511149
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1644511149
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1644511149
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_625
timestamp 1644511149
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1644511149
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1644511149
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_645
timestamp 1644511149
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_657
timestamp 1644511149
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_669
timestamp 1644511149
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_681
timestamp 1644511149
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1644511149
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1644511149
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_701
timestamp 1644511149
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_713
timestamp 1644511149
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_725
timestamp 1644511149
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_737
timestamp 1644511149
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1644511149
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1644511149
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_757
timestamp 1644511149
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_769
timestamp 1644511149
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_781
timestamp 1644511149
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_793
timestamp 1644511149
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1644511149
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1644511149
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_813
timestamp 1644511149
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_825
timestamp 1644511149
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_837
timestamp 1644511149
transform 1 0 78108 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_849
timestamp 1644511149
transform 1 0 79212 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_861
timestamp 1644511149
transform 1 0 80316 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_867
timestamp 1644511149
transform 1 0 80868 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_869
timestamp 1644511149
transform 1 0 81052 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_881
timestamp 1644511149
transform 1 0 82156 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_893
timestamp 1644511149
transform 1 0 83260 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_905
timestamp 1644511149
transform 1 0 84364 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_917
timestamp 1644511149
transform 1 0 85468 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_923
timestamp 1644511149
transform 1 0 86020 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_925
timestamp 1644511149
transform 1 0 86204 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_937
timestamp 1644511149
transform 1 0 87308 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_949
timestamp 1644511149
transform 1 0 88412 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_961
timestamp 1644511149
transform 1 0 89516 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_973
timestamp 1644511149
transform 1 0 90620 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_979
timestamp 1644511149
transform 1 0 91172 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_981
timestamp 1644511149
transform 1 0 91356 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_993
timestamp 1644511149
transform 1 0 92460 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1005
timestamp 1644511149
transform 1 0 93564 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1017
timestamp 1644511149
transform 1 0 94668 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1029
timestamp 1644511149
transform 1 0 95772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1035
timestamp 1644511149
transform 1 0 96324 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1037
timestamp 1644511149
transform 1 0 96508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1049
timestamp 1644511149
transform 1 0 97612 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1061
timestamp 1644511149
transform 1 0 98716 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1073
timestamp 1644511149
transform 1 0 99820 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1085
timestamp 1644511149
transform 1 0 100924 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1091
timestamp 1644511149
transform 1 0 101476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1093
timestamp 1644511149
transform 1 0 101660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1105
timestamp 1644511149
transform 1 0 102764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1117
timestamp 1644511149
transform 1 0 103868 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1129
timestamp 1644511149
transform 1 0 104972 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1141
timestamp 1644511149
transform 1 0 106076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1147
timestamp 1644511149
transform 1 0 106628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1149
timestamp 1644511149
transform 1 0 106812 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1161
timestamp 1644511149
transform 1 0 107916 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1173
timestamp 1644511149
transform 1 0 109020 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1185
timestamp 1644511149
transform 1 0 110124 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1197
timestamp 1644511149
transform 1 0 111228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1203
timestamp 1644511149
transform 1 0 111780 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1205
timestamp 1644511149
transform 1 0 111964 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1217
timestamp 1644511149
transform 1 0 113068 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_1229
timestamp 1644511149
transform 1 0 114172 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_1241
timestamp 1644511149
transform 1 0 115276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_1249
timestamp 1644511149
transform 1 0 116012 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1255
timestamp 1644511149
transform 1 0 116564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1259
timestamp 1644511149
transform 1 0 116932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_1261
timestamp 1644511149
transform 1 0 117116 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_1273
timestamp 1644511149
transform 1 0 118220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1644511149
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_585
timestamp 1644511149
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_597
timestamp 1644511149
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1644511149
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1644511149
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_629
timestamp 1644511149
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_641
timestamp 1644511149
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_653
timestamp 1644511149
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1644511149
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1644511149
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_673
timestamp 1644511149
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_685
timestamp 1644511149
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_697
timestamp 1644511149
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_709
timestamp 1644511149
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1644511149
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1644511149
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_729
timestamp 1644511149
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_741
timestamp 1644511149
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_753
timestamp 1644511149
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_765
timestamp 1644511149
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1644511149
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1644511149
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_785
timestamp 1644511149
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_797
timestamp 1644511149
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_809
timestamp 1644511149
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_821
timestamp 1644511149
transform 1 0 76636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_833
timestamp 1644511149
transform 1 0 77740 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_839
timestamp 1644511149
transform 1 0 78292 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_841
timestamp 1644511149
transform 1 0 78476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_853
timestamp 1644511149
transform 1 0 79580 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_865
timestamp 1644511149
transform 1 0 80684 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_877
timestamp 1644511149
transform 1 0 81788 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_889
timestamp 1644511149
transform 1 0 82892 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_895
timestamp 1644511149
transform 1 0 83444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_897
timestamp 1644511149
transform 1 0 83628 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_909
timestamp 1644511149
transform 1 0 84732 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_921
timestamp 1644511149
transform 1 0 85836 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_933
timestamp 1644511149
transform 1 0 86940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_945
timestamp 1644511149
transform 1 0 88044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_951
timestamp 1644511149
transform 1 0 88596 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_953
timestamp 1644511149
transform 1 0 88780 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_965
timestamp 1644511149
transform 1 0 89884 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_977
timestamp 1644511149
transform 1 0 90988 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_989
timestamp 1644511149
transform 1 0 92092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1001
timestamp 1644511149
transform 1 0 93196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1007
timestamp 1644511149
transform 1 0 93748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1009
timestamp 1644511149
transform 1 0 93932 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1021
timestamp 1644511149
transform 1 0 95036 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1033
timestamp 1644511149
transform 1 0 96140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1045
timestamp 1644511149
transform 1 0 97244 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1057
timestamp 1644511149
transform 1 0 98348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1063
timestamp 1644511149
transform 1 0 98900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1065
timestamp 1644511149
transform 1 0 99084 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1077
timestamp 1644511149
transform 1 0 100188 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1089
timestamp 1644511149
transform 1 0 101292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1101
timestamp 1644511149
transform 1 0 102396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1113
timestamp 1644511149
transform 1 0 103500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1119
timestamp 1644511149
transform 1 0 104052 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1121
timestamp 1644511149
transform 1 0 104236 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1133
timestamp 1644511149
transform 1 0 105340 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1145
timestamp 1644511149
transform 1 0 106444 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1157
timestamp 1644511149
transform 1 0 107548 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1169
timestamp 1644511149
transform 1 0 108652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1175
timestamp 1644511149
transform 1 0 109204 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1177
timestamp 1644511149
transform 1 0 109388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1189
timestamp 1644511149
transform 1 0 110492 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1201
timestamp 1644511149
transform 1 0 111596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1213
timestamp 1644511149
transform 1 0 112700 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_1225
timestamp 1644511149
transform 1 0 113804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1231
timestamp 1644511149
transform 1 0 114356 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1233
timestamp 1644511149
transform 1 0 114540 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_1245
timestamp 1644511149
transform 1 0 115644 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_1257
timestamp 1644511149
transform 1 0 116748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_1265
timestamp 1644511149
transform 1 0 117484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_1273
timestamp 1644511149
transform 1 0 118220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1644511149
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_601
timestamp 1644511149
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_613
timestamp 1644511149
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_625
timestamp 1644511149
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1644511149
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1644511149
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_645
timestamp 1644511149
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_657
timestamp 1644511149
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_669
timestamp 1644511149
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_681
timestamp 1644511149
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1644511149
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1644511149
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_701
timestamp 1644511149
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_713
timestamp 1644511149
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_725
timestamp 1644511149
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_737
timestamp 1644511149
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1644511149
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1644511149
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_757
timestamp 1644511149
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_769
timestamp 1644511149
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_781
timestamp 1644511149
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_793
timestamp 1644511149
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1644511149
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1644511149
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_813
timestamp 1644511149
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_825
timestamp 1644511149
transform 1 0 77004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_837
timestamp 1644511149
transform 1 0 78108 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_849
timestamp 1644511149
transform 1 0 79212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_861
timestamp 1644511149
transform 1 0 80316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_867
timestamp 1644511149
transform 1 0 80868 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_869
timestamp 1644511149
transform 1 0 81052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_881
timestamp 1644511149
transform 1 0 82156 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_893
timestamp 1644511149
transform 1 0 83260 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_905
timestamp 1644511149
transform 1 0 84364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_917
timestamp 1644511149
transform 1 0 85468 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_923
timestamp 1644511149
transform 1 0 86020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_925
timestamp 1644511149
transform 1 0 86204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_937
timestamp 1644511149
transform 1 0 87308 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_949
timestamp 1644511149
transform 1 0 88412 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_961
timestamp 1644511149
transform 1 0 89516 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_973
timestamp 1644511149
transform 1 0 90620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_979
timestamp 1644511149
transform 1 0 91172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_981
timestamp 1644511149
transform 1 0 91356 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_993
timestamp 1644511149
transform 1 0 92460 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1005
timestamp 1644511149
transform 1 0 93564 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1017
timestamp 1644511149
transform 1 0 94668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1029
timestamp 1644511149
transform 1 0 95772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1035
timestamp 1644511149
transform 1 0 96324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1037
timestamp 1644511149
transform 1 0 96508 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1049
timestamp 1644511149
transform 1 0 97612 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1061
timestamp 1644511149
transform 1 0 98716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1073
timestamp 1644511149
transform 1 0 99820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1085
timestamp 1644511149
transform 1 0 100924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1091
timestamp 1644511149
transform 1 0 101476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1093
timestamp 1644511149
transform 1 0 101660 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1105
timestamp 1644511149
transform 1 0 102764 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1117
timestamp 1644511149
transform 1 0 103868 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1129
timestamp 1644511149
transform 1 0 104972 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1141
timestamp 1644511149
transform 1 0 106076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1147
timestamp 1644511149
transform 1 0 106628 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1149
timestamp 1644511149
transform 1 0 106812 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1161
timestamp 1644511149
transform 1 0 107916 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1173
timestamp 1644511149
transform 1 0 109020 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1185
timestamp 1644511149
transform 1 0 110124 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1197
timestamp 1644511149
transform 1 0 111228 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1203
timestamp 1644511149
transform 1 0 111780 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1205
timestamp 1644511149
transform 1 0 111964 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1217
timestamp 1644511149
transform 1 0 113068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1229
timestamp 1644511149
transform 1 0 114172 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_1241
timestamp 1644511149
transform 1 0 115276 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1253
timestamp 1644511149
transform 1 0 116380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1259
timestamp 1644511149
transform 1 0 116932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1261
timestamp 1644511149
transform 1 0 117116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1267
timestamp 1644511149
transform 1 0 117668 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_1271
timestamp 1644511149
transform 1 0 118036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_517
timestamp 1644511149
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_529
timestamp 1644511149
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_541
timestamp 1644511149
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1644511149
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1644511149
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_573
timestamp 1644511149
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_585
timestamp 1644511149
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_597
timestamp 1644511149
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1644511149
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_617
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_629
timestamp 1644511149
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_641
timestamp 1644511149
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_653
timestamp 1644511149
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1644511149
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1644511149
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_673
timestamp 1644511149
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_685
timestamp 1644511149
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_697
timestamp 1644511149
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_709
timestamp 1644511149
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1644511149
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1644511149
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_729
timestamp 1644511149
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_741
timestamp 1644511149
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_753
timestamp 1644511149
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_765
timestamp 1644511149
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1644511149
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1644511149
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_785
timestamp 1644511149
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_797
timestamp 1644511149
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_809
timestamp 1644511149
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_821
timestamp 1644511149
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1644511149
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1644511149
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_841
timestamp 1644511149
transform 1 0 78476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_853
timestamp 1644511149
transform 1 0 79580 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_865
timestamp 1644511149
transform 1 0 80684 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_877
timestamp 1644511149
transform 1 0 81788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_889
timestamp 1644511149
transform 1 0 82892 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_895
timestamp 1644511149
transform 1 0 83444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_897
timestamp 1644511149
transform 1 0 83628 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_909
timestamp 1644511149
transform 1 0 84732 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_921
timestamp 1644511149
transform 1 0 85836 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_933
timestamp 1644511149
transform 1 0 86940 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_945
timestamp 1644511149
transform 1 0 88044 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_951
timestamp 1644511149
transform 1 0 88596 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_957
timestamp 1644511149
transform 1 0 89148 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_969
timestamp 1644511149
transform 1 0 90252 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_979
timestamp 1644511149
transform 1 0 91172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_991
timestamp 1644511149
transform 1 0 92276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1003
timestamp 1644511149
transform 1 0 93380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1007
timestamp 1644511149
transform 1 0 93748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1009
timestamp 1644511149
transform 1 0 93932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1021
timestamp 1644511149
transform 1 0 95036 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1033
timestamp 1644511149
transform 1 0 96140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1045
timestamp 1644511149
transform 1 0 97244 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1057
timestamp 1644511149
transform 1 0 98348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1063
timestamp 1644511149
transform 1 0 98900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1065
timestamp 1644511149
transform 1 0 99084 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1077
timestamp 1644511149
transform 1 0 100188 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1089
timestamp 1644511149
transform 1 0 101292 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1101
timestamp 1644511149
transform 1 0 102396 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1113
timestamp 1644511149
transform 1 0 103500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1119
timestamp 1644511149
transform 1 0 104052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1121
timestamp 1644511149
transform 1 0 104236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1133
timestamp 1644511149
transform 1 0 105340 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1145
timestamp 1644511149
transform 1 0 106444 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1157
timestamp 1644511149
transform 1 0 107548 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1169
timestamp 1644511149
transform 1 0 108652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1175
timestamp 1644511149
transform 1 0 109204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1177
timestamp 1644511149
transform 1 0 109388 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1189
timestamp 1644511149
transform 1 0 110492 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1201
timestamp 1644511149
transform 1 0 111596 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1213
timestamp 1644511149
transform 1 0 112700 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_1225
timestamp 1644511149
transform 1 0 113804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1231
timestamp 1644511149
transform 1 0 114356 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1233
timestamp 1644511149
transform 1 0 114540 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_1245
timestamp 1644511149
transform 1 0 115644 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_1257
timestamp 1644511149
transform 1 0 116748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_1265
timestamp 1644511149
transform 1 0 117484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_1273
timestamp 1644511149
transform 1 0 118220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_501
timestamp 1644511149
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1644511149
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1644511149
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_589
timestamp 1644511149
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_601
timestamp 1644511149
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_613
timestamp 1644511149
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_625
timestamp 1644511149
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1644511149
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1644511149
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_645
timestamp 1644511149
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_657
timestamp 1644511149
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_669
timestamp 1644511149
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_681
timestamp 1644511149
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1644511149
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1644511149
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_701
timestamp 1644511149
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_713
timestamp 1644511149
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_725
timestamp 1644511149
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_737
timestamp 1644511149
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1644511149
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1644511149
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_757
timestamp 1644511149
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_769
timestamp 1644511149
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_781
timestamp 1644511149
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_793
timestamp 1644511149
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1644511149
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1644511149
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_813
timestamp 1644511149
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_825
timestamp 1644511149
transform 1 0 77004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_837
timestamp 1644511149
transform 1 0 78108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_849
timestamp 1644511149
transform 1 0 79212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_861
timestamp 1644511149
transform 1 0 80316 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_867
timestamp 1644511149
transform 1 0 80868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_869
timestamp 1644511149
transform 1 0 81052 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_881
timestamp 1644511149
transform 1 0 82156 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_893
timestamp 1644511149
transform 1 0 83260 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_905
timestamp 1644511149
transform 1 0 84364 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_917
timestamp 1644511149
transform 1 0 85468 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_923
timestamp 1644511149
transform 1 0 86020 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_925
timestamp 1644511149
transform 1 0 86204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_937
timestamp 1644511149
transform 1 0 87308 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_949
timestamp 1644511149
transform 1 0 88412 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_961
timestamp 1644511149
transform 1 0 89516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_973
timestamp 1644511149
transform 1 0 90620 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_979
timestamp 1644511149
transform 1 0 91172 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_981
timestamp 1644511149
transform 1 0 91356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_993
timestamp 1644511149
transform 1 0 92460 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1005
timestamp 1644511149
transform 1 0 93564 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1017
timestamp 1644511149
transform 1 0 94668 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1029
timestamp 1644511149
transform 1 0 95772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1035
timestamp 1644511149
transform 1 0 96324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1037
timestamp 1644511149
transform 1 0 96508 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1049
timestamp 1644511149
transform 1 0 97612 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1061
timestamp 1644511149
transform 1 0 98716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1073
timestamp 1644511149
transform 1 0 99820 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1085
timestamp 1644511149
transform 1 0 100924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1091
timestamp 1644511149
transform 1 0 101476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1093
timestamp 1644511149
transform 1 0 101660 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1105
timestamp 1644511149
transform 1 0 102764 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1117
timestamp 1644511149
transform 1 0 103868 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1129
timestamp 1644511149
transform 1 0 104972 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1141
timestamp 1644511149
transform 1 0 106076 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1147
timestamp 1644511149
transform 1 0 106628 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1149
timestamp 1644511149
transform 1 0 106812 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1161
timestamp 1644511149
transform 1 0 107916 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1173
timestamp 1644511149
transform 1 0 109020 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1185
timestamp 1644511149
transform 1 0 110124 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1197
timestamp 1644511149
transform 1 0 111228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1203
timestamp 1644511149
transform 1 0 111780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1205
timestamp 1644511149
transform 1 0 111964 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1217
timestamp 1644511149
transform 1 0 113068 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1229
timestamp 1644511149
transform 1 0 114172 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1241
timestamp 1644511149
transform 1 0 115276 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_1253
timestamp 1644511149
transform 1 0 116380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1259
timestamp 1644511149
transform 1 0 116932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_1261
timestamp 1644511149
transform 1 0 117116 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_1273
timestamp 1644511149
transform 1 0 118220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1644511149
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1644511149
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1644511149
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1644511149
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_597
timestamp 1644511149
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1644511149
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1644511149
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_629
timestamp 1644511149
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_641
timestamp 1644511149
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_653
timestamp 1644511149
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1644511149
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1644511149
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_673
timestamp 1644511149
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_685
timestamp 1644511149
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_697
timestamp 1644511149
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_709
timestamp 1644511149
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1644511149
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1644511149
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_729
timestamp 1644511149
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_741
timestamp 1644511149
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_753
timestamp 1644511149
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_765
timestamp 1644511149
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1644511149
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1644511149
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_785
timestamp 1644511149
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_797
timestamp 1644511149
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_809
timestamp 1644511149
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_821
timestamp 1644511149
transform 1 0 76636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_833
timestamp 1644511149
transform 1 0 77740 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_839
timestamp 1644511149
transform 1 0 78292 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_841
timestamp 1644511149
transform 1 0 78476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_853
timestamp 1644511149
transform 1 0 79580 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_865
timestamp 1644511149
transform 1 0 80684 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_877
timestamp 1644511149
transform 1 0 81788 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_889
timestamp 1644511149
transform 1 0 82892 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_895
timestamp 1644511149
transform 1 0 83444 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_897
timestamp 1644511149
transform 1 0 83628 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_909
timestamp 1644511149
transform 1 0 84732 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_921
timestamp 1644511149
transform 1 0 85836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_933
timestamp 1644511149
transform 1 0 86940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_945
timestamp 1644511149
transform 1 0 88044 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_951
timestamp 1644511149
transform 1 0 88596 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_953
timestamp 1644511149
transform 1 0 88780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_965
timestamp 1644511149
transform 1 0 89884 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_977
timestamp 1644511149
transform 1 0 90988 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_989
timestamp 1644511149
transform 1 0 92092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1001
timestamp 1644511149
transform 1 0 93196 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1007
timestamp 1644511149
transform 1 0 93748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1009
timestamp 1644511149
transform 1 0 93932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1021
timestamp 1644511149
transform 1 0 95036 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1033
timestamp 1644511149
transform 1 0 96140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1045
timestamp 1644511149
transform 1 0 97244 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1057
timestamp 1644511149
transform 1 0 98348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1063
timestamp 1644511149
transform 1 0 98900 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1065
timestamp 1644511149
transform 1 0 99084 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1077
timestamp 1644511149
transform 1 0 100188 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1089
timestamp 1644511149
transform 1 0 101292 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1101
timestamp 1644511149
transform 1 0 102396 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1113
timestamp 1644511149
transform 1 0 103500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1119
timestamp 1644511149
transform 1 0 104052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1121
timestamp 1644511149
transform 1 0 104236 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1133
timestamp 1644511149
transform 1 0 105340 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1145
timestamp 1644511149
transform 1 0 106444 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1157
timestamp 1644511149
transform 1 0 107548 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1169
timestamp 1644511149
transform 1 0 108652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1175
timestamp 1644511149
transform 1 0 109204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1177
timestamp 1644511149
transform 1 0 109388 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1189
timestamp 1644511149
transform 1 0 110492 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1201
timestamp 1644511149
transform 1 0 111596 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1213
timestamp 1644511149
transform 1 0 112700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_1225
timestamp 1644511149
transform 1 0 113804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1231
timestamp 1644511149
transform 1 0 114356 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1233
timestamp 1644511149
transform 1 0 114540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_1245
timestamp 1644511149
transform 1 0 115644 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_1257
timestamp 1644511149
transform 1 0 116748 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_1265
timestamp 1644511149
transform 1 0 117484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_1273
timestamp 1644511149
transform 1 0 118220 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1644511149
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1644511149
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_557
timestamp 1644511149
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_569
timestamp 1644511149
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1644511149
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_613
timestamp 1644511149
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_625
timestamp 1644511149
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1644511149
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1644511149
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_645
timestamp 1644511149
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_657
timestamp 1644511149
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_669
timestamp 1644511149
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_681
timestamp 1644511149
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1644511149
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1644511149
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_701
timestamp 1644511149
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_713
timestamp 1644511149
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_725
timestamp 1644511149
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_737
timestamp 1644511149
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1644511149
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1644511149
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_757
timestamp 1644511149
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_769
timestamp 1644511149
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_781
timestamp 1644511149
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_793
timestamp 1644511149
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1644511149
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1644511149
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_813
timestamp 1644511149
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_825
timestamp 1644511149
transform 1 0 77004 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_837
timestamp 1644511149
transform 1 0 78108 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_849
timestamp 1644511149
transform 1 0 79212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_861
timestamp 1644511149
transform 1 0 80316 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_867
timestamp 1644511149
transform 1 0 80868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_869
timestamp 1644511149
transform 1 0 81052 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_881
timestamp 1644511149
transform 1 0 82156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_893
timestamp 1644511149
transform 1 0 83260 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_905
timestamp 1644511149
transform 1 0 84364 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_917
timestamp 1644511149
transform 1 0 85468 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_923
timestamp 1644511149
transform 1 0 86020 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_925
timestamp 1644511149
transform 1 0 86204 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_937
timestamp 1644511149
transform 1 0 87308 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_949
timestamp 1644511149
transform 1 0 88412 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_961
timestamp 1644511149
transform 1 0 89516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_973
timestamp 1644511149
transform 1 0 90620 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_979
timestamp 1644511149
transform 1 0 91172 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_981
timestamp 1644511149
transform 1 0 91356 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_993
timestamp 1644511149
transform 1 0 92460 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1005
timestamp 1644511149
transform 1 0 93564 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1017
timestamp 1644511149
transform 1 0 94668 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1029
timestamp 1644511149
transform 1 0 95772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1035
timestamp 1644511149
transform 1 0 96324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1037
timestamp 1644511149
transform 1 0 96508 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1049
timestamp 1644511149
transform 1 0 97612 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1061
timestamp 1644511149
transform 1 0 98716 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1073
timestamp 1644511149
transform 1 0 99820 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1085
timestamp 1644511149
transform 1 0 100924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1091
timestamp 1644511149
transform 1 0 101476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1093
timestamp 1644511149
transform 1 0 101660 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1105
timestamp 1644511149
transform 1 0 102764 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1117
timestamp 1644511149
transform 1 0 103868 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1129
timestamp 1644511149
transform 1 0 104972 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1141
timestamp 1644511149
transform 1 0 106076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1147
timestamp 1644511149
transform 1 0 106628 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1149
timestamp 1644511149
transform 1 0 106812 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1161
timestamp 1644511149
transform 1 0 107916 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1173
timestamp 1644511149
transform 1 0 109020 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1185
timestamp 1644511149
transform 1 0 110124 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1197
timestamp 1644511149
transform 1 0 111228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1203
timestamp 1644511149
transform 1 0 111780 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1205
timestamp 1644511149
transform 1 0 111964 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1217
timestamp 1644511149
transform 1 0 113068 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1229
timestamp 1644511149
transform 1 0 114172 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_1241
timestamp 1644511149
transform 1 0 115276 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1253
timestamp 1644511149
transform 1 0 116380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1259
timestamp 1644511149
transform 1 0 116932 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_1261
timestamp 1644511149
transform 1 0 117116 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_1273
timestamp 1644511149
transform 1 0 118220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_517
timestamp 1644511149
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_529
timestamp 1644511149
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_541
timestamp 1644511149
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1644511149
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1644511149
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_561
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_573
timestamp 1644511149
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1644511149
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1644511149
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_629
timestamp 1644511149
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_641
timestamp 1644511149
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_653
timestamp 1644511149
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1644511149
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1644511149
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_673
timestamp 1644511149
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_685
timestamp 1644511149
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_697
timestamp 1644511149
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_709
timestamp 1644511149
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1644511149
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1644511149
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_729
timestamp 1644511149
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_741
timestamp 1644511149
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_753
timestamp 1644511149
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_765
timestamp 1644511149
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1644511149
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1644511149
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_785
timestamp 1644511149
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_797
timestamp 1644511149
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_809
timestamp 1644511149
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_821
timestamp 1644511149
transform 1 0 76636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_833
timestamp 1644511149
transform 1 0 77740 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_839
timestamp 1644511149
transform 1 0 78292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_841
timestamp 1644511149
transform 1 0 78476 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_853
timestamp 1644511149
transform 1 0 79580 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_865
timestamp 1644511149
transform 1 0 80684 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_877
timestamp 1644511149
transform 1 0 81788 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_889
timestamp 1644511149
transform 1 0 82892 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_895
timestamp 1644511149
transform 1 0 83444 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_897
timestamp 1644511149
transform 1 0 83628 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_909
timestamp 1644511149
transform 1 0 84732 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_921
timestamp 1644511149
transform 1 0 85836 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_933
timestamp 1644511149
transform 1 0 86940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_945
timestamp 1644511149
transform 1 0 88044 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_951
timestamp 1644511149
transform 1 0 88596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_953
timestamp 1644511149
transform 1 0 88780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_965
timestamp 1644511149
transform 1 0 89884 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_977
timestamp 1644511149
transform 1 0 90988 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_989
timestamp 1644511149
transform 1 0 92092 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1001
timestamp 1644511149
transform 1 0 93196 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1007
timestamp 1644511149
transform 1 0 93748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1009
timestamp 1644511149
transform 1 0 93932 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1021
timestamp 1644511149
transform 1 0 95036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1033
timestamp 1644511149
transform 1 0 96140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1045
timestamp 1644511149
transform 1 0 97244 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1057
timestamp 1644511149
transform 1 0 98348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1063
timestamp 1644511149
transform 1 0 98900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1065
timestamp 1644511149
transform 1 0 99084 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1077
timestamp 1644511149
transform 1 0 100188 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1089
timestamp 1644511149
transform 1 0 101292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1101
timestamp 1644511149
transform 1 0 102396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1113
timestamp 1644511149
transform 1 0 103500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1119
timestamp 1644511149
transform 1 0 104052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1121
timestamp 1644511149
transform 1 0 104236 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1133
timestamp 1644511149
transform 1 0 105340 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1145
timestamp 1644511149
transform 1 0 106444 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1157
timestamp 1644511149
transform 1 0 107548 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1169
timestamp 1644511149
transform 1 0 108652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1175
timestamp 1644511149
transform 1 0 109204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1177
timestamp 1644511149
transform 1 0 109388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1189
timestamp 1644511149
transform 1 0 110492 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1201
timestamp 1644511149
transform 1 0 111596 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1213
timestamp 1644511149
transform 1 0 112700 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_1225
timestamp 1644511149
transform 1 0 113804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1231
timestamp 1644511149
transform 1 0 114356 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1233
timestamp 1644511149
transform 1 0 114540 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1245
timestamp 1644511149
transform 1 0 115644 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_1257
timestamp 1644511149
transform 1 0 116748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_1269
timestamp 1644511149
transform 1 0 117852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_513
timestamp 1644511149
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1644511149
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1644511149
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_557
timestamp 1644511149
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_569
timestamp 1644511149
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_601
timestamp 1644511149
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_613
timestamp 1644511149
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_625
timestamp 1644511149
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1644511149
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1644511149
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_645
timestamp 1644511149
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_657
timestamp 1644511149
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_669
timestamp 1644511149
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_681
timestamp 1644511149
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1644511149
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1644511149
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_701
timestamp 1644511149
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_713
timestamp 1644511149
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_725
timestamp 1644511149
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_737
timestamp 1644511149
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1644511149
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1644511149
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_757
timestamp 1644511149
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_769
timestamp 1644511149
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_781
timestamp 1644511149
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_793
timestamp 1644511149
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1644511149
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1644511149
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_813
timestamp 1644511149
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_825
timestamp 1644511149
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_837
timestamp 1644511149
transform 1 0 78108 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_849
timestamp 1644511149
transform 1 0 79212 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_861
timestamp 1644511149
transform 1 0 80316 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_867
timestamp 1644511149
transform 1 0 80868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_869
timestamp 1644511149
transform 1 0 81052 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_881
timestamp 1644511149
transform 1 0 82156 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_893
timestamp 1644511149
transform 1 0 83260 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_905
timestamp 1644511149
transform 1 0 84364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_917
timestamp 1644511149
transform 1 0 85468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_923
timestamp 1644511149
transform 1 0 86020 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_925
timestamp 1644511149
transform 1 0 86204 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_937
timestamp 1644511149
transform 1 0 87308 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_949
timestamp 1644511149
transform 1 0 88412 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_961
timestamp 1644511149
transform 1 0 89516 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_973
timestamp 1644511149
transform 1 0 90620 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_979
timestamp 1644511149
transform 1 0 91172 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_981
timestamp 1644511149
transform 1 0 91356 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_993
timestamp 1644511149
transform 1 0 92460 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1005
timestamp 1644511149
transform 1 0 93564 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1017
timestamp 1644511149
transform 1 0 94668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1029
timestamp 1644511149
transform 1 0 95772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1035
timestamp 1644511149
transform 1 0 96324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1037
timestamp 1644511149
transform 1 0 96508 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1049
timestamp 1644511149
transform 1 0 97612 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1061
timestamp 1644511149
transform 1 0 98716 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1073
timestamp 1644511149
transform 1 0 99820 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1085
timestamp 1644511149
transform 1 0 100924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1091
timestamp 1644511149
transform 1 0 101476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1093
timestamp 1644511149
transform 1 0 101660 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1105
timestamp 1644511149
transform 1 0 102764 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1117
timestamp 1644511149
transform 1 0 103868 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1129
timestamp 1644511149
transform 1 0 104972 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1141
timestamp 1644511149
transform 1 0 106076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1147
timestamp 1644511149
transform 1 0 106628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1149
timestamp 1644511149
transform 1 0 106812 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1161
timestamp 1644511149
transform 1 0 107916 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1173
timestamp 1644511149
transform 1 0 109020 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1185
timestamp 1644511149
transform 1 0 110124 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1197
timestamp 1644511149
transform 1 0 111228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1203
timestamp 1644511149
transform 1 0 111780 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1205
timestamp 1644511149
transform 1 0 111964 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1217
timestamp 1644511149
transform 1 0 113068 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1229
timestamp 1644511149
transform 1 0 114172 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_1241
timestamp 1644511149
transform 1 0 115276 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1253
timestamp 1644511149
transform 1 0 116380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1259
timestamp 1644511149
transform 1 0 116932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_1261
timestamp 1644511149
transform 1 0 117116 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_1273
timestamp 1644511149
transform 1 0 118220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_585
timestamp 1644511149
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_597
timestamp 1644511149
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1644511149
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1644511149
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_629
timestamp 1644511149
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_641
timestamp 1644511149
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_653
timestamp 1644511149
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1644511149
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1644511149
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_673
timestamp 1644511149
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_685
timestamp 1644511149
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_697
timestamp 1644511149
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_709
timestamp 1644511149
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1644511149
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1644511149
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_729
timestamp 1644511149
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_741
timestamp 1644511149
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_753
timestamp 1644511149
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_765
timestamp 1644511149
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1644511149
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1644511149
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_785
timestamp 1644511149
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_797
timestamp 1644511149
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_809
timestamp 1644511149
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_821
timestamp 1644511149
transform 1 0 76636 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_833
timestamp 1644511149
transform 1 0 77740 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_839
timestamp 1644511149
transform 1 0 78292 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_841
timestamp 1644511149
transform 1 0 78476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_853
timestamp 1644511149
transform 1 0 79580 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_865
timestamp 1644511149
transform 1 0 80684 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_877
timestamp 1644511149
transform 1 0 81788 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_889
timestamp 1644511149
transform 1 0 82892 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_895
timestamp 1644511149
transform 1 0 83444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_897
timestamp 1644511149
transform 1 0 83628 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_909
timestamp 1644511149
transform 1 0 84732 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_921
timestamp 1644511149
transform 1 0 85836 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_933
timestamp 1644511149
transform 1 0 86940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_945
timestamp 1644511149
transform 1 0 88044 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_951
timestamp 1644511149
transform 1 0 88596 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_953
timestamp 1644511149
transform 1 0 88780 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_965
timestamp 1644511149
transform 1 0 89884 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_977
timestamp 1644511149
transform 1 0 90988 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_989
timestamp 1644511149
transform 1 0 92092 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1001
timestamp 1644511149
transform 1 0 93196 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1007
timestamp 1644511149
transform 1 0 93748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1009
timestamp 1644511149
transform 1 0 93932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1021
timestamp 1644511149
transform 1 0 95036 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1033
timestamp 1644511149
transform 1 0 96140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1045
timestamp 1644511149
transform 1 0 97244 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1057
timestamp 1644511149
transform 1 0 98348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1063
timestamp 1644511149
transform 1 0 98900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1065
timestamp 1644511149
transform 1 0 99084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1077
timestamp 1644511149
transform 1 0 100188 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1089
timestamp 1644511149
transform 1 0 101292 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1101
timestamp 1644511149
transform 1 0 102396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1113
timestamp 1644511149
transform 1 0 103500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1119
timestamp 1644511149
transform 1 0 104052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1121
timestamp 1644511149
transform 1 0 104236 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1133
timestamp 1644511149
transform 1 0 105340 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1145
timestamp 1644511149
transform 1 0 106444 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1157
timestamp 1644511149
transform 1 0 107548 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1169
timestamp 1644511149
transform 1 0 108652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1175
timestamp 1644511149
transform 1 0 109204 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1177
timestamp 1644511149
transform 1 0 109388 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1189
timestamp 1644511149
transform 1 0 110492 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1201
timestamp 1644511149
transform 1 0 111596 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1213
timestamp 1644511149
transform 1 0 112700 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_1225
timestamp 1644511149
transform 1 0 113804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1231
timestamp 1644511149
transform 1 0 114356 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1233
timestamp 1644511149
transform 1 0 114540 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1245
timestamp 1644511149
transform 1 0 115644 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_1257
timestamp 1644511149
transform 1 0 116748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_1269
timestamp 1644511149
transform 1 0 117852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1644511149
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_545
timestamp 1644511149
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_557
timestamp 1644511149
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_569
timestamp 1644511149
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1644511149
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_601
timestamp 1644511149
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_613
timestamp 1644511149
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_625
timestamp 1644511149
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1644511149
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1644511149
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_645
timestamp 1644511149
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_657
timestamp 1644511149
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_669
timestamp 1644511149
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_681
timestamp 1644511149
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1644511149
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1644511149
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_701
timestamp 1644511149
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_713
timestamp 1644511149
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_725
timestamp 1644511149
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_737
timestamp 1644511149
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1644511149
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1644511149
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_757
timestamp 1644511149
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_769
timestamp 1644511149
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_781
timestamp 1644511149
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_793
timestamp 1644511149
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1644511149
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1644511149
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_817
timestamp 1644511149
transform 1 0 76268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_829
timestamp 1644511149
transform 1 0 77372 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_841
timestamp 1644511149
transform 1 0 78476 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_853
timestamp 1644511149
transform 1 0 79580 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_865
timestamp 1644511149
transform 1 0 80684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_869
timestamp 1644511149
transform 1 0 81052 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_881
timestamp 1644511149
transform 1 0 82156 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_893
timestamp 1644511149
transform 1 0 83260 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_905
timestamp 1644511149
transform 1 0 84364 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_917
timestamp 1644511149
transform 1 0 85468 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_923
timestamp 1644511149
transform 1 0 86020 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_925
timestamp 1644511149
transform 1 0 86204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_937
timestamp 1644511149
transform 1 0 87308 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_949
timestamp 1644511149
transform 1 0 88412 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_961
timestamp 1644511149
transform 1 0 89516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_973
timestamp 1644511149
transform 1 0 90620 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_979
timestamp 1644511149
transform 1 0 91172 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_981
timestamp 1644511149
transform 1 0 91356 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_993
timestamp 1644511149
transform 1 0 92460 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1005
timestamp 1644511149
transform 1 0 93564 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1017
timestamp 1644511149
transform 1 0 94668 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1029
timestamp 1644511149
transform 1 0 95772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1035
timestamp 1644511149
transform 1 0 96324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1037
timestamp 1644511149
transform 1 0 96508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1049
timestamp 1644511149
transform 1 0 97612 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1061
timestamp 1644511149
transform 1 0 98716 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1073
timestamp 1644511149
transform 1 0 99820 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1085
timestamp 1644511149
transform 1 0 100924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1091
timestamp 1644511149
transform 1 0 101476 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1093
timestamp 1644511149
transform 1 0 101660 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1105
timestamp 1644511149
transform 1 0 102764 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1117
timestamp 1644511149
transform 1 0 103868 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1129
timestamp 1644511149
transform 1 0 104972 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1141
timestamp 1644511149
transform 1 0 106076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1147
timestamp 1644511149
transform 1 0 106628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1149
timestamp 1644511149
transform 1 0 106812 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1161
timestamp 1644511149
transform 1 0 107916 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1173
timestamp 1644511149
transform 1 0 109020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1185
timestamp 1644511149
transform 1 0 110124 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1197
timestamp 1644511149
transform 1 0 111228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1203
timestamp 1644511149
transform 1 0 111780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1205
timestamp 1644511149
transform 1 0 111964 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1217
timestamp 1644511149
transform 1 0 113068 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1229
timestamp 1644511149
transform 1 0 114172 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_1241
timestamp 1644511149
transform 1 0 115276 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1253
timestamp 1644511149
transform 1 0 116380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1259
timestamp 1644511149
transform 1 0 116932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_1261
timestamp 1644511149
transform 1 0 117116 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_1273
timestamp 1644511149
transform 1 0 118220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_517
timestamp 1644511149
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_529
timestamp 1644511149
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_541
timestamp 1644511149
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1644511149
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1644511149
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_561
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_573
timestamp 1644511149
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_585
timestamp 1644511149
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_597
timestamp 1644511149
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1644511149
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1644511149
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_617
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_629
timestamp 1644511149
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_641
timestamp 1644511149
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_653
timestamp 1644511149
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1644511149
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1644511149
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_673
timestamp 1644511149
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_685
timestamp 1644511149
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_697
timestamp 1644511149
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_709
timestamp 1644511149
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1644511149
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1644511149
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_729
timestamp 1644511149
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_741
timestamp 1644511149
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_753
timestamp 1644511149
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_765
timestamp 1644511149
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1644511149
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1644511149
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_785
timestamp 1644511149
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_797
timestamp 1644511149
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_809
timestamp 1644511149
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_821
timestamp 1644511149
transform 1 0 76636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_833
timestamp 1644511149
transform 1 0 77740 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_839
timestamp 1644511149
transform 1 0 78292 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_841
timestamp 1644511149
transform 1 0 78476 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_853
timestamp 1644511149
transform 1 0 79580 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_865
timestamp 1644511149
transform 1 0 80684 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_877
timestamp 1644511149
transform 1 0 81788 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_889
timestamp 1644511149
transform 1 0 82892 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_895
timestamp 1644511149
transform 1 0 83444 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_897
timestamp 1644511149
transform 1 0 83628 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_909
timestamp 1644511149
transform 1 0 84732 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_921
timestamp 1644511149
transform 1 0 85836 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_933
timestamp 1644511149
transform 1 0 86940 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_945
timestamp 1644511149
transform 1 0 88044 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_951
timestamp 1644511149
transform 1 0 88596 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_953
timestamp 1644511149
transform 1 0 88780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_965
timestamp 1644511149
transform 1 0 89884 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_977
timestamp 1644511149
transform 1 0 90988 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_989
timestamp 1644511149
transform 1 0 92092 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1001
timestamp 1644511149
transform 1 0 93196 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1007
timestamp 1644511149
transform 1 0 93748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1009
timestamp 1644511149
transform 1 0 93932 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1021
timestamp 1644511149
transform 1 0 95036 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1033
timestamp 1644511149
transform 1 0 96140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1045
timestamp 1644511149
transform 1 0 97244 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1057
timestamp 1644511149
transform 1 0 98348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1063
timestamp 1644511149
transform 1 0 98900 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1065
timestamp 1644511149
transform 1 0 99084 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1077
timestamp 1644511149
transform 1 0 100188 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1089
timestamp 1644511149
transform 1 0 101292 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1101
timestamp 1644511149
transform 1 0 102396 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1113
timestamp 1644511149
transform 1 0 103500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1119
timestamp 1644511149
transform 1 0 104052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1121
timestamp 1644511149
transform 1 0 104236 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1133
timestamp 1644511149
transform 1 0 105340 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1145
timestamp 1644511149
transform 1 0 106444 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1157
timestamp 1644511149
transform 1 0 107548 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1169
timestamp 1644511149
transform 1 0 108652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1175
timestamp 1644511149
transform 1 0 109204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1177
timestamp 1644511149
transform 1 0 109388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1189
timestamp 1644511149
transform 1 0 110492 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1201
timestamp 1644511149
transform 1 0 111596 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1213
timestamp 1644511149
transform 1 0 112700 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_1225
timestamp 1644511149
transform 1 0 113804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1231
timestamp 1644511149
transform 1 0 114356 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1233
timestamp 1644511149
transform 1 0 114540 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1245
timestamp 1644511149
transform 1 0 115644 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_1257
timestamp 1644511149
transform 1 0 116748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_1269
timestamp 1644511149
transform 1 0 117852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_501
timestamp 1644511149
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_513
timestamp 1644511149
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_557
timestamp 1644511149
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_569
timestamp 1644511149
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1644511149
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1644511149
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_601
timestamp 1644511149
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_613
timestamp 1644511149
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_625
timestamp 1644511149
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1644511149
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1644511149
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_645
timestamp 1644511149
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_657
timestamp 1644511149
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_669
timestamp 1644511149
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_681
timestamp 1644511149
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1644511149
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1644511149
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_701
timestamp 1644511149
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_713
timestamp 1644511149
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_725
timestamp 1644511149
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_737
timestamp 1644511149
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1644511149
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1644511149
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_757
timestamp 1644511149
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_769
timestamp 1644511149
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_781
timestamp 1644511149
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_793
timestamp 1644511149
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1644511149
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1644511149
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_813
timestamp 1644511149
transform 1 0 75900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_825
timestamp 1644511149
transform 1 0 77004 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_837
timestamp 1644511149
transform 1 0 78108 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_849
timestamp 1644511149
transform 1 0 79212 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_861
timestamp 1644511149
transform 1 0 80316 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_867
timestamp 1644511149
transform 1 0 80868 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_869
timestamp 1644511149
transform 1 0 81052 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_881
timestamp 1644511149
transform 1 0 82156 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_893
timestamp 1644511149
transform 1 0 83260 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_905
timestamp 1644511149
transform 1 0 84364 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_917
timestamp 1644511149
transform 1 0 85468 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_923
timestamp 1644511149
transform 1 0 86020 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_925
timestamp 1644511149
transform 1 0 86204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_937
timestamp 1644511149
transform 1 0 87308 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_949
timestamp 1644511149
transform 1 0 88412 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_961
timestamp 1644511149
transform 1 0 89516 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_973
timestamp 1644511149
transform 1 0 90620 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_979
timestamp 1644511149
transform 1 0 91172 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_981
timestamp 1644511149
transform 1 0 91356 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_993
timestamp 1644511149
transform 1 0 92460 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1005
timestamp 1644511149
transform 1 0 93564 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1017
timestamp 1644511149
transform 1 0 94668 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1029
timestamp 1644511149
transform 1 0 95772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1035
timestamp 1644511149
transform 1 0 96324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1037
timestamp 1644511149
transform 1 0 96508 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1049
timestamp 1644511149
transform 1 0 97612 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1061
timestamp 1644511149
transform 1 0 98716 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1073
timestamp 1644511149
transform 1 0 99820 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1085
timestamp 1644511149
transform 1 0 100924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1091
timestamp 1644511149
transform 1 0 101476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1093
timestamp 1644511149
transform 1 0 101660 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1105
timestamp 1644511149
transform 1 0 102764 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1117
timestamp 1644511149
transform 1 0 103868 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1129
timestamp 1644511149
transform 1 0 104972 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1141
timestamp 1644511149
transform 1 0 106076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1147
timestamp 1644511149
transform 1 0 106628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1149
timestamp 1644511149
transform 1 0 106812 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1161
timestamp 1644511149
transform 1 0 107916 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1173
timestamp 1644511149
transform 1 0 109020 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1185
timestamp 1644511149
transform 1 0 110124 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1197
timestamp 1644511149
transform 1 0 111228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1203
timestamp 1644511149
transform 1 0 111780 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1205
timestamp 1644511149
transform 1 0 111964 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1217
timestamp 1644511149
transform 1 0 113068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1229
timestamp 1644511149
transform 1 0 114172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_1241
timestamp 1644511149
transform 1 0 115276 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_1253
timestamp 1644511149
transform 1 0 116380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1259
timestamp 1644511149
transform 1 0 116932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1261
timestamp 1644511149
transform 1 0 117116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_1267
timestamp 1644511149
transform 1 0 117668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_1273
timestamp 1644511149
transform 1 0 118220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_517
timestamp 1644511149
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_529
timestamp 1644511149
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_541
timestamp 1644511149
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1644511149
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1644511149
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_573
timestamp 1644511149
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_585
timestamp 1644511149
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_597
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1644511149
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_629
timestamp 1644511149
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_641
timestamp 1644511149
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_653
timestamp 1644511149
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1644511149
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1644511149
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_673
timestamp 1644511149
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_685
timestamp 1644511149
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_697
timestamp 1644511149
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_709
timestamp 1644511149
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1644511149
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1644511149
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_729
timestamp 1644511149
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_741
timestamp 1644511149
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_753
timestamp 1644511149
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_765
timestamp 1644511149
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1644511149
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1644511149
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_785
timestamp 1644511149
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_797
timestamp 1644511149
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_809
timestamp 1644511149
transform 1 0 75532 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_821
timestamp 1644511149
transform 1 0 76636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_833
timestamp 1644511149
transform 1 0 77740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_839
timestamp 1644511149
transform 1 0 78292 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_841
timestamp 1644511149
transform 1 0 78476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_853
timestamp 1644511149
transform 1 0 79580 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_865
timestamp 1644511149
transform 1 0 80684 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_877
timestamp 1644511149
transform 1 0 81788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_889
timestamp 1644511149
transform 1 0 82892 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_895
timestamp 1644511149
transform 1 0 83444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_897
timestamp 1644511149
transform 1 0 83628 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_909
timestamp 1644511149
transform 1 0 84732 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_921
timestamp 1644511149
transform 1 0 85836 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_933
timestamp 1644511149
transform 1 0 86940 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_945
timestamp 1644511149
transform 1 0 88044 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_951
timestamp 1644511149
transform 1 0 88596 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_953
timestamp 1644511149
transform 1 0 88780 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_965
timestamp 1644511149
transform 1 0 89884 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_977
timestamp 1644511149
transform 1 0 90988 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_989
timestamp 1644511149
transform 1 0 92092 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1001
timestamp 1644511149
transform 1 0 93196 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1007
timestamp 1644511149
transform 1 0 93748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1009
timestamp 1644511149
transform 1 0 93932 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1021
timestamp 1644511149
transform 1 0 95036 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1033
timestamp 1644511149
transform 1 0 96140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1045
timestamp 1644511149
transform 1 0 97244 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1057
timestamp 1644511149
transform 1 0 98348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1063
timestamp 1644511149
transform 1 0 98900 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1065
timestamp 1644511149
transform 1 0 99084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1077
timestamp 1644511149
transform 1 0 100188 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1089
timestamp 1644511149
transform 1 0 101292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1101
timestamp 1644511149
transform 1 0 102396 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1113
timestamp 1644511149
transform 1 0 103500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1119
timestamp 1644511149
transform 1 0 104052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1121
timestamp 1644511149
transform 1 0 104236 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1133
timestamp 1644511149
transform 1 0 105340 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1145
timestamp 1644511149
transform 1 0 106444 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1157
timestamp 1644511149
transform 1 0 107548 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1169
timestamp 1644511149
transform 1 0 108652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1175
timestamp 1644511149
transform 1 0 109204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1177
timestamp 1644511149
transform 1 0 109388 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1189
timestamp 1644511149
transform 1 0 110492 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1201
timestamp 1644511149
transform 1 0 111596 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1213
timestamp 1644511149
transform 1 0 112700 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_1225
timestamp 1644511149
transform 1 0 113804 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1231
timestamp 1644511149
transform 1 0 114356 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1233
timestamp 1644511149
transform 1 0 114540 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_1245
timestamp 1644511149
transform 1 0 115644 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_1257
timestamp 1644511149
transform 1 0 116748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_1267
timestamp 1644511149
transform 1 0 117668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_1273
timestamp 1644511149
transform 1 0 118220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1644511149
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1644511149
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_545
timestamp 1644511149
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_601
timestamp 1644511149
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_613
timestamp 1644511149
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_625
timestamp 1644511149
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1644511149
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1644511149
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_645
timestamp 1644511149
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_657
timestamp 1644511149
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_669
timestamp 1644511149
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_681
timestamp 1644511149
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1644511149
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1644511149
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_701
timestamp 1644511149
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_713
timestamp 1644511149
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_725
timestamp 1644511149
transform 1 0 67804 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_737
timestamp 1644511149
transform 1 0 68908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1644511149
transform 1 0 70012 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1644511149
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_757
timestamp 1644511149
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_769
timestamp 1644511149
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_781
timestamp 1644511149
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_793
timestamp 1644511149
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 1644511149
transform 1 0 75164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 1644511149
transform 1 0 75716 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_813
timestamp 1644511149
transform 1 0 75900 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_825
timestamp 1644511149
transform 1 0 77004 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_837
timestamp 1644511149
transform 1 0 78108 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_849
timestamp 1644511149
transform 1 0 79212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_861
timestamp 1644511149
transform 1 0 80316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_867
timestamp 1644511149
transform 1 0 80868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_869
timestamp 1644511149
transform 1 0 81052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_881
timestamp 1644511149
transform 1 0 82156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_893
timestamp 1644511149
transform 1 0 83260 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_905
timestamp 1644511149
transform 1 0 84364 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_917
timestamp 1644511149
transform 1 0 85468 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_923
timestamp 1644511149
transform 1 0 86020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_925
timestamp 1644511149
transform 1 0 86204 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_937
timestamp 1644511149
transform 1 0 87308 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_949
timestamp 1644511149
transform 1 0 88412 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_961
timestamp 1644511149
transform 1 0 89516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_973
timestamp 1644511149
transform 1 0 90620 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_979
timestamp 1644511149
transform 1 0 91172 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_981
timestamp 1644511149
transform 1 0 91356 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_993
timestamp 1644511149
transform 1 0 92460 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1005
timestamp 1644511149
transform 1 0 93564 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1017
timestamp 1644511149
transform 1 0 94668 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1029
timestamp 1644511149
transform 1 0 95772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1035
timestamp 1644511149
transform 1 0 96324 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1037
timestamp 1644511149
transform 1 0 96508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1049
timestamp 1644511149
transform 1 0 97612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1061
timestamp 1644511149
transform 1 0 98716 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1073
timestamp 1644511149
transform 1 0 99820 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1085
timestamp 1644511149
transform 1 0 100924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1091
timestamp 1644511149
transform 1 0 101476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1093
timestamp 1644511149
transform 1 0 101660 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1105
timestamp 1644511149
transform 1 0 102764 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1117
timestamp 1644511149
transform 1 0 103868 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1129
timestamp 1644511149
transform 1 0 104972 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1141
timestamp 1644511149
transform 1 0 106076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1147
timestamp 1644511149
transform 1 0 106628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1149
timestamp 1644511149
transform 1 0 106812 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1161
timestamp 1644511149
transform 1 0 107916 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1173
timestamp 1644511149
transform 1 0 109020 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1185
timestamp 1644511149
transform 1 0 110124 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1197
timestamp 1644511149
transform 1 0 111228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1203
timestamp 1644511149
transform 1 0 111780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1205
timestamp 1644511149
transform 1 0 111964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1217
timestamp 1644511149
transform 1 0 113068 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1229
timestamp 1644511149
transform 1 0 114172 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1241
timestamp 1644511149
transform 1 0 115276 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_1253
timestamp 1644511149
transform 1 0 116380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1259
timestamp 1644511149
transform 1 0 116932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_1261
timestamp 1644511149
transform 1 0 117116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_1273
timestamp 1644511149
transform 1 0 118220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_405
timestamp 1644511149
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_417
timestamp 1644511149
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_429
timestamp 1644511149
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1644511149
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1644511149
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_517
timestamp 1644511149
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_529
timestamp 1644511149
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_541
timestamp 1644511149
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1644511149
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_585
timestamp 1644511149
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_597
timestamp 1644511149
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_629
timestamp 1644511149
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_641
timestamp 1644511149
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_653
timestamp 1644511149
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1644511149
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1644511149
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_673
timestamp 1644511149
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_685
timestamp 1644511149
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_697
timestamp 1644511149
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_709
timestamp 1644511149
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1644511149
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1644511149
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_729
timestamp 1644511149
transform 1 0 68172 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_741
timestamp 1644511149
transform 1 0 69276 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_753
timestamp 1644511149
transform 1 0 70380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_765
timestamp 1644511149
transform 1 0 71484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 1644511149
transform 1 0 72588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1644511149
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_785
timestamp 1644511149
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_797
timestamp 1644511149
transform 1 0 74428 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_809
timestamp 1644511149
transform 1 0 75532 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_821
timestamp 1644511149
transform 1 0 76636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_833
timestamp 1644511149
transform 1 0 77740 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_839
timestamp 1644511149
transform 1 0 78292 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_841
timestamp 1644511149
transform 1 0 78476 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_853
timestamp 1644511149
transform 1 0 79580 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_865
timestamp 1644511149
transform 1 0 80684 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_877
timestamp 1644511149
transform 1 0 81788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_889
timestamp 1644511149
transform 1 0 82892 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_895
timestamp 1644511149
transform 1 0 83444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_897
timestamp 1644511149
transform 1 0 83628 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_909
timestamp 1644511149
transform 1 0 84732 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_921
timestamp 1644511149
transform 1 0 85836 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_933
timestamp 1644511149
transform 1 0 86940 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_945
timestamp 1644511149
transform 1 0 88044 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_951
timestamp 1644511149
transform 1 0 88596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_953
timestamp 1644511149
transform 1 0 88780 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_957
timestamp 1644511149
transform 1 0 89148 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_962
timestamp 1644511149
transform 1 0 89608 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_974
timestamp 1644511149
transform 1 0 90712 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_986
timestamp 1644511149
transform 1 0 91816 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_998
timestamp 1644511149
transform 1 0 92920 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1006
timestamp 1644511149
transform 1 0 93656 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1009
timestamp 1644511149
transform 1 0 93932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1021
timestamp 1644511149
transform 1 0 95036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1033
timestamp 1644511149
transform 1 0 96140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1045
timestamp 1644511149
transform 1 0 97244 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1057
timestamp 1644511149
transform 1 0 98348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1063
timestamp 1644511149
transform 1 0 98900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1065
timestamp 1644511149
transform 1 0 99084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1077
timestamp 1644511149
transform 1 0 100188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1089
timestamp 1644511149
transform 1 0 101292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1101
timestamp 1644511149
transform 1 0 102396 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1113
timestamp 1644511149
transform 1 0 103500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1119
timestamp 1644511149
transform 1 0 104052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1121
timestamp 1644511149
transform 1 0 104236 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1133
timestamp 1644511149
transform 1 0 105340 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1145
timestamp 1644511149
transform 1 0 106444 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1157
timestamp 1644511149
transform 1 0 107548 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1169
timestamp 1644511149
transform 1 0 108652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1175
timestamp 1644511149
transform 1 0 109204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1177
timestamp 1644511149
transform 1 0 109388 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1189
timestamp 1644511149
transform 1 0 110492 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1201
timestamp 1644511149
transform 1 0 111596 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1213
timestamp 1644511149
transform 1 0 112700 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_1225
timestamp 1644511149
transform 1 0 113804 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1231
timestamp 1644511149
transform 1 0 114356 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1233
timestamp 1644511149
transform 1 0 114540 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_1245
timestamp 1644511149
transform 1 0 115644 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_1257
timestamp 1644511149
transform 1 0 116748 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_1267
timestamp 1644511149
transform 1 0 117668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_1273
timestamp 1644511149
transform 1 0 118220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_569
timestamp 1644511149
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1644511149
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1644511149
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_613
timestamp 1644511149
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_625
timestamp 1644511149
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1644511149
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1644511149
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_645
timestamp 1644511149
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_657
timestamp 1644511149
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_669
timestamp 1644511149
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_681
timestamp 1644511149
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1644511149
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1644511149
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_701
timestamp 1644511149
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_713
timestamp 1644511149
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_725
timestamp 1644511149
transform 1 0 67804 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_737
timestamp 1644511149
transform 1 0 68908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_749
timestamp 1644511149
transform 1 0 70012 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_755
timestamp 1644511149
transform 1 0 70564 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_757
timestamp 1644511149
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_769
timestamp 1644511149
transform 1 0 71852 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_781
timestamp 1644511149
transform 1 0 72956 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_793
timestamp 1644511149
transform 1 0 74060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 1644511149
transform 1 0 75164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 1644511149
transform 1 0 75716 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_813
timestamp 1644511149
transform 1 0 75900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_825
timestamp 1644511149
transform 1 0 77004 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_837
timestamp 1644511149
transform 1 0 78108 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_849
timestamp 1644511149
transform 1 0 79212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_861
timestamp 1644511149
transform 1 0 80316 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_867
timestamp 1644511149
transform 1 0 80868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_869
timestamp 1644511149
transform 1 0 81052 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_881
timestamp 1644511149
transform 1 0 82156 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_893
timestamp 1644511149
transform 1 0 83260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_905
timestamp 1644511149
transform 1 0 84364 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_917
timestamp 1644511149
transform 1 0 85468 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_923
timestamp 1644511149
transform 1 0 86020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_925
timestamp 1644511149
transform 1 0 86204 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_937
timestamp 1644511149
transform 1 0 87308 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_949
timestamp 1644511149
transform 1 0 88412 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_961
timestamp 1644511149
transform 1 0 89516 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_973
timestamp 1644511149
transform 1 0 90620 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_979
timestamp 1644511149
transform 1 0 91172 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_981
timestamp 1644511149
transform 1 0 91356 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_993
timestamp 1644511149
transform 1 0 92460 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1005
timestamp 1644511149
transform 1 0 93564 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1017
timestamp 1644511149
transform 1 0 94668 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1029
timestamp 1644511149
transform 1 0 95772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1035
timestamp 1644511149
transform 1 0 96324 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1037
timestamp 1644511149
transform 1 0 96508 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1049
timestamp 1644511149
transform 1 0 97612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1061
timestamp 1644511149
transform 1 0 98716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1073
timestamp 1644511149
transform 1 0 99820 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1085
timestamp 1644511149
transform 1 0 100924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1091
timestamp 1644511149
transform 1 0 101476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1093
timestamp 1644511149
transform 1 0 101660 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1105
timestamp 1644511149
transform 1 0 102764 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1117
timestamp 1644511149
transform 1 0 103868 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1129
timestamp 1644511149
transform 1 0 104972 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1141
timestamp 1644511149
transform 1 0 106076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1147
timestamp 1644511149
transform 1 0 106628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1149
timestamp 1644511149
transform 1 0 106812 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1161
timestamp 1644511149
transform 1 0 107916 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1173
timestamp 1644511149
transform 1 0 109020 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1185
timestamp 1644511149
transform 1 0 110124 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1197
timestamp 1644511149
transform 1 0 111228 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1203
timestamp 1644511149
transform 1 0 111780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1205
timestamp 1644511149
transform 1 0 111964 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1217
timestamp 1644511149
transform 1 0 113068 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1229
timestamp 1644511149
transform 1 0 114172 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1241
timestamp 1644511149
transform 1 0 115276 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_1253
timestamp 1644511149
transform 1 0 116380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1259
timestamp 1644511149
transform 1 0 116932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_1261
timestamp 1644511149
transform 1 0 117116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_1273
timestamp 1644511149
transform 1 0 118220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1644511149
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_541
timestamp 1644511149
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1644511149
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1644511149
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_561
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_573
timestamp 1644511149
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_585
timestamp 1644511149
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_597
timestamp 1644511149
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1644511149
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_617
timestamp 1644511149
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_629
timestamp 1644511149
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_641
timestamp 1644511149
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_653
timestamp 1644511149
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1644511149
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1644511149
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_673
timestamp 1644511149
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_685
timestamp 1644511149
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_697
timestamp 1644511149
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_709
timestamp 1644511149
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1644511149
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1644511149
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_729
timestamp 1644511149
transform 1 0 68172 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_741
timestamp 1644511149
transform 1 0 69276 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_753
timestamp 1644511149
transform 1 0 70380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_765
timestamp 1644511149
transform 1 0 71484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 1644511149
transform 1 0 72588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 1644511149
transform 1 0 73140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_785
timestamp 1644511149
transform 1 0 73324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_797
timestamp 1644511149
transform 1 0 74428 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_809
timestamp 1644511149
transform 1 0 75532 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_821
timestamp 1644511149
transform 1 0 76636 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_833
timestamp 1644511149
transform 1 0 77740 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_839
timestamp 1644511149
transform 1 0 78292 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_841
timestamp 1644511149
transform 1 0 78476 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_853
timestamp 1644511149
transform 1 0 79580 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_865
timestamp 1644511149
transform 1 0 80684 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_877
timestamp 1644511149
transform 1 0 81788 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_889
timestamp 1644511149
transform 1 0 82892 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_895
timestamp 1644511149
transform 1 0 83444 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_897
timestamp 1644511149
transform 1 0 83628 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_909
timestamp 1644511149
transform 1 0 84732 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_921
timestamp 1644511149
transform 1 0 85836 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_933
timestamp 1644511149
transform 1 0 86940 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_945
timestamp 1644511149
transform 1 0 88044 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_951
timestamp 1644511149
transform 1 0 88596 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_953
timestamp 1644511149
transform 1 0 88780 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_965
timestamp 1644511149
transform 1 0 89884 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_977
timestamp 1644511149
transform 1 0 90988 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_989
timestamp 1644511149
transform 1 0 92092 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1001
timestamp 1644511149
transform 1 0 93196 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1007
timestamp 1644511149
transform 1 0 93748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1009
timestamp 1644511149
transform 1 0 93932 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1021
timestamp 1644511149
transform 1 0 95036 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1033
timestamp 1644511149
transform 1 0 96140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1045
timestamp 1644511149
transform 1 0 97244 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1057
timestamp 1644511149
transform 1 0 98348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1063
timestamp 1644511149
transform 1 0 98900 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1065
timestamp 1644511149
transform 1 0 99084 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1077
timestamp 1644511149
transform 1 0 100188 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1089
timestamp 1644511149
transform 1 0 101292 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1101
timestamp 1644511149
transform 1 0 102396 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1113
timestamp 1644511149
transform 1 0 103500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1119
timestamp 1644511149
transform 1 0 104052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1121
timestamp 1644511149
transform 1 0 104236 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1133
timestamp 1644511149
transform 1 0 105340 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1145
timestamp 1644511149
transform 1 0 106444 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1157
timestamp 1644511149
transform 1 0 107548 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1169
timestamp 1644511149
transform 1 0 108652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1175
timestamp 1644511149
transform 1 0 109204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1177
timestamp 1644511149
transform 1 0 109388 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1189
timestamp 1644511149
transform 1 0 110492 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1201
timestamp 1644511149
transform 1 0 111596 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1213
timestamp 1644511149
transform 1 0 112700 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_1225
timestamp 1644511149
transform 1 0 113804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1231
timestamp 1644511149
transform 1 0 114356 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1233
timestamp 1644511149
transform 1 0 114540 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_1245
timestamp 1644511149
transform 1 0 115644 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_1257
timestamp 1644511149
transform 1 0 116748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_1267
timestamp 1644511149
transform 1 0 117668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_1273
timestamp 1644511149
transform 1 0 118220 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_501
timestamp 1644511149
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_513
timestamp 1644511149
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1644511149
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1644511149
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_533
timestamp 1644511149
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_545
timestamp 1644511149
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_557
timestamp 1644511149
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_569
timestamp 1644511149
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1644511149
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1644511149
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_601
timestamp 1644511149
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_613
timestamp 1644511149
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_625
timestamp 1644511149
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1644511149
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1644511149
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_645
timestamp 1644511149
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_657
timestamp 1644511149
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_669
timestamp 1644511149
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_681
timestamp 1644511149
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1644511149
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1644511149
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_701
timestamp 1644511149
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_713
timestamp 1644511149
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_725
timestamp 1644511149
transform 1 0 67804 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_737
timestamp 1644511149
transform 1 0 68908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 1644511149
transform 1 0 70012 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 1644511149
transform 1 0 70564 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_757
timestamp 1644511149
transform 1 0 70748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_769
timestamp 1644511149
transform 1 0 71852 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_781
timestamp 1644511149
transform 1 0 72956 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_793
timestamp 1644511149
transform 1 0 74060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_805
timestamp 1644511149
transform 1 0 75164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_811
timestamp 1644511149
transform 1 0 75716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_813
timestamp 1644511149
transform 1 0 75900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_825
timestamp 1644511149
transform 1 0 77004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_837
timestamp 1644511149
transform 1 0 78108 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_849
timestamp 1644511149
transform 1 0 79212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_861
timestamp 1644511149
transform 1 0 80316 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_867
timestamp 1644511149
transform 1 0 80868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_869
timestamp 1644511149
transform 1 0 81052 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_881
timestamp 1644511149
transform 1 0 82156 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_893
timestamp 1644511149
transform 1 0 83260 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_905
timestamp 1644511149
transform 1 0 84364 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_917
timestamp 1644511149
transform 1 0 85468 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_923
timestamp 1644511149
transform 1 0 86020 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_925
timestamp 1644511149
transform 1 0 86204 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_937
timestamp 1644511149
transform 1 0 87308 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_949
timestamp 1644511149
transform 1 0 88412 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_961
timestamp 1644511149
transform 1 0 89516 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_973
timestamp 1644511149
transform 1 0 90620 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_979
timestamp 1644511149
transform 1 0 91172 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_981
timestamp 1644511149
transform 1 0 91356 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_993
timestamp 1644511149
transform 1 0 92460 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1005
timestamp 1644511149
transform 1 0 93564 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1017
timestamp 1644511149
transform 1 0 94668 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1029
timestamp 1644511149
transform 1 0 95772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1035
timestamp 1644511149
transform 1 0 96324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1037
timestamp 1644511149
transform 1 0 96508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1049
timestamp 1644511149
transform 1 0 97612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1061
timestamp 1644511149
transform 1 0 98716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1073
timestamp 1644511149
transform 1 0 99820 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1085
timestamp 1644511149
transform 1 0 100924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1091
timestamp 1644511149
transform 1 0 101476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1093
timestamp 1644511149
transform 1 0 101660 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1105
timestamp 1644511149
transform 1 0 102764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1117
timestamp 1644511149
transform 1 0 103868 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1129
timestamp 1644511149
transform 1 0 104972 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1141
timestamp 1644511149
transform 1 0 106076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1147
timestamp 1644511149
transform 1 0 106628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1149
timestamp 1644511149
transform 1 0 106812 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1161
timestamp 1644511149
transform 1 0 107916 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1173
timestamp 1644511149
transform 1 0 109020 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1185
timestamp 1644511149
transform 1 0 110124 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1197
timestamp 1644511149
transform 1 0 111228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1203
timestamp 1644511149
transform 1 0 111780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1205
timestamp 1644511149
transform 1 0 111964 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1217
timestamp 1644511149
transform 1 0 113068 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1229
timestamp 1644511149
transform 1 0 114172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_1241
timestamp 1644511149
transform 1 0 115276 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_1253
timestamp 1644511149
transform 1 0 116380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1259
timestamp 1644511149
transform 1 0 116932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_1261
timestamp 1644511149
transform 1 0 117116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_1267
timestamp 1644511149
transform 1 0 117668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_1273
timestamp 1644511149
transform 1 0 118220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1644511149
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_517
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_529
timestamp 1644511149
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_541
timestamp 1644511149
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1644511149
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1644511149
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_561
timestamp 1644511149
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_573
timestamp 1644511149
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_585
timestamp 1644511149
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_597
timestamp 1644511149
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1644511149
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1644511149
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_629
timestamp 1644511149
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_641
timestamp 1644511149
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_653
timestamp 1644511149
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1644511149
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1644511149
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_673
timestamp 1644511149
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_685
timestamp 1644511149
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_697
timestamp 1644511149
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_709
timestamp 1644511149
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1644511149
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1644511149
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_729
timestamp 1644511149
transform 1 0 68172 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_741
timestamp 1644511149
transform 1 0 69276 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_753
timestamp 1644511149
transform 1 0 70380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_765
timestamp 1644511149
transform 1 0 71484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_777
timestamp 1644511149
transform 1 0 72588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 1644511149
transform 1 0 73140 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_785
timestamp 1644511149
transform 1 0 73324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_797
timestamp 1644511149
transform 1 0 74428 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_809
timestamp 1644511149
transform 1 0 75532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_821
timestamp 1644511149
transform 1 0 76636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_833
timestamp 1644511149
transform 1 0 77740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_839
timestamp 1644511149
transform 1 0 78292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_841
timestamp 1644511149
transform 1 0 78476 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_853
timestamp 1644511149
transform 1 0 79580 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_865
timestamp 1644511149
transform 1 0 80684 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_877
timestamp 1644511149
transform 1 0 81788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_889
timestamp 1644511149
transform 1 0 82892 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_895
timestamp 1644511149
transform 1 0 83444 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_897
timestamp 1644511149
transform 1 0 83628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_909
timestamp 1644511149
transform 1 0 84732 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_921
timestamp 1644511149
transform 1 0 85836 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_933
timestamp 1644511149
transform 1 0 86940 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_945
timestamp 1644511149
transform 1 0 88044 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_951
timestamp 1644511149
transform 1 0 88596 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_953
timestamp 1644511149
transform 1 0 88780 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_965
timestamp 1644511149
transform 1 0 89884 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_977
timestamp 1644511149
transform 1 0 90988 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_989
timestamp 1644511149
transform 1 0 92092 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1001
timestamp 1644511149
transform 1 0 93196 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1007
timestamp 1644511149
transform 1 0 93748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1009
timestamp 1644511149
transform 1 0 93932 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1021
timestamp 1644511149
transform 1 0 95036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1033
timestamp 1644511149
transform 1 0 96140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1045
timestamp 1644511149
transform 1 0 97244 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1057
timestamp 1644511149
transform 1 0 98348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1063
timestamp 1644511149
transform 1 0 98900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1065
timestamp 1644511149
transform 1 0 99084 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1077
timestamp 1644511149
transform 1 0 100188 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1089
timestamp 1644511149
transform 1 0 101292 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1101
timestamp 1644511149
transform 1 0 102396 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1113
timestamp 1644511149
transform 1 0 103500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1119
timestamp 1644511149
transform 1 0 104052 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1121
timestamp 1644511149
transform 1 0 104236 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1133
timestamp 1644511149
transform 1 0 105340 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1145
timestamp 1644511149
transform 1 0 106444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1157
timestamp 1644511149
transform 1 0 107548 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1169
timestamp 1644511149
transform 1 0 108652 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1175
timestamp 1644511149
transform 1 0 109204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1177
timestamp 1644511149
transform 1 0 109388 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1189
timestamp 1644511149
transform 1 0 110492 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1201
timestamp 1644511149
transform 1 0 111596 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1213
timestamp 1644511149
transform 1 0 112700 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_1225
timestamp 1644511149
transform 1 0 113804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1231
timestamp 1644511149
transform 1 0 114356 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1233
timestamp 1644511149
transform 1 0 114540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1245
timestamp 1644511149
transform 1 0 115644 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_1257
timestamp 1644511149
transform 1 0 116748 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_1269
timestamp 1644511149
transform 1 0 117852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_501
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_513
timestamp 1644511149
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1644511149
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1644511149
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_533
timestamp 1644511149
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_545
timestamp 1644511149
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_557
timestamp 1644511149
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_569
timestamp 1644511149
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1644511149
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1644511149
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_613
timestamp 1644511149
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_625
timestamp 1644511149
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1644511149
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1644511149
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_645
timestamp 1644511149
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_657
timestamp 1644511149
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_669
timestamp 1644511149
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_681
timestamp 1644511149
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1644511149
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1644511149
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_701
timestamp 1644511149
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_713
timestamp 1644511149
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_725
timestamp 1644511149
transform 1 0 67804 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_737
timestamp 1644511149
transform 1 0 68908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_749
timestamp 1644511149
transform 1 0 70012 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_755
timestamp 1644511149
transform 1 0 70564 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_757
timestamp 1644511149
transform 1 0 70748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_769
timestamp 1644511149
transform 1 0 71852 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_781
timestamp 1644511149
transform 1 0 72956 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_793
timestamp 1644511149
transform 1 0 74060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_805
timestamp 1644511149
transform 1 0 75164 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_811
timestamp 1644511149
transform 1 0 75716 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_813
timestamp 1644511149
transform 1 0 75900 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_825
timestamp 1644511149
transform 1 0 77004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_837
timestamp 1644511149
transform 1 0 78108 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_849
timestamp 1644511149
transform 1 0 79212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_861
timestamp 1644511149
transform 1 0 80316 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_867
timestamp 1644511149
transform 1 0 80868 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_869
timestamp 1644511149
transform 1 0 81052 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_881
timestamp 1644511149
transform 1 0 82156 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_893
timestamp 1644511149
transform 1 0 83260 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_905
timestamp 1644511149
transform 1 0 84364 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_917
timestamp 1644511149
transform 1 0 85468 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_923
timestamp 1644511149
transform 1 0 86020 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_925
timestamp 1644511149
transform 1 0 86204 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_937
timestamp 1644511149
transform 1 0 87308 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_949
timestamp 1644511149
transform 1 0 88412 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_961
timestamp 1644511149
transform 1 0 89516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_973
timestamp 1644511149
transform 1 0 90620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_979
timestamp 1644511149
transform 1 0 91172 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_981
timestamp 1644511149
transform 1 0 91356 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_993
timestamp 1644511149
transform 1 0 92460 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1005
timestamp 1644511149
transform 1 0 93564 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1017
timestamp 1644511149
transform 1 0 94668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1029
timestamp 1644511149
transform 1 0 95772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1035
timestamp 1644511149
transform 1 0 96324 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1037
timestamp 1644511149
transform 1 0 96508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1049
timestamp 1644511149
transform 1 0 97612 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1061
timestamp 1644511149
transform 1 0 98716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1073
timestamp 1644511149
transform 1 0 99820 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1085
timestamp 1644511149
transform 1 0 100924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1091
timestamp 1644511149
transform 1 0 101476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1093
timestamp 1644511149
transform 1 0 101660 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1105
timestamp 1644511149
transform 1 0 102764 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1117
timestamp 1644511149
transform 1 0 103868 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1129
timestamp 1644511149
transform 1 0 104972 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1141
timestamp 1644511149
transform 1 0 106076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1147
timestamp 1644511149
transform 1 0 106628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1149
timestamp 1644511149
transform 1 0 106812 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1161
timestamp 1644511149
transform 1 0 107916 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1173
timestamp 1644511149
transform 1 0 109020 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1185
timestamp 1644511149
transform 1 0 110124 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1197
timestamp 1644511149
transform 1 0 111228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1203
timestamp 1644511149
transform 1 0 111780 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1205
timestamp 1644511149
transform 1 0 111964 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1217
timestamp 1644511149
transform 1 0 113068 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1229
timestamp 1644511149
transform 1 0 114172 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_1241
timestamp 1644511149
transform 1 0 115276 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_1253
timestamp 1644511149
transform 1 0 116380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1259
timestamp 1644511149
transform 1 0 116932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_1261
timestamp 1644511149
transform 1 0 117116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_1267
timestamp 1644511149
transform 1 0 117668 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_1273
timestamp 1644511149
transform 1 0 118220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_561
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_573
timestamp 1644511149
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_585
timestamp 1644511149
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1644511149
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1644511149
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_629
timestamp 1644511149
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_641
timestamp 1644511149
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_653
timestamp 1644511149
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1644511149
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1644511149
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_673
timestamp 1644511149
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_685
timestamp 1644511149
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_697
timestamp 1644511149
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_709
timestamp 1644511149
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1644511149
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1644511149
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_729
timestamp 1644511149
transform 1 0 68172 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_741
timestamp 1644511149
transform 1 0 69276 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_753
timestamp 1644511149
transform 1 0 70380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_765
timestamp 1644511149
transform 1 0 71484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_777
timestamp 1644511149
transform 1 0 72588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 1644511149
transform 1 0 73140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_785
timestamp 1644511149
transform 1 0 73324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_797
timestamp 1644511149
transform 1 0 74428 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_809
timestamp 1644511149
transform 1 0 75532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_821
timestamp 1644511149
transform 1 0 76636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_833
timestamp 1644511149
transform 1 0 77740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_839
timestamp 1644511149
transform 1 0 78292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_841
timestamp 1644511149
transform 1 0 78476 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_853
timestamp 1644511149
transform 1 0 79580 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_865
timestamp 1644511149
transform 1 0 80684 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_877
timestamp 1644511149
transform 1 0 81788 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_889
timestamp 1644511149
transform 1 0 82892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_895
timestamp 1644511149
transform 1 0 83444 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_897
timestamp 1644511149
transform 1 0 83628 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_909
timestamp 1644511149
transform 1 0 84732 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_921
timestamp 1644511149
transform 1 0 85836 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_933
timestamp 1644511149
transform 1 0 86940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_945
timestamp 1644511149
transform 1 0 88044 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_951
timestamp 1644511149
transform 1 0 88596 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_953
timestamp 1644511149
transform 1 0 88780 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_965
timestamp 1644511149
transform 1 0 89884 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_977
timestamp 1644511149
transform 1 0 90988 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_989
timestamp 1644511149
transform 1 0 92092 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1001
timestamp 1644511149
transform 1 0 93196 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1007
timestamp 1644511149
transform 1 0 93748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1009
timestamp 1644511149
transform 1 0 93932 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1021
timestamp 1644511149
transform 1 0 95036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1033
timestamp 1644511149
transform 1 0 96140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1045
timestamp 1644511149
transform 1 0 97244 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1057
timestamp 1644511149
transform 1 0 98348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1063
timestamp 1644511149
transform 1 0 98900 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1065
timestamp 1644511149
transform 1 0 99084 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1077
timestamp 1644511149
transform 1 0 100188 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1089
timestamp 1644511149
transform 1 0 101292 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1101
timestamp 1644511149
transform 1 0 102396 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1113
timestamp 1644511149
transform 1 0 103500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1119
timestamp 1644511149
transform 1 0 104052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1121
timestamp 1644511149
transform 1 0 104236 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1133
timestamp 1644511149
transform 1 0 105340 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1145
timestamp 1644511149
transform 1 0 106444 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1157
timestamp 1644511149
transform 1 0 107548 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1169
timestamp 1644511149
transform 1 0 108652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1175
timestamp 1644511149
transform 1 0 109204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1177
timestamp 1644511149
transform 1 0 109388 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1189
timestamp 1644511149
transform 1 0 110492 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1201
timestamp 1644511149
transform 1 0 111596 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1213
timestamp 1644511149
transform 1 0 112700 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_1225
timestamp 1644511149
transform 1 0 113804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1231
timestamp 1644511149
transform 1 0 114356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1233
timestamp 1644511149
transform 1 0 114540 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1245
timestamp 1644511149
transform 1 0 115644 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_1257
timestamp 1644511149
transform 1 0 116748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_1269
timestamp 1644511149
transform 1 0 117852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_533
timestamp 1644511149
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_557
timestamp 1644511149
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_569
timestamp 1644511149
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_601
timestamp 1644511149
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_613
timestamp 1644511149
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_625
timestamp 1644511149
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1644511149
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1644511149
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_645
timestamp 1644511149
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_657
timestamp 1644511149
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_669
timestamp 1644511149
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_681
timestamp 1644511149
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1644511149
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1644511149
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_701
timestamp 1644511149
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_713
timestamp 1644511149
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_725
timestamp 1644511149
transform 1 0 67804 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_737
timestamp 1644511149
transform 1 0 68908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_749
timestamp 1644511149
transform 1 0 70012 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 1644511149
transform 1 0 70564 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_757
timestamp 1644511149
transform 1 0 70748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_769
timestamp 1644511149
transform 1 0 71852 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_781
timestamp 1644511149
transform 1 0 72956 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_793
timestamp 1644511149
transform 1 0 74060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_805
timestamp 1644511149
transform 1 0 75164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 1644511149
transform 1 0 75716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_813
timestamp 1644511149
transform 1 0 75900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_825
timestamp 1644511149
transform 1 0 77004 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_837
timestamp 1644511149
transform 1 0 78108 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_849
timestamp 1644511149
transform 1 0 79212 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_861
timestamp 1644511149
transform 1 0 80316 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_867
timestamp 1644511149
transform 1 0 80868 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_869
timestamp 1644511149
transform 1 0 81052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_881
timestamp 1644511149
transform 1 0 82156 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_893
timestamp 1644511149
transform 1 0 83260 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_905
timestamp 1644511149
transform 1 0 84364 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_917
timestamp 1644511149
transform 1 0 85468 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_923
timestamp 1644511149
transform 1 0 86020 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_925
timestamp 1644511149
transform 1 0 86204 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_937
timestamp 1644511149
transform 1 0 87308 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_949
timestamp 1644511149
transform 1 0 88412 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_961
timestamp 1644511149
transform 1 0 89516 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_973
timestamp 1644511149
transform 1 0 90620 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_979
timestamp 1644511149
transform 1 0 91172 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_981
timestamp 1644511149
transform 1 0 91356 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_993
timestamp 1644511149
transform 1 0 92460 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1005
timestamp 1644511149
transform 1 0 93564 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1017
timestamp 1644511149
transform 1 0 94668 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1029
timestamp 1644511149
transform 1 0 95772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1035
timestamp 1644511149
transform 1 0 96324 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1037
timestamp 1644511149
transform 1 0 96508 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1049
timestamp 1644511149
transform 1 0 97612 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1061
timestamp 1644511149
transform 1 0 98716 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1073
timestamp 1644511149
transform 1 0 99820 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1085
timestamp 1644511149
transform 1 0 100924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1091
timestamp 1644511149
transform 1 0 101476 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1093
timestamp 1644511149
transform 1 0 101660 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1105
timestamp 1644511149
transform 1 0 102764 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1117
timestamp 1644511149
transform 1 0 103868 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1129
timestamp 1644511149
transform 1 0 104972 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1141
timestamp 1644511149
transform 1 0 106076 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1147
timestamp 1644511149
transform 1 0 106628 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1149
timestamp 1644511149
transform 1 0 106812 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1161
timestamp 1644511149
transform 1 0 107916 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1173
timestamp 1644511149
transform 1 0 109020 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1185
timestamp 1644511149
transform 1 0 110124 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1197
timestamp 1644511149
transform 1 0 111228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1203
timestamp 1644511149
transform 1 0 111780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1205
timestamp 1644511149
transform 1 0 111964 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1217
timestamp 1644511149
transform 1 0 113068 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1229
timestamp 1644511149
transform 1 0 114172 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_1241
timestamp 1644511149
transform 1 0 115276 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_1253
timestamp 1644511149
transform 1 0 116380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1259
timestamp 1644511149
transform 1 0 116932 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_1261
timestamp 1644511149
transform 1 0 117116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_1267
timestamp 1644511149
transform 1 0 117668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_1273
timestamp 1644511149
transform 1 0 118220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_517
timestamp 1644511149
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_529
timestamp 1644511149
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1644511149
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1644511149
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_561
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_573
timestamp 1644511149
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_585
timestamp 1644511149
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_597
timestamp 1644511149
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1644511149
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1644511149
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_629
timestamp 1644511149
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_641
timestamp 1644511149
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_653
timestamp 1644511149
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1644511149
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1644511149
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_673
timestamp 1644511149
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_685
timestamp 1644511149
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_697
timestamp 1644511149
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_709
timestamp 1644511149
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1644511149
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1644511149
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_729
timestamp 1644511149
transform 1 0 68172 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_741
timestamp 1644511149
transform 1 0 69276 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_753
timestamp 1644511149
transform 1 0 70380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_765
timestamp 1644511149
transform 1 0 71484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 1644511149
transform 1 0 72588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 1644511149
transform 1 0 73140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_785
timestamp 1644511149
transform 1 0 73324 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_797
timestamp 1644511149
transform 1 0 74428 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_809
timestamp 1644511149
transform 1 0 75532 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_821
timestamp 1644511149
transform 1 0 76636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_833
timestamp 1644511149
transform 1 0 77740 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_839
timestamp 1644511149
transform 1 0 78292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_841
timestamp 1644511149
transform 1 0 78476 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_853
timestamp 1644511149
transform 1 0 79580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_865
timestamp 1644511149
transform 1 0 80684 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_877
timestamp 1644511149
transform 1 0 81788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_889
timestamp 1644511149
transform 1 0 82892 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_895
timestamp 1644511149
transform 1 0 83444 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_897
timestamp 1644511149
transform 1 0 83628 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_909
timestamp 1644511149
transform 1 0 84732 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_921
timestamp 1644511149
transform 1 0 85836 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_933
timestamp 1644511149
transform 1 0 86940 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_945
timestamp 1644511149
transform 1 0 88044 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_951
timestamp 1644511149
transform 1 0 88596 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_953
timestamp 1644511149
transform 1 0 88780 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_965
timestamp 1644511149
transform 1 0 89884 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_977
timestamp 1644511149
transform 1 0 90988 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_989
timestamp 1644511149
transform 1 0 92092 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1001
timestamp 1644511149
transform 1 0 93196 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1007
timestamp 1644511149
transform 1 0 93748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1009
timestamp 1644511149
transform 1 0 93932 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1021
timestamp 1644511149
transform 1 0 95036 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1033
timestamp 1644511149
transform 1 0 96140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1045
timestamp 1644511149
transform 1 0 97244 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1057
timestamp 1644511149
transform 1 0 98348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1063
timestamp 1644511149
transform 1 0 98900 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1065
timestamp 1644511149
transform 1 0 99084 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1077
timestamp 1644511149
transform 1 0 100188 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1089
timestamp 1644511149
transform 1 0 101292 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1101
timestamp 1644511149
transform 1 0 102396 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1113
timestamp 1644511149
transform 1 0 103500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1119
timestamp 1644511149
transform 1 0 104052 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1121
timestamp 1644511149
transform 1 0 104236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1133
timestamp 1644511149
transform 1 0 105340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1145
timestamp 1644511149
transform 1 0 106444 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1157
timestamp 1644511149
transform 1 0 107548 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1169
timestamp 1644511149
transform 1 0 108652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1175
timestamp 1644511149
transform 1 0 109204 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1177
timestamp 1644511149
transform 1 0 109388 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1189
timestamp 1644511149
transform 1 0 110492 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1201
timestamp 1644511149
transform 1 0 111596 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1213
timestamp 1644511149
transform 1 0 112700 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_1225
timestamp 1644511149
transform 1 0 113804 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1231
timestamp 1644511149
transform 1 0 114356 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1233
timestamp 1644511149
transform 1 0 114540 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1245
timestamp 1644511149
transform 1 0 115644 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_1257
timestamp 1644511149
transform 1 0 116748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_1269
timestamp 1644511149
transform 1 0 117852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_277
timestamp 1644511149
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_321
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_333
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_345
timestamp 1644511149
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1644511149
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_513
timestamp 1644511149
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1644511149
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1644511149
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_569
timestamp 1644511149
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1644511149
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_613
timestamp 1644511149
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_625
timestamp 1644511149
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1644511149
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1644511149
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_645
timestamp 1644511149
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_657
timestamp 1644511149
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_669
timestamp 1644511149
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_681
timestamp 1644511149
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1644511149
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1644511149
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_701
timestamp 1644511149
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_713
timestamp 1644511149
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_725
timestamp 1644511149
transform 1 0 67804 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_737
timestamp 1644511149
transform 1 0 68908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 1644511149
transform 1 0 70012 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 1644511149
transform 1 0 70564 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_757
timestamp 1644511149
transform 1 0 70748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_769
timestamp 1644511149
transform 1 0 71852 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_781
timestamp 1644511149
transform 1 0 72956 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_793
timestamp 1644511149
transform 1 0 74060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 1644511149
transform 1 0 75164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 1644511149
transform 1 0 75716 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_813
timestamp 1644511149
transform 1 0 75900 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_825
timestamp 1644511149
transform 1 0 77004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_837
timestamp 1644511149
transform 1 0 78108 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_849
timestamp 1644511149
transform 1 0 79212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_861
timestamp 1644511149
transform 1 0 80316 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_867
timestamp 1644511149
transform 1 0 80868 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_869
timestamp 1644511149
transform 1 0 81052 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_881
timestamp 1644511149
transform 1 0 82156 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_893
timestamp 1644511149
transform 1 0 83260 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_905
timestamp 1644511149
transform 1 0 84364 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_917
timestamp 1644511149
transform 1 0 85468 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_923
timestamp 1644511149
transform 1 0 86020 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_925
timestamp 1644511149
transform 1 0 86204 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_937
timestamp 1644511149
transform 1 0 87308 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_949
timestamp 1644511149
transform 1 0 88412 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_961
timestamp 1644511149
transform 1 0 89516 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_973
timestamp 1644511149
transform 1 0 90620 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_979
timestamp 1644511149
transform 1 0 91172 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_981
timestamp 1644511149
transform 1 0 91356 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_993
timestamp 1644511149
transform 1 0 92460 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1005
timestamp 1644511149
transform 1 0 93564 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1017
timestamp 1644511149
transform 1 0 94668 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1029
timestamp 1644511149
transform 1 0 95772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1035
timestamp 1644511149
transform 1 0 96324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1037
timestamp 1644511149
transform 1 0 96508 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1049
timestamp 1644511149
transform 1 0 97612 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1061
timestamp 1644511149
transform 1 0 98716 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1073
timestamp 1644511149
transform 1 0 99820 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1085
timestamp 1644511149
transform 1 0 100924 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1091
timestamp 1644511149
transform 1 0 101476 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1093
timestamp 1644511149
transform 1 0 101660 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1105
timestamp 1644511149
transform 1 0 102764 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1117
timestamp 1644511149
transform 1 0 103868 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1129
timestamp 1644511149
transform 1 0 104972 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1141
timestamp 1644511149
transform 1 0 106076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1147
timestamp 1644511149
transform 1 0 106628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1149
timestamp 1644511149
transform 1 0 106812 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1161
timestamp 1644511149
transform 1 0 107916 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1173
timestamp 1644511149
transform 1 0 109020 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1185
timestamp 1644511149
transform 1 0 110124 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1197
timestamp 1644511149
transform 1 0 111228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1203
timestamp 1644511149
transform 1 0 111780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1205
timestamp 1644511149
transform 1 0 111964 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1217
timestamp 1644511149
transform 1 0 113068 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1229
timestamp 1644511149
transform 1 0 114172 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_1241
timestamp 1644511149
transform 1 0 115276 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_1253
timestamp 1644511149
transform 1 0 116380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1259
timestamp 1644511149
transform 1 0 116932 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_1261
timestamp 1644511149
transform 1 0 117116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_1267
timestamp 1644511149
transform 1 0 117668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_1273
timestamp 1644511149
transform 1 0 118220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_193
timestamp 1644511149
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_205
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_305
timestamp 1644511149
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1644511149
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_529
timestamp 1644511149
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_541
timestamp 1644511149
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1644511149
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1644511149
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_573
timestamp 1644511149
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_585
timestamp 1644511149
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_597
timestamp 1644511149
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1644511149
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1644511149
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_617
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_629
timestamp 1644511149
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_641
timestamp 1644511149
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_653
timestamp 1644511149
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1644511149
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1644511149
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_673
timestamp 1644511149
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_685
timestamp 1644511149
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_697
timestamp 1644511149
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_709
timestamp 1644511149
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1644511149
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1644511149
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_729
timestamp 1644511149
transform 1 0 68172 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_741
timestamp 1644511149
transform 1 0 69276 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_753
timestamp 1644511149
transform 1 0 70380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_765
timestamp 1644511149
transform 1 0 71484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 1644511149
transform 1 0 72588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 1644511149
transform 1 0 73140 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_785
timestamp 1644511149
transform 1 0 73324 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_797
timestamp 1644511149
transform 1 0 74428 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_809
timestamp 1644511149
transform 1 0 75532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_821
timestamp 1644511149
transform 1 0 76636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_833
timestamp 1644511149
transform 1 0 77740 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_839
timestamp 1644511149
transform 1 0 78292 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_841
timestamp 1644511149
transform 1 0 78476 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_853
timestamp 1644511149
transform 1 0 79580 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_865
timestamp 1644511149
transform 1 0 80684 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_877
timestamp 1644511149
transform 1 0 81788 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_889
timestamp 1644511149
transform 1 0 82892 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_895
timestamp 1644511149
transform 1 0 83444 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_897
timestamp 1644511149
transform 1 0 83628 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_909
timestamp 1644511149
transform 1 0 84732 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_921
timestamp 1644511149
transform 1 0 85836 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_933
timestamp 1644511149
transform 1 0 86940 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_945
timestamp 1644511149
transform 1 0 88044 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_951
timestamp 1644511149
transform 1 0 88596 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_953
timestamp 1644511149
transform 1 0 88780 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_965
timestamp 1644511149
transform 1 0 89884 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_977
timestamp 1644511149
transform 1 0 90988 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_989
timestamp 1644511149
transform 1 0 92092 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1001
timestamp 1644511149
transform 1 0 93196 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1007
timestamp 1644511149
transform 1 0 93748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1009
timestamp 1644511149
transform 1 0 93932 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1021
timestamp 1644511149
transform 1 0 95036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1033
timestamp 1644511149
transform 1 0 96140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1045
timestamp 1644511149
transform 1 0 97244 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1057
timestamp 1644511149
transform 1 0 98348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1063
timestamp 1644511149
transform 1 0 98900 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1065
timestamp 1644511149
transform 1 0 99084 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1077
timestamp 1644511149
transform 1 0 100188 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1089
timestamp 1644511149
transform 1 0 101292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1101
timestamp 1644511149
transform 1 0 102396 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1113
timestamp 1644511149
transform 1 0 103500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1119
timestamp 1644511149
transform 1 0 104052 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1121
timestamp 1644511149
transform 1 0 104236 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1133
timestamp 1644511149
transform 1 0 105340 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1145
timestamp 1644511149
transform 1 0 106444 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1157
timestamp 1644511149
transform 1 0 107548 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1169
timestamp 1644511149
transform 1 0 108652 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1175
timestamp 1644511149
transform 1 0 109204 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1177
timestamp 1644511149
transform 1 0 109388 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1189
timestamp 1644511149
transform 1 0 110492 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1201
timestamp 1644511149
transform 1 0 111596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1213
timestamp 1644511149
transform 1 0 112700 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1225
timestamp 1644511149
transform 1 0 113804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_1231
timestamp 1644511149
transform 1 0 114356 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1233
timestamp 1644511149
transform 1 0 114540 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_1245
timestamp 1644511149
transform 1 0 115644 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_1257
timestamp 1644511149
transform 1 0 116748 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_1267
timestamp 1644511149
transform 1 0 117668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_1273
timestamp 1644511149
transform 1 0 118220 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1644511149
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1644511149
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_333
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_345
timestamp 1644511149
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1644511149
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_533
timestamp 1644511149
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_545
timestamp 1644511149
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_557
timestamp 1644511149
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_569
timestamp 1644511149
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1644511149
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1644511149
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_601
timestamp 1644511149
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_625
timestamp 1644511149
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1644511149
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1644511149
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_645
timestamp 1644511149
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_657
timestamp 1644511149
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_669
timestamp 1644511149
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_681
timestamp 1644511149
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1644511149
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1644511149
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_701
timestamp 1644511149
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_713
timestamp 1644511149
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_725
timestamp 1644511149
transform 1 0 67804 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_737
timestamp 1644511149
transform 1 0 68908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 1644511149
transform 1 0 70012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 1644511149
transform 1 0 70564 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_757
timestamp 1644511149
transform 1 0 70748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_769
timestamp 1644511149
transform 1 0 71852 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_781
timestamp 1644511149
transform 1 0 72956 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_793
timestamp 1644511149
transform 1 0 74060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 1644511149
transform 1 0 75164 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 1644511149
transform 1 0 75716 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_813
timestamp 1644511149
transform 1 0 75900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_825
timestamp 1644511149
transform 1 0 77004 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_837
timestamp 1644511149
transform 1 0 78108 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_849
timestamp 1644511149
transform 1 0 79212 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_861
timestamp 1644511149
transform 1 0 80316 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_867
timestamp 1644511149
transform 1 0 80868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_869
timestamp 1644511149
transform 1 0 81052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_881
timestamp 1644511149
transform 1 0 82156 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_893
timestamp 1644511149
transform 1 0 83260 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_905
timestamp 1644511149
transform 1 0 84364 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_917
timestamp 1644511149
transform 1 0 85468 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_923
timestamp 1644511149
transform 1 0 86020 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_925
timestamp 1644511149
transform 1 0 86204 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_937
timestamp 1644511149
transform 1 0 87308 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_949
timestamp 1644511149
transform 1 0 88412 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_961
timestamp 1644511149
transform 1 0 89516 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_973
timestamp 1644511149
transform 1 0 90620 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_979
timestamp 1644511149
transform 1 0 91172 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_981
timestamp 1644511149
transform 1 0 91356 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_993
timestamp 1644511149
transform 1 0 92460 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1005
timestamp 1644511149
transform 1 0 93564 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1017
timestamp 1644511149
transform 1 0 94668 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1029
timestamp 1644511149
transform 1 0 95772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1035
timestamp 1644511149
transform 1 0 96324 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1037
timestamp 1644511149
transform 1 0 96508 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1049
timestamp 1644511149
transform 1 0 97612 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1061
timestamp 1644511149
transform 1 0 98716 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1073
timestamp 1644511149
transform 1 0 99820 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1085
timestamp 1644511149
transform 1 0 100924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1091
timestamp 1644511149
transform 1 0 101476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1093
timestamp 1644511149
transform 1 0 101660 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1105
timestamp 1644511149
transform 1 0 102764 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1117
timestamp 1644511149
transform 1 0 103868 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1129
timestamp 1644511149
transform 1 0 104972 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1141
timestamp 1644511149
transform 1 0 106076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1147
timestamp 1644511149
transform 1 0 106628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1149
timestamp 1644511149
transform 1 0 106812 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1161
timestamp 1644511149
transform 1 0 107916 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1173
timestamp 1644511149
transform 1 0 109020 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1185
timestamp 1644511149
transform 1 0 110124 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1197
timestamp 1644511149
transform 1 0 111228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1203
timestamp 1644511149
transform 1 0 111780 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1205
timestamp 1644511149
transform 1 0 111964 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1217
timestamp 1644511149
transform 1 0 113068 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1229
timestamp 1644511149
transform 1 0 114172 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1241
timestamp 1644511149
transform 1 0 115276 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_1253
timestamp 1644511149
transform 1 0 116380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1259
timestamp 1644511149
transform 1 0 116932 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_1261
timestamp 1644511149
transform 1 0 117116 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_1273
timestamp 1644511149
transform 1 0 118220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1644511149
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_181
timestamp 1644511149
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_205
timestamp 1644511149
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1644511149
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1644511149
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1644511149
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_305
timestamp 1644511149
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1644511149
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_361
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_373
timestamp 1644511149
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1644511149
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1644511149
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_505
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_517
timestamp 1644511149
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_529
timestamp 1644511149
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_541
timestamp 1644511149
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1644511149
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1644511149
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_573
timestamp 1644511149
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_585
timestamp 1644511149
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_597
timestamp 1644511149
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1644511149
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1644511149
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_629
timestamp 1644511149
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_641
timestamp 1644511149
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_653
timestamp 1644511149
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1644511149
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1644511149
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_673
timestamp 1644511149
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_685
timestamp 1644511149
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_697
timestamp 1644511149
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_709
timestamp 1644511149
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1644511149
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1644511149
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_729
timestamp 1644511149
transform 1 0 68172 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_741
timestamp 1644511149
transform 1 0 69276 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_753
timestamp 1644511149
transform 1 0 70380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_765
timestamp 1644511149
transform 1 0 71484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 1644511149
transform 1 0 72588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 1644511149
transform 1 0 73140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_785
timestamp 1644511149
transform 1 0 73324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_797
timestamp 1644511149
transform 1 0 74428 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_809
timestamp 1644511149
transform 1 0 75532 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_821
timestamp 1644511149
transform 1 0 76636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_833
timestamp 1644511149
transform 1 0 77740 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_839
timestamp 1644511149
transform 1 0 78292 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_841
timestamp 1644511149
transform 1 0 78476 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_853
timestamp 1644511149
transform 1 0 79580 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_865
timestamp 1644511149
transform 1 0 80684 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_877
timestamp 1644511149
transform 1 0 81788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_889
timestamp 1644511149
transform 1 0 82892 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_895
timestamp 1644511149
transform 1 0 83444 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_897
timestamp 1644511149
transform 1 0 83628 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_909
timestamp 1644511149
transform 1 0 84732 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_921
timestamp 1644511149
transform 1 0 85836 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_933
timestamp 1644511149
transform 1 0 86940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_945
timestamp 1644511149
transform 1 0 88044 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_951
timestamp 1644511149
transform 1 0 88596 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_953
timestamp 1644511149
transform 1 0 88780 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_965
timestamp 1644511149
transform 1 0 89884 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_977
timestamp 1644511149
transform 1 0 90988 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_989
timestamp 1644511149
transform 1 0 92092 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1001
timestamp 1644511149
transform 1 0 93196 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1007
timestamp 1644511149
transform 1 0 93748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1009
timestamp 1644511149
transform 1 0 93932 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1021
timestamp 1644511149
transform 1 0 95036 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1033
timestamp 1644511149
transform 1 0 96140 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1045
timestamp 1644511149
transform 1 0 97244 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1057
timestamp 1644511149
transform 1 0 98348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1063
timestamp 1644511149
transform 1 0 98900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1065
timestamp 1644511149
transform 1 0 99084 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1077
timestamp 1644511149
transform 1 0 100188 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1089
timestamp 1644511149
transform 1 0 101292 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1101
timestamp 1644511149
transform 1 0 102396 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1113
timestamp 1644511149
transform 1 0 103500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1119
timestamp 1644511149
transform 1 0 104052 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1121
timestamp 1644511149
transform 1 0 104236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1133
timestamp 1644511149
transform 1 0 105340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1145
timestamp 1644511149
transform 1 0 106444 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1157
timestamp 1644511149
transform 1 0 107548 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1169
timestamp 1644511149
transform 1 0 108652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1175
timestamp 1644511149
transform 1 0 109204 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1177
timestamp 1644511149
transform 1 0 109388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1189
timestamp 1644511149
transform 1 0 110492 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1201
timestamp 1644511149
transform 1 0 111596 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1213
timestamp 1644511149
transform 1 0 112700 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_1225
timestamp 1644511149
transform 1 0 113804 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_1231
timestamp 1644511149
transform 1 0 114356 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1233
timestamp 1644511149
transform 1 0 114540 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_1245
timestamp 1644511149
transform 1 0 115644 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_1257
timestamp 1644511149
transform 1 0 116748 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_1267
timestamp 1644511149
transform 1 0 117668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_1273
timestamp 1644511149
transform 1 0 118220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1644511149
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1644511149
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_209
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_221
timestamp 1644511149
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1644511149
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1644511149
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1644511149
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1644511149
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_389
timestamp 1644511149
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_401
timestamp 1644511149
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1644511149
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1644511149
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_501
timestamp 1644511149
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_513
timestamp 1644511149
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1644511149
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1644511149
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_533
timestamp 1644511149
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_545
timestamp 1644511149
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_557
timestamp 1644511149
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_569
timestamp 1644511149
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1644511149
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_613
timestamp 1644511149
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_625
timestamp 1644511149
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1644511149
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1644511149
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_645
timestamp 1644511149
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_657
timestamp 1644511149
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_669
timestamp 1644511149
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_681
timestamp 1644511149
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1644511149
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1644511149
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_701
timestamp 1644511149
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_713
timestamp 1644511149
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_725
timestamp 1644511149
transform 1 0 67804 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_737
timestamp 1644511149
transform 1 0 68908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 1644511149
transform 1 0 70012 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 1644511149
transform 1 0 70564 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_757
timestamp 1644511149
transform 1 0 70748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_769
timestamp 1644511149
transform 1 0 71852 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_781
timestamp 1644511149
transform 1 0 72956 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_793
timestamp 1644511149
transform 1 0 74060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 1644511149
transform 1 0 75164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 1644511149
transform 1 0 75716 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_813
timestamp 1644511149
transform 1 0 75900 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_825
timestamp 1644511149
transform 1 0 77004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_837
timestamp 1644511149
transform 1 0 78108 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_849
timestamp 1644511149
transform 1 0 79212 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_861
timestamp 1644511149
transform 1 0 80316 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_867
timestamp 1644511149
transform 1 0 80868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_869
timestamp 1644511149
transform 1 0 81052 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_881
timestamp 1644511149
transform 1 0 82156 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_893
timestamp 1644511149
transform 1 0 83260 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_905
timestamp 1644511149
transform 1 0 84364 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_917
timestamp 1644511149
transform 1 0 85468 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_923
timestamp 1644511149
transform 1 0 86020 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_925
timestamp 1644511149
transform 1 0 86204 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_937
timestamp 1644511149
transform 1 0 87308 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_949
timestamp 1644511149
transform 1 0 88412 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_961
timestamp 1644511149
transform 1 0 89516 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_973
timestamp 1644511149
transform 1 0 90620 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_979
timestamp 1644511149
transform 1 0 91172 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_981
timestamp 1644511149
transform 1 0 91356 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_993
timestamp 1644511149
transform 1 0 92460 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1005
timestamp 1644511149
transform 1 0 93564 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1017
timestamp 1644511149
transform 1 0 94668 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1029
timestamp 1644511149
transform 1 0 95772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1035
timestamp 1644511149
transform 1 0 96324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1037
timestamp 1644511149
transform 1 0 96508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1049
timestamp 1644511149
transform 1 0 97612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1061
timestamp 1644511149
transform 1 0 98716 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1073
timestamp 1644511149
transform 1 0 99820 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1085
timestamp 1644511149
transform 1 0 100924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1091
timestamp 1644511149
transform 1 0 101476 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1093
timestamp 1644511149
transform 1 0 101660 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1105
timestamp 1644511149
transform 1 0 102764 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1117
timestamp 1644511149
transform 1 0 103868 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1129
timestamp 1644511149
transform 1 0 104972 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1141
timestamp 1644511149
transform 1 0 106076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1147
timestamp 1644511149
transform 1 0 106628 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1149
timestamp 1644511149
transform 1 0 106812 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1161
timestamp 1644511149
transform 1 0 107916 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1173
timestamp 1644511149
transform 1 0 109020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1185
timestamp 1644511149
transform 1 0 110124 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1197
timestamp 1644511149
transform 1 0 111228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1203
timestamp 1644511149
transform 1 0 111780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1205
timestamp 1644511149
transform 1 0 111964 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1217
timestamp 1644511149
transform 1 0 113068 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1229
timestamp 1644511149
transform 1 0 114172 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1241
timestamp 1644511149
transform 1 0 115276 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_1253
timestamp 1644511149
transform 1 0 116380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_1259
timestamp 1644511149
transform 1 0 116932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_1261
timestamp 1644511149
transform 1 0 117116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_1273
timestamp 1644511149
transform 1 0 118220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1644511149
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1644511149
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_193
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_205
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_249
timestamp 1644511149
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_261
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_305
timestamp 1644511149
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_349
timestamp 1644511149
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_361
timestamp 1644511149
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_373
timestamp 1644511149
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1644511149
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1644511149
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1644511149
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1644511149
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1644511149
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_629
timestamp 1644511149
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_641
timestamp 1644511149
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_653
timestamp 1644511149
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1644511149
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1644511149
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_673
timestamp 1644511149
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_685
timestamp 1644511149
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_697
timestamp 1644511149
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_709
timestamp 1644511149
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1644511149
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1644511149
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_729
timestamp 1644511149
transform 1 0 68172 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_741
timestamp 1644511149
transform 1 0 69276 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_753
timestamp 1644511149
transform 1 0 70380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_765
timestamp 1644511149
transform 1 0 71484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_777
timestamp 1644511149
transform 1 0 72588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_783
timestamp 1644511149
transform 1 0 73140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_785
timestamp 1644511149
transform 1 0 73324 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_797
timestamp 1644511149
transform 1 0 74428 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_809
timestamp 1644511149
transform 1 0 75532 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_821
timestamp 1644511149
transform 1 0 76636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_833
timestamp 1644511149
transform 1 0 77740 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_839
timestamp 1644511149
transform 1 0 78292 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_841
timestamp 1644511149
transform 1 0 78476 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_853
timestamp 1644511149
transform 1 0 79580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_865
timestamp 1644511149
transform 1 0 80684 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_877
timestamp 1644511149
transform 1 0 81788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_889
timestamp 1644511149
transform 1 0 82892 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_895
timestamp 1644511149
transform 1 0 83444 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_897
timestamp 1644511149
transform 1 0 83628 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_909
timestamp 1644511149
transform 1 0 84732 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_921
timestamp 1644511149
transform 1 0 85836 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_933
timestamp 1644511149
transform 1 0 86940 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_945
timestamp 1644511149
transform 1 0 88044 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_951
timestamp 1644511149
transform 1 0 88596 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_953
timestamp 1644511149
transform 1 0 88780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_965
timestamp 1644511149
transform 1 0 89884 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_977
timestamp 1644511149
transform 1 0 90988 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_989
timestamp 1644511149
transform 1 0 92092 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1001
timestamp 1644511149
transform 1 0 93196 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1007
timestamp 1644511149
transform 1 0 93748 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1009
timestamp 1644511149
transform 1 0 93932 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1021
timestamp 1644511149
transform 1 0 95036 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1033
timestamp 1644511149
transform 1 0 96140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1045
timestamp 1644511149
transform 1 0 97244 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1057
timestamp 1644511149
transform 1 0 98348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1063
timestamp 1644511149
transform 1 0 98900 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1065
timestamp 1644511149
transform 1 0 99084 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1077
timestamp 1644511149
transform 1 0 100188 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1089
timestamp 1644511149
transform 1 0 101292 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1101
timestamp 1644511149
transform 1 0 102396 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1113
timestamp 1644511149
transform 1 0 103500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1119
timestamp 1644511149
transform 1 0 104052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1121
timestamp 1644511149
transform 1 0 104236 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1133
timestamp 1644511149
transform 1 0 105340 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1145
timestamp 1644511149
transform 1 0 106444 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1157
timestamp 1644511149
transform 1 0 107548 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1169
timestamp 1644511149
transform 1 0 108652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1175
timestamp 1644511149
transform 1 0 109204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1177
timestamp 1644511149
transform 1 0 109388 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1189
timestamp 1644511149
transform 1 0 110492 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1201
timestamp 1644511149
transform 1 0 111596 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1213
timestamp 1644511149
transform 1 0 112700 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_1225
timestamp 1644511149
transform 1 0 113804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1231
timestamp 1644511149
transform 1 0 114356 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1233
timestamp 1644511149
transform 1 0 114540 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_1245
timestamp 1644511149
transform 1 0 115644 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_1257
timestamp 1644511149
transform 1 0 116748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_1267
timestamp 1644511149
transform 1 0 117668 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_1273
timestamp 1644511149
transform 1 0 118220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_165
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_177
timestamp 1644511149
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1644511149
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_221
timestamp 1644511149
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_233
timestamp 1644511149
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1644511149
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_277
timestamp 1644511149
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_289
timestamp 1644511149
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_333
timestamp 1644511149
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1644511149
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1644511149
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1644511149
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1644511149
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_545
timestamp 1644511149
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_557
timestamp 1644511149
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_569
timestamp 1644511149
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1644511149
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_601
timestamp 1644511149
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_613
timestamp 1644511149
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_625
timestamp 1644511149
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1644511149
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1644511149
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_645
timestamp 1644511149
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_657
timestamp 1644511149
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_669
timestamp 1644511149
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_681
timestamp 1644511149
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1644511149
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1644511149
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_701
timestamp 1644511149
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_713
timestamp 1644511149
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_725
timestamp 1644511149
transform 1 0 67804 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_737
timestamp 1644511149
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 1644511149
transform 1 0 70012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 1644511149
transform 1 0 70564 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_757
timestamp 1644511149
transform 1 0 70748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_769
timestamp 1644511149
transform 1 0 71852 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_781
timestamp 1644511149
transform 1 0 72956 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_793
timestamp 1644511149
transform 1 0 74060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 1644511149
transform 1 0 75164 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 1644511149
transform 1 0 75716 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_813
timestamp 1644511149
transform 1 0 75900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_825
timestamp 1644511149
transform 1 0 77004 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_837
timestamp 1644511149
transform 1 0 78108 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_849
timestamp 1644511149
transform 1 0 79212 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_861
timestamp 1644511149
transform 1 0 80316 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_867
timestamp 1644511149
transform 1 0 80868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_869
timestamp 1644511149
transform 1 0 81052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_881
timestamp 1644511149
transform 1 0 82156 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_893
timestamp 1644511149
transform 1 0 83260 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_905
timestamp 1644511149
transform 1 0 84364 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_917
timestamp 1644511149
transform 1 0 85468 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_923
timestamp 1644511149
transform 1 0 86020 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_925
timestamp 1644511149
transform 1 0 86204 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_937
timestamp 1644511149
transform 1 0 87308 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_949
timestamp 1644511149
transform 1 0 88412 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_961
timestamp 1644511149
transform 1 0 89516 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_973
timestamp 1644511149
transform 1 0 90620 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_979
timestamp 1644511149
transform 1 0 91172 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_981
timestamp 1644511149
transform 1 0 91356 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_993
timestamp 1644511149
transform 1 0 92460 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1005
timestamp 1644511149
transform 1 0 93564 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1017
timestamp 1644511149
transform 1 0 94668 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1029
timestamp 1644511149
transform 1 0 95772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1035
timestamp 1644511149
transform 1 0 96324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1037
timestamp 1644511149
transform 1 0 96508 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1049
timestamp 1644511149
transform 1 0 97612 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1061
timestamp 1644511149
transform 1 0 98716 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1073
timestamp 1644511149
transform 1 0 99820 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1085
timestamp 1644511149
transform 1 0 100924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1091
timestamp 1644511149
transform 1 0 101476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1093
timestamp 1644511149
transform 1 0 101660 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1105
timestamp 1644511149
transform 1 0 102764 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1117
timestamp 1644511149
transform 1 0 103868 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1129
timestamp 1644511149
transform 1 0 104972 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1141
timestamp 1644511149
transform 1 0 106076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1147
timestamp 1644511149
transform 1 0 106628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1149
timestamp 1644511149
transform 1 0 106812 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1161
timestamp 1644511149
transform 1 0 107916 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1173
timestamp 1644511149
transform 1 0 109020 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1185
timestamp 1644511149
transform 1 0 110124 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1197
timestamp 1644511149
transform 1 0 111228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1203
timestamp 1644511149
transform 1 0 111780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1205
timestamp 1644511149
transform 1 0 111964 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1217
timestamp 1644511149
transform 1 0 113068 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1229
timestamp 1644511149
transform 1 0 114172 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_1241
timestamp 1644511149
transform 1 0 115276 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_1253
timestamp 1644511149
transform 1 0 116380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1259
timestamp 1644511149
transform 1 0 116932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_1261
timestamp 1644511149
transform 1 0 117116 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_1267
timestamp 1644511149
transform 1 0 117668 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_1273
timestamp 1644511149
transform 1 0 118220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1644511149
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_93
timestamp 1644511149
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_205
timestamp 1644511149
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1644511149
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1644511149
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_305
timestamp 1644511149
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_317
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_361
timestamp 1644511149
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_373
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_517
timestamp 1644511149
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_529
timestamp 1644511149
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_541
timestamp 1644511149
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1644511149
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1644511149
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_561
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_573
timestamp 1644511149
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_585
timestamp 1644511149
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_597
timestamp 1644511149
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1644511149
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1644511149
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_617
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_629
timestamp 1644511149
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_641
timestamp 1644511149
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_653
timestamp 1644511149
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1644511149
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1644511149
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_673
timestamp 1644511149
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_685
timestamp 1644511149
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_697
timestamp 1644511149
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_709
timestamp 1644511149
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1644511149
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1644511149
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_729
timestamp 1644511149
transform 1 0 68172 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_741
timestamp 1644511149
transform 1 0 69276 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_753
timestamp 1644511149
transform 1 0 70380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_765
timestamp 1644511149
transform 1 0 71484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 1644511149
transform 1 0 72588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 1644511149
transform 1 0 73140 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_785
timestamp 1644511149
transform 1 0 73324 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_797
timestamp 1644511149
transform 1 0 74428 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_809
timestamp 1644511149
transform 1 0 75532 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_821
timestamp 1644511149
transform 1 0 76636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_833
timestamp 1644511149
transform 1 0 77740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_839
timestamp 1644511149
transform 1 0 78292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_841
timestamp 1644511149
transform 1 0 78476 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_853
timestamp 1644511149
transform 1 0 79580 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_865
timestamp 1644511149
transform 1 0 80684 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_877
timestamp 1644511149
transform 1 0 81788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_889
timestamp 1644511149
transform 1 0 82892 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_895
timestamp 1644511149
transform 1 0 83444 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_897
timestamp 1644511149
transform 1 0 83628 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_909
timestamp 1644511149
transform 1 0 84732 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_921
timestamp 1644511149
transform 1 0 85836 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_933
timestamp 1644511149
transform 1 0 86940 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_945
timestamp 1644511149
transform 1 0 88044 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_951
timestamp 1644511149
transform 1 0 88596 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_953
timestamp 1644511149
transform 1 0 88780 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_965
timestamp 1644511149
transform 1 0 89884 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_977
timestamp 1644511149
transform 1 0 90988 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_989
timestamp 1644511149
transform 1 0 92092 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1001
timestamp 1644511149
transform 1 0 93196 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1007
timestamp 1644511149
transform 1 0 93748 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1009
timestamp 1644511149
transform 1 0 93932 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1021
timestamp 1644511149
transform 1 0 95036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1033
timestamp 1644511149
transform 1 0 96140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1045
timestamp 1644511149
transform 1 0 97244 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1057
timestamp 1644511149
transform 1 0 98348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1063
timestamp 1644511149
transform 1 0 98900 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1065
timestamp 1644511149
transform 1 0 99084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1077
timestamp 1644511149
transform 1 0 100188 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1089
timestamp 1644511149
transform 1 0 101292 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1101
timestamp 1644511149
transform 1 0 102396 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1113
timestamp 1644511149
transform 1 0 103500 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1119
timestamp 1644511149
transform 1 0 104052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1121
timestamp 1644511149
transform 1 0 104236 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1133
timestamp 1644511149
transform 1 0 105340 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1145
timestamp 1644511149
transform 1 0 106444 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1157
timestamp 1644511149
transform 1 0 107548 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1169
timestamp 1644511149
transform 1 0 108652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1175
timestamp 1644511149
transform 1 0 109204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1177
timestamp 1644511149
transform 1 0 109388 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1189
timestamp 1644511149
transform 1 0 110492 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1201
timestamp 1644511149
transform 1 0 111596 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1213
timestamp 1644511149
transform 1 0 112700 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_1225
timestamp 1644511149
transform 1 0 113804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1231
timestamp 1644511149
transform 1 0 114356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1233
timestamp 1644511149
transform 1 0 114540 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1245
timestamp 1644511149
transform 1 0 115644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_1257
timestamp 1644511149
transform 1 0 116748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_1269
timestamp 1644511149
transform 1 0 117852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_165
timestamp 1644511149
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_177
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_221
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_233
timestamp 1644511149
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_277
timestamp 1644511149
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_289
timestamp 1644511149
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1644511149
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1644511149
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_345
timestamp 1644511149
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1644511149
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1644511149
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_377
timestamp 1644511149
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_389
timestamp 1644511149
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_401
timestamp 1644511149
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1644511149
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1644511149
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_513
timestamp 1644511149
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1644511149
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1644511149
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_613
timestamp 1644511149
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_625
timestamp 1644511149
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1644511149
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1644511149
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_645
timestamp 1644511149
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_657
timestamp 1644511149
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_669
timestamp 1644511149
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_681
timestamp 1644511149
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1644511149
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1644511149
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_701
timestamp 1644511149
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_713
timestamp 1644511149
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_725
timestamp 1644511149
transform 1 0 67804 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_737
timestamp 1644511149
transform 1 0 68908 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 1644511149
transform 1 0 70012 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 1644511149
transform 1 0 70564 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_757
timestamp 1644511149
transform 1 0 70748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_769
timestamp 1644511149
transform 1 0 71852 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_781
timestamp 1644511149
transform 1 0 72956 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_793
timestamp 1644511149
transform 1 0 74060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 1644511149
transform 1 0 75164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 1644511149
transform 1 0 75716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_813
timestamp 1644511149
transform 1 0 75900 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_825
timestamp 1644511149
transform 1 0 77004 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_837
timestamp 1644511149
transform 1 0 78108 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_849
timestamp 1644511149
transform 1 0 79212 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_861
timestamp 1644511149
transform 1 0 80316 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_867
timestamp 1644511149
transform 1 0 80868 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_869
timestamp 1644511149
transform 1 0 81052 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_881
timestamp 1644511149
transform 1 0 82156 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_893
timestamp 1644511149
transform 1 0 83260 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_905
timestamp 1644511149
transform 1 0 84364 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_917
timestamp 1644511149
transform 1 0 85468 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_923
timestamp 1644511149
transform 1 0 86020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_925
timestamp 1644511149
transform 1 0 86204 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_937
timestamp 1644511149
transform 1 0 87308 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_949
timestamp 1644511149
transform 1 0 88412 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_961
timestamp 1644511149
transform 1 0 89516 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_973
timestamp 1644511149
transform 1 0 90620 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_979
timestamp 1644511149
transform 1 0 91172 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_981
timestamp 1644511149
transform 1 0 91356 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_993
timestamp 1644511149
transform 1 0 92460 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1005
timestamp 1644511149
transform 1 0 93564 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1017
timestamp 1644511149
transform 1 0 94668 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1029
timestamp 1644511149
transform 1 0 95772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1035
timestamp 1644511149
transform 1 0 96324 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1037
timestamp 1644511149
transform 1 0 96508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1049
timestamp 1644511149
transform 1 0 97612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1061
timestamp 1644511149
transform 1 0 98716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1073
timestamp 1644511149
transform 1 0 99820 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1085
timestamp 1644511149
transform 1 0 100924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1091
timestamp 1644511149
transform 1 0 101476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1093
timestamp 1644511149
transform 1 0 101660 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1105
timestamp 1644511149
transform 1 0 102764 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1117
timestamp 1644511149
transform 1 0 103868 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1129
timestamp 1644511149
transform 1 0 104972 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1141
timestamp 1644511149
transform 1 0 106076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1147
timestamp 1644511149
transform 1 0 106628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1149
timestamp 1644511149
transform 1 0 106812 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1161
timestamp 1644511149
transform 1 0 107916 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1173
timestamp 1644511149
transform 1 0 109020 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1185
timestamp 1644511149
transform 1 0 110124 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1197
timestamp 1644511149
transform 1 0 111228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1203
timestamp 1644511149
transform 1 0 111780 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1205
timestamp 1644511149
transform 1 0 111964 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1217
timestamp 1644511149
transform 1 0 113068 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1229
timestamp 1644511149
transform 1 0 114172 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_1241
timestamp 1644511149
transform 1 0 115276 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_1253
timestamp 1644511149
transform 1 0 116380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_1259
timestamp 1644511149
transform 1 0 116932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_1261
timestamp 1644511149
transform 1 0 117116 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_1267
timestamp 1644511149
transform 1 0 117668 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_1273
timestamp 1644511149
transform 1 0 118220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_181
timestamp 1644511149
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_205
timestamp 1644511149
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_237
timestamp 1644511149
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1644511149
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_305
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_361
timestamp 1644511149
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_373
timestamp 1644511149
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_529
timestamp 1644511149
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_541
timestamp 1644511149
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1644511149
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1644511149
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_561
timestamp 1644511149
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_573
timestamp 1644511149
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_585
timestamp 1644511149
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_597
timestamp 1644511149
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1644511149
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1644511149
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_629
timestamp 1644511149
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_641
timestamp 1644511149
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_653
timestamp 1644511149
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1644511149
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1644511149
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_673
timestamp 1644511149
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_685
timestamp 1644511149
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_697
timestamp 1644511149
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_709
timestamp 1644511149
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1644511149
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1644511149
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_729
timestamp 1644511149
transform 1 0 68172 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_741
timestamp 1644511149
transform 1 0 69276 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_753
timestamp 1644511149
transform 1 0 70380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_765
timestamp 1644511149
transform 1 0 71484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 1644511149
transform 1 0 72588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 1644511149
transform 1 0 73140 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_785
timestamp 1644511149
transform 1 0 73324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_797
timestamp 1644511149
transform 1 0 74428 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_809
timestamp 1644511149
transform 1 0 75532 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_821
timestamp 1644511149
transform 1 0 76636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_833
timestamp 1644511149
transform 1 0 77740 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_839
timestamp 1644511149
transform 1 0 78292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_841
timestamp 1644511149
transform 1 0 78476 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_853
timestamp 1644511149
transform 1 0 79580 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_865
timestamp 1644511149
transform 1 0 80684 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_877
timestamp 1644511149
transform 1 0 81788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_889
timestamp 1644511149
transform 1 0 82892 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_895
timestamp 1644511149
transform 1 0 83444 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_897
timestamp 1644511149
transform 1 0 83628 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_909
timestamp 1644511149
transform 1 0 84732 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_921
timestamp 1644511149
transform 1 0 85836 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_933
timestamp 1644511149
transform 1 0 86940 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_945
timestamp 1644511149
transform 1 0 88044 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_951
timestamp 1644511149
transform 1 0 88596 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_953
timestamp 1644511149
transform 1 0 88780 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_965
timestamp 1644511149
transform 1 0 89884 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_977
timestamp 1644511149
transform 1 0 90988 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_989
timestamp 1644511149
transform 1 0 92092 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1001
timestamp 1644511149
transform 1 0 93196 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1007
timestamp 1644511149
transform 1 0 93748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1009
timestamp 1644511149
transform 1 0 93932 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1021
timestamp 1644511149
transform 1 0 95036 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1033
timestamp 1644511149
transform 1 0 96140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1045
timestamp 1644511149
transform 1 0 97244 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1057
timestamp 1644511149
transform 1 0 98348 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1063
timestamp 1644511149
transform 1 0 98900 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1065
timestamp 1644511149
transform 1 0 99084 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1077
timestamp 1644511149
transform 1 0 100188 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1089
timestamp 1644511149
transform 1 0 101292 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1101
timestamp 1644511149
transform 1 0 102396 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1113
timestamp 1644511149
transform 1 0 103500 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1119
timestamp 1644511149
transform 1 0 104052 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1121
timestamp 1644511149
transform 1 0 104236 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1133
timestamp 1644511149
transform 1 0 105340 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1145
timestamp 1644511149
transform 1 0 106444 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1157
timestamp 1644511149
transform 1 0 107548 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1169
timestamp 1644511149
transform 1 0 108652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1175
timestamp 1644511149
transform 1 0 109204 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1177
timestamp 1644511149
transform 1 0 109388 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1189
timestamp 1644511149
transform 1 0 110492 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1201
timestamp 1644511149
transform 1 0 111596 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1213
timestamp 1644511149
transform 1 0 112700 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_1225
timestamp 1644511149
transform 1 0 113804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_1231
timestamp 1644511149
transform 1 0 114356 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1233
timestamp 1644511149
transform 1 0 114540 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1245
timestamp 1644511149
transform 1 0 115644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_1257
timestamp 1644511149
transform 1 0 116748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1269
timestamp 1644511149
transform 1 0 117852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_165
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_177
timestamp 1644511149
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1644511149
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_277
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_333
timestamp 1644511149
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_345
timestamp 1644511149
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1644511149
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1644511149
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_533
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_545
timestamp 1644511149
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_557
timestamp 1644511149
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_569
timestamp 1644511149
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1644511149
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1644511149
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_589
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_601
timestamp 1644511149
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_613
timestamp 1644511149
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_625
timestamp 1644511149
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1644511149
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1644511149
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_645
timestamp 1644511149
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_657
timestamp 1644511149
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_669
timestamp 1644511149
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_681
timestamp 1644511149
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1644511149
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1644511149
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_701
timestamp 1644511149
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_713
timestamp 1644511149
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_725
timestamp 1644511149
transform 1 0 67804 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_737
timestamp 1644511149
transform 1 0 68908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 1644511149
transform 1 0 70012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 1644511149
transform 1 0 70564 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_757
timestamp 1644511149
transform 1 0 70748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_769
timestamp 1644511149
transform 1 0 71852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_781
timestamp 1644511149
transform 1 0 72956 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_793
timestamp 1644511149
transform 1 0 74060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 1644511149
transform 1 0 75164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 1644511149
transform 1 0 75716 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_813
timestamp 1644511149
transform 1 0 75900 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_825
timestamp 1644511149
transform 1 0 77004 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_837
timestamp 1644511149
transform 1 0 78108 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_849
timestamp 1644511149
transform 1 0 79212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_861
timestamp 1644511149
transform 1 0 80316 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_867
timestamp 1644511149
transform 1 0 80868 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_869
timestamp 1644511149
transform 1 0 81052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_881
timestamp 1644511149
transform 1 0 82156 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_893
timestamp 1644511149
transform 1 0 83260 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_905
timestamp 1644511149
transform 1 0 84364 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_917
timestamp 1644511149
transform 1 0 85468 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_923
timestamp 1644511149
transform 1 0 86020 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_925
timestamp 1644511149
transform 1 0 86204 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_937
timestamp 1644511149
transform 1 0 87308 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_949
timestamp 1644511149
transform 1 0 88412 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_961
timestamp 1644511149
transform 1 0 89516 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_973
timestamp 1644511149
transform 1 0 90620 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_979
timestamp 1644511149
transform 1 0 91172 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_981
timestamp 1644511149
transform 1 0 91356 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_993
timestamp 1644511149
transform 1 0 92460 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1005
timestamp 1644511149
transform 1 0 93564 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1017
timestamp 1644511149
transform 1 0 94668 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1029
timestamp 1644511149
transform 1 0 95772 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1035
timestamp 1644511149
transform 1 0 96324 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1037
timestamp 1644511149
transform 1 0 96508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1049
timestamp 1644511149
transform 1 0 97612 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1061
timestamp 1644511149
transform 1 0 98716 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1073
timestamp 1644511149
transform 1 0 99820 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1085
timestamp 1644511149
transform 1 0 100924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1091
timestamp 1644511149
transform 1 0 101476 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1093
timestamp 1644511149
transform 1 0 101660 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1105
timestamp 1644511149
transform 1 0 102764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1117
timestamp 1644511149
transform 1 0 103868 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1129
timestamp 1644511149
transform 1 0 104972 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1141
timestamp 1644511149
transform 1 0 106076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1147
timestamp 1644511149
transform 1 0 106628 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1149
timestamp 1644511149
transform 1 0 106812 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1161
timestamp 1644511149
transform 1 0 107916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1173
timestamp 1644511149
transform 1 0 109020 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1185
timestamp 1644511149
transform 1 0 110124 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1197
timestamp 1644511149
transform 1 0 111228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1203
timestamp 1644511149
transform 1 0 111780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1205
timestamp 1644511149
transform 1 0 111964 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1217
timestamp 1644511149
transform 1 0 113068 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1229
timestamp 1644511149
transform 1 0 114172 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_1241
timestamp 1644511149
transform 1 0 115276 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_1253
timestamp 1644511149
transform 1 0 116380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1259
timestamp 1644511149
transform 1 0 116932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_1261
timestamp 1644511149
transform 1 0 117116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_1267
timestamp 1644511149
transform 1 0 117668 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_1273
timestamp 1644511149
transform 1 0 118220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_205
timestamp 1644511149
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_237
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_249
timestamp 1644511149
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_261
timestamp 1644511149
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1644511149
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_373
timestamp 1644511149
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1644511149
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_517
timestamp 1644511149
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_529
timestamp 1644511149
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_541
timestamp 1644511149
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1644511149
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_561
timestamp 1644511149
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_573
timestamp 1644511149
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_585
timestamp 1644511149
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_597
timestamp 1644511149
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1644511149
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_629
timestamp 1644511149
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_641
timestamp 1644511149
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_653
timestamp 1644511149
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1644511149
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1644511149
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_673
timestamp 1644511149
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_685
timestamp 1644511149
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_697
timestamp 1644511149
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_709
timestamp 1644511149
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1644511149
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1644511149
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_729
timestamp 1644511149
transform 1 0 68172 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_741
timestamp 1644511149
transform 1 0 69276 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_753
timestamp 1644511149
transform 1 0 70380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_765
timestamp 1644511149
transform 1 0 71484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 1644511149
transform 1 0 72588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 1644511149
transform 1 0 73140 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_785
timestamp 1644511149
transform 1 0 73324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_797
timestamp 1644511149
transform 1 0 74428 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_809
timestamp 1644511149
transform 1 0 75532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_821
timestamp 1644511149
transform 1 0 76636 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_833
timestamp 1644511149
transform 1 0 77740 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_839
timestamp 1644511149
transform 1 0 78292 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_841
timestamp 1644511149
transform 1 0 78476 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_853
timestamp 1644511149
transform 1 0 79580 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_865
timestamp 1644511149
transform 1 0 80684 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_877
timestamp 1644511149
transform 1 0 81788 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_889
timestamp 1644511149
transform 1 0 82892 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_895
timestamp 1644511149
transform 1 0 83444 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_897
timestamp 1644511149
transform 1 0 83628 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_909
timestamp 1644511149
transform 1 0 84732 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_921
timestamp 1644511149
transform 1 0 85836 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_933
timestamp 1644511149
transform 1 0 86940 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_945
timestamp 1644511149
transform 1 0 88044 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_951
timestamp 1644511149
transform 1 0 88596 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_953
timestamp 1644511149
transform 1 0 88780 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_965
timestamp 1644511149
transform 1 0 89884 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_977
timestamp 1644511149
transform 1 0 90988 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_989
timestamp 1644511149
transform 1 0 92092 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1001
timestamp 1644511149
transform 1 0 93196 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1007
timestamp 1644511149
transform 1 0 93748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1009
timestamp 1644511149
transform 1 0 93932 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1021
timestamp 1644511149
transform 1 0 95036 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1033
timestamp 1644511149
transform 1 0 96140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1045
timestamp 1644511149
transform 1 0 97244 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1057
timestamp 1644511149
transform 1 0 98348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1063
timestamp 1644511149
transform 1 0 98900 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1065
timestamp 1644511149
transform 1 0 99084 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1077
timestamp 1644511149
transform 1 0 100188 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1089
timestamp 1644511149
transform 1 0 101292 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1101
timestamp 1644511149
transform 1 0 102396 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1113
timestamp 1644511149
transform 1 0 103500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1119
timestamp 1644511149
transform 1 0 104052 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1121
timestamp 1644511149
transform 1 0 104236 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1133
timestamp 1644511149
transform 1 0 105340 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1145
timestamp 1644511149
transform 1 0 106444 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1157
timestamp 1644511149
transform 1 0 107548 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1169
timestamp 1644511149
transform 1 0 108652 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1175
timestamp 1644511149
transform 1 0 109204 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1177
timestamp 1644511149
transform 1 0 109388 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1189
timestamp 1644511149
transform 1 0 110492 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1201
timestamp 1644511149
transform 1 0 111596 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1213
timestamp 1644511149
transform 1 0 112700 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_1225
timestamp 1644511149
transform 1 0 113804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1231
timestamp 1644511149
transform 1 0 114356 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1233
timestamp 1644511149
transform 1 0 114540 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_1245
timestamp 1644511149
transform 1 0 115644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_1257
timestamp 1644511149
transform 1 0 116748 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_1267
timestamp 1644511149
transform 1 0 117668 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_1273
timestamp 1644511149
transform 1 0 118220 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_209
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_277
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_333
timestamp 1644511149
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_345
timestamp 1644511149
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_389
timestamp 1644511149
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_401
timestamp 1644511149
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1644511149
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1644511149
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_433
timestamp 1644511149
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_445
timestamp 1644511149
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_457
timestamp 1644511149
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1644511149
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_501
timestamp 1644511149
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_513
timestamp 1644511149
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1644511149
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1644511149
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_569
timestamp 1644511149
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1644511149
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1644511149
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_589
timestamp 1644511149
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_601
timestamp 1644511149
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_625
timestamp 1644511149
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1644511149
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1644511149
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_645
timestamp 1644511149
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_657
timestamp 1644511149
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_669
timestamp 1644511149
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_681
timestamp 1644511149
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1644511149
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1644511149
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_701
timestamp 1644511149
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_713
timestamp 1644511149
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_725
timestamp 1644511149
transform 1 0 67804 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_737
timestamp 1644511149
transform 1 0 68908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 1644511149
transform 1 0 70012 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 1644511149
transform 1 0 70564 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_757
timestamp 1644511149
transform 1 0 70748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_769
timestamp 1644511149
transform 1 0 71852 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_781
timestamp 1644511149
transform 1 0 72956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_793
timestamp 1644511149
transform 1 0 74060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 1644511149
transform 1 0 75164 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 1644511149
transform 1 0 75716 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_813
timestamp 1644511149
transform 1 0 75900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_825
timestamp 1644511149
transform 1 0 77004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_837
timestamp 1644511149
transform 1 0 78108 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_849
timestamp 1644511149
transform 1 0 79212 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_861
timestamp 1644511149
transform 1 0 80316 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_867
timestamp 1644511149
transform 1 0 80868 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_869
timestamp 1644511149
transform 1 0 81052 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_881
timestamp 1644511149
transform 1 0 82156 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_893
timestamp 1644511149
transform 1 0 83260 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_905
timestamp 1644511149
transform 1 0 84364 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_917
timestamp 1644511149
transform 1 0 85468 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_923
timestamp 1644511149
transform 1 0 86020 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_925
timestamp 1644511149
transform 1 0 86204 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_937
timestamp 1644511149
transform 1 0 87308 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_949
timestamp 1644511149
transform 1 0 88412 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_961
timestamp 1644511149
transform 1 0 89516 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_973
timestamp 1644511149
transform 1 0 90620 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_979
timestamp 1644511149
transform 1 0 91172 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_981
timestamp 1644511149
transform 1 0 91356 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_993
timestamp 1644511149
transform 1 0 92460 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1005
timestamp 1644511149
transform 1 0 93564 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1017
timestamp 1644511149
transform 1 0 94668 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1029
timestamp 1644511149
transform 1 0 95772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1035
timestamp 1644511149
transform 1 0 96324 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1037
timestamp 1644511149
transform 1 0 96508 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1049
timestamp 1644511149
transform 1 0 97612 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1061
timestamp 1644511149
transform 1 0 98716 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1073
timestamp 1644511149
transform 1 0 99820 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1085
timestamp 1644511149
transform 1 0 100924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1091
timestamp 1644511149
transform 1 0 101476 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1093
timestamp 1644511149
transform 1 0 101660 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1105
timestamp 1644511149
transform 1 0 102764 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1117
timestamp 1644511149
transform 1 0 103868 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1129
timestamp 1644511149
transform 1 0 104972 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1141
timestamp 1644511149
transform 1 0 106076 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1147
timestamp 1644511149
transform 1 0 106628 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1149
timestamp 1644511149
transform 1 0 106812 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1161
timestamp 1644511149
transform 1 0 107916 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1173
timestamp 1644511149
transform 1 0 109020 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1185
timestamp 1644511149
transform 1 0 110124 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1197
timestamp 1644511149
transform 1 0 111228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1203
timestamp 1644511149
transform 1 0 111780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1205
timestamp 1644511149
transform 1 0 111964 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1217
timestamp 1644511149
transform 1 0 113068 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1229
timestamp 1644511149
transform 1 0 114172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1241
timestamp 1644511149
transform 1 0 115276 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_1253
timestamp 1644511149
transform 1 0 116380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1259
timestamp 1644511149
transform 1 0 116932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_1261
timestamp 1644511149
transform 1 0 117116 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_1273
timestamp 1644511149
transform 1 0 118220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1644511149
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_249
timestamp 1644511149
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_261
timestamp 1644511149
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1644511149
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1644511149
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1644511149
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_305
timestamp 1644511149
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1644511149
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1644511149
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_349
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_361
timestamp 1644511149
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1644511149
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_405
timestamp 1644511149
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_417
timestamp 1644511149
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_429
timestamp 1644511149
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1644511149
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_529
timestamp 1644511149
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_541
timestamp 1644511149
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1644511149
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1644511149
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_597
timestamp 1644511149
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1644511149
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1644511149
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_617
timestamp 1644511149
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_629
timestamp 1644511149
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_641
timestamp 1644511149
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_653
timestamp 1644511149
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1644511149
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1644511149
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_673
timestamp 1644511149
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_685
timestamp 1644511149
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_697
timestamp 1644511149
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_709
timestamp 1644511149
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1644511149
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1644511149
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_729
timestamp 1644511149
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_741
timestamp 1644511149
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_753
timestamp 1644511149
transform 1 0 70380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_765
timestamp 1644511149
transform 1 0 71484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 1644511149
transform 1 0 72588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 1644511149
transform 1 0 73140 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_785
timestamp 1644511149
transform 1 0 73324 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_797
timestamp 1644511149
transform 1 0 74428 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_809
timestamp 1644511149
transform 1 0 75532 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_821
timestamp 1644511149
transform 1 0 76636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_833
timestamp 1644511149
transform 1 0 77740 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_839
timestamp 1644511149
transform 1 0 78292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_841
timestamp 1644511149
transform 1 0 78476 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_853
timestamp 1644511149
transform 1 0 79580 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_865
timestamp 1644511149
transform 1 0 80684 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_877
timestamp 1644511149
transform 1 0 81788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_889
timestamp 1644511149
transform 1 0 82892 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_895
timestamp 1644511149
transform 1 0 83444 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_897
timestamp 1644511149
transform 1 0 83628 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_909
timestamp 1644511149
transform 1 0 84732 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_921
timestamp 1644511149
transform 1 0 85836 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_933
timestamp 1644511149
transform 1 0 86940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_945
timestamp 1644511149
transform 1 0 88044 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_951
timestamp 1644511149
transform 1 0 88596 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_953
timestamp 1644511149
transform 1 0 88780 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_965
timestamp 1644511149
transform 1 0 89884 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_977
timestamp 1644511149
transform 1 0 90988 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_989
timestamp 1644511149
transform 1 0 92092 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1001
timestamp 1644511149
transform 1 0 93196 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1007
timestamp 1644511149
transform 1 0 93748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1009
timestamp 1644511149
transform 1 0 93932 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1021
timestamp 1644511149
transform 1 0 95036 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1033
timestamp 1644511149
transform 1 0 96140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1045
timestamp 1644511149
transform 1 0 97244 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1057
timestamp 1644511149
transform 1 0 98348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1063
timestamp 1644511149
transform 1 0 98900 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1065
timestamp 1644511149
transform 1 0 99084 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1077
timestamp 1644511149
transform 1 0 100188 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1089
timestamp 1644511149
transform 1 0 101292 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1101
timestamp 1644511149
transform 1 0 102396 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1113
timestamp 1644511149
transform 1 0 103500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1119
timestamp 1644511149
transform 1 0 104052 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1121
timestamp 1644511149
transform 1 0 104236 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1133
timestamp 1644511149
transform 1 0 105340 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1145
timestamp 1644511149
transform 1 0 106444 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1157
timestamp 1644511149
transform 1 0 107548 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1169
timestamp 1644511149
transform 1 0 108652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1175
timestamp 1644511149
transform 1 0 109204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1177
timestamp 1644511149
transform 1 0 109388 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1189
timestamp 1644511149
transform 1 0 110492 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1201
timestamp 1644511149
transform 1 0 111596 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1213
timestamp 1644511149
transform 1 0 112700 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_1225
timestamp 1644511149
transform 1 0 113804 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1231
timestamp 1644511149
transform 1 0 114356 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1233
timestamp 1644511149
transform 1 0 114540 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_1245
timestamp 1644511149
transform 1 0 115644 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_1257
timestamp 1644511149
transform 1 0 116748 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_1267
timestamp 1644511149
transform 1 0 117668 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_1273
timestamp 1644511149
transform 1 0 118220 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_177
timestamp 1644511149
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1644511149
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_233
timestamp 1644511149
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_277
timestamp 1644511149
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_289
timestamp 1644511149
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1644511149
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_345
timestamp 1644511149
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_365
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_377
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_389
timestamp 1644511149
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_401
timestamp 1644511149
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1644511149
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_513
timestamp 1644511149
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1644511149
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1644511149
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_533
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_545
timestamp 1644511149
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_557
timestamp 1644511149
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_569
timestamp 1644511149
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1644511149
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_601
timestamp 1644511149
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_613
timestamp 1644511149
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_625
timestamp 1644511149
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1644511149
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1644511149
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_645
timestamp 1644511149
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_657
timestamp 1644511149
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_669
timestamp 1644511149
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_681
timestamp 1644511149
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1644511149
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1644511149
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_701
timestamp 1644511149
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_713
timestamp 1644511149
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_725
timestamp 1644511149
transform 1 0 67804 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_737
timestamp 1644511149
transform 1 0 68908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 1644511149
transform 1 0 70012 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 1644511149
transform 1 0 70564 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_757
timestamp 1644511149
transform 1 0 70748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_769
timestamp 1644511149
transform 1 0 71852 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_781
timestamp 1644511149
transform 1 0 72956 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_793
timestamp 1644511149
transform 1 0 74060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 1644511149
transform 1 0 75164 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 1644511149
transform 1 0 75716 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_813
timestamp 1644511149
transform 1 0 75900 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_825
timestamp 1644511149
transform 1 0 77004 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_837
timestamp 1644511149
transform 1 0 78108 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_849
timestamp 1644511149
transform 1 0 79212 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_861
timestamp 1644511149
transform 1 0 80316 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_867
timestamp 1644511149
transform 1 0 80868 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_869
timestamp 1644511149
transform 1 0 81052 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_881
timestamp 1644511149
transform 1 0 82156 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_893
timestamp 1644511149
transform 1 0 83260 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_905
timestamp 1644511149
transform 1 0 84364 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_917
timestamp 1644511149
transform 1 0 85468 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_923
timestamp 1644511149
transform 1 0 86020 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_925
timestamp 1644511149
transform 1 0 86204 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_937
timestamp 1644511149
transform 1 0 87308 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_949
timestamp 1644511149
transform 1 0 88412 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_961
timestamp 1644511149
transform 1 0 89516 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_973
timestamp 1644511149
transform 1 0 90620 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_979
timestamp 1644511149
transform 1 0 91172 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_981
timestamp 1644511149
transform 1 0 91356 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_993
timestamp 1644511149
transform 1 0 92460 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1005
timestamp 1644511149
transform 1 0 93564 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1017
timestamp 1644511149
transform 1 0 94668 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1029
timestamp 1644511149
transform 1 0 95772 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1035
timestamp 1644511149
transform 1 0 96324 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1037
timestamp 1644511149
transform 1 0 96508 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1049
timestamp 1644511149
transform 1 0 97612 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1061
timestamp 1644511149
transform 1 0 98716 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1073
timestamp 1644511149
transform 1 0 99820 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1085
timestamp 1644511149
transform 1 0 100924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1091
timestamp 1644511149
transform 1 0 101476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1093
timestamp 1644511149
transform 1 0 101660 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1105
timestamp 1644511149
transform 1 0 102764 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1117
timestamp 1644511149
transform 1 0 103868 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1129
timestamp 1644511149
transform 1 0 104972 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1141
timestamp 1644511149
transform 1 0 106076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1147
timestamp 1644511149
transform 1 0 106628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1149
timestamp 1644511149
transform 1 0 106812 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1161
timestamp 1644511149
transform 1 0 107916 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1173
timestamp 1644511149
transform 1 0 109020 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1185
timestamp 1644511149
transform 1 0 110124 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1197
timestamp 1644511149
transform 1 0 111228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1203
timestamp 1644511149
transform 1 0 111780 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1205
timestamp 1644511149
transform 1 0 111964 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1217
timestamp 1644511149
transform 1 0 113068 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1229
timestamp 1644511149
transform 1 0 114172 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1241
timestamp 1644511149
transform 1 0 115276 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_1253
timestamp 1644511149
transform 1 0 116380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_1259
timestamp 1644511149
transform 1 0 116932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_1261
timestamp 1644511149
transform 1 0 117116 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_1273
timestamp 1644511149
transform 1 0 118220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1644511149
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1644511149
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_261
timestamp 1644511149
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1644511149
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_305
timestamp 1644511149
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_317
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_517
timestamp 1644511149
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_529
timestamp 1644511149
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_541
timestamp 1644511149
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1644511149
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1644511149
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_561
timestamp 1644511149
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_573
timestamp 1644511149
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_585
timestamp 1644511149
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_597
timestamp 1644511149
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1644511149
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1644511149
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_629
timestamp 1644511149
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_641
timestamp 1644511149
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_653
timestamp 1644511149
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1644511149
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1644511149
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_673
timestamp 1644511149
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_685
timestamp 1644511149
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_697
timestamp 1644511149
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_709
timestamp 1644511149
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1644511149
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1644511149
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_729
timestamp 1644511149
transform 1 0 68172 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_741
timestamp 1644511149
transform 1 0 69276 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_753
timestamp 1644511149
transform 1 0 70380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_765
timestamp 1644511149
transform 1 0 71484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 1644511149
transform 1 0 72588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 1644511149
transform 1 0 73140 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_785
timestamp 1644511149
transform 1 0 73324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_797
timestamp 1644511149
transform 1 0 74428 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_809
timestamp 1644511149
transform 1 0 75532 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_821
timestamp 1644511149
transform 1 0 76636 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_833
timestamp 1644511149
transform 1 0 77740 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_839
timestamp 1644511149
transform 1 0 78292 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_841
timestamp 1644511149
transform 1 0 78476 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_853
timestamp 1644511149
transform 1 0 79580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_865
timestamp 1644511149
transform 1 0 80684 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_877
timestamp 1644511149
transform 1 0 81788 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_889
timestamp 1644511149
transform 1 0 82892 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_895
timestamp 1644511149
transform 1 0 83444 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_897
timestamp 1644511149
transform 1 0 83628 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_909
timestamp 1644511149
transform 1 0 84732 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_921
timestamp 1644511149
transform 1 0 85836 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_933
timestamp 1644511149
transform 1 0 86940 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_945
timestamp 1644511149
transform 1 0 88044 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_951
timestamp 1644511149
transform 1 0 88596 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_953
timestamp 1644511149
transform 1 0 88780 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_965
timestamp 1644511149
transform 1 0 89884 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_977
timestamp 1644511149
transform 1 0 90988 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_989
timestamp 1644511149
transform 1 0 92092 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1001
timestamp 1644511149
transform 1 0 93196 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1007
timestamp 1644511149
transform 1 0 93748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1009
timestamp 1644511149
transform 1 0 93932 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1021
timestamp 1644511149
transform 1 0 95036 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1033
timestamp 1644511149
transform 1 0 96140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1045
timestamp 1644511149
transform 1 0 97244 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1057
timestamp 1644511149
transform 1 0 98348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1063
timestamp 1644511149
transform 1 0 98900 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1065
timestamp 1644511149
transform 1 0 99084 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1077
timestamp 1644511149
transform 1 0 100188 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1089
timestamp 1644511149
transform 1 0 101292 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1101
timestamp 1644511149
transform 1 0 102396 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1113
timestamp 1644511149
transform 1 0 103500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1119
timestamp 1644511149
transform 1 0 104052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1121
timestamp 1644511149
transform 1 0 104236 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1133
timestamp 1644511149
transform 1 0 105340 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1145
timestamp 1644511149
transform 1 0 106444 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1157
timestamp 1644511149
transform 1 0 107548 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1169
timestamp 1644511149
transform 1 0 108652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1175
timestamp 1644511149
transform 1 0 109204 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1177
timestamp 1644511149
transform 1 0 109388 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1189
timestamp 1644511149
transform 1 0 110492 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1201
timestamp 1644511149
transform 1 0 111596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1213
timestamp 1644511149
transform 1 0 112700 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_1225
timestamp 1644511149
transform 1 0 113804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1231
timestamp 1644511149
transform 1 0 114356 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1233
timestamp 1644511149
transform 1 0 114540 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_1245
timestamp 1644511149
transform 1 0 115644 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1257
timestamp 1644511149
transform 1 0 116748 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_1267
timestamp 1644511149
transform 1 0 117668 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_1273
timestamp 1644511149
transform 1 0 118220 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_165
timestamp 1644511149
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1644511149
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_221
timestamp 1644511149
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_233
timestamp 1644511149
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1644511149
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1644511149
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_277
timestamp 1644511149
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_289
timestamp 1644511149
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1644511149
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_321
timestamp 1644511149
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_333
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_345
timestamp 1644511149
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1644511149
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1644511149
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_365
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_377
timestamp 1644511149
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_389
timestamp 1644511149
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_401
timestamp 1644511149
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1644511149
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_533
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_545
timestamp 1644511149
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_557
timestamp 1644511149
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_569
timestamp 1644511149
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1644511149
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1644511149
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_601
timestamp 1644511149
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_613
timestamp 1644511149
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_625
timestamp 1644511149
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1644511149
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1644511149
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_645
timestamp 1644511149
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_657
timestamp 1644511149
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_669
timestamp 1644511149
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_681
timestamp 1644511149
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1644511149
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1644511149
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_701
timestamp 1644511149
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_713
timestamp 1644511149
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_725
timestamp 1644511149
transform 1 0 67804 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_737
timestamp 1644511149
transform 1 0 68908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 1644511149
transform 1 0 70012 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 1644511149
transform 1 0 70564 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_757
timestamp 1644511149
transform 1 0 70748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_769
timestamp 1644511149
transform 1 0 71852 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_781
timestamp 1644511149
transform 1 0 72956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_793
timestamp 1644511149
transform 1 0 74060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 1644511149
transform 1 0 75164 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 1644511149
transform 1 0 75716 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_813
timestamp 1644511149
transform 1 0 75900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_825
timestamp 1644511149
transform 1 0 77004 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_837
timestamp 1644511149
transform 1 0 78108 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_849
timestamp 1644511149
transform 1 0 79212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_861
timestamp 1644511149
transform 1 0 80316 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_867
timestamp 1644511149
transform 1 0 80868 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_869
timestamp 1644511149
transform 1 0 81052 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_881
timestamp 1644511149
transform 1 0 82156 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_893
timestamp 1644511149
transform 1 0 83260 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_905
timestamp 1644511149
transform 1 0 84364 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_917
timestamp 1644511149
transform 1 0 85468 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_923
timestamp 1644511149
transform 1 0 86020 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_925
timestamp 1644511149
transform 1 0 86204 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_937
timestamp 1644511149
transform 1 0 87308 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_949
timestamp 1644511149
transform 1 0 88412 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_961
timestamp 1644511149
transform 1 0 89516 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_973
timestamp 1644511149
transform 1 0 90620 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_979
timestamp 1644511149
transform 1 0 91172 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_981
timestamp 1644511149
transform 1 0 91356 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_993
timestamp 1644511149
transform 1 0 92460 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1005
timestamp 1644511149
transform 1 0 93564 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1017
timestamp 1644511149
transform 1 0 94668 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1029
timestamp 1644511149
transform 1 0 95772 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1035
timestamp 1644511149
transform 1 0 96324 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1037
timestamp 1644511149
transform 1 0 96508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1049
timestamp 1644511149
transform 1 0 97612 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1061
timestamp 1644511149
transform 1 0 98716 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1073
timestamp 1644511149
transform 1 0 99820 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1085
timestamp 1644511149
transform 1 0 100924 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1091
timestamp 1644511149
transform 1 0 101476 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1093
timestamp 1644511149
transform 1 0 101660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1105
timestamp 1644511149
transform 1 0 102764 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1117
timestamp 1644511149
transform 1 0 103868 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1129
timestamp 1644511149
transform 1 0 104972 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1141
timestamp 1644511149
transform 1 0 106076 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1147
timestamp 1644511149
transform 1 0 106628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1149
timestamp 1644511149
transform 1 0 106812 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1161
timestamp 1644511149
transform 1 0 107916 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1173
timestamp 1644511149
transform 1 0 109020 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1185
timestamp 1644511149
transform 1 0 110124 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1197
timestamp 1644511149
transform 1 0 111228 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1203
timestamp 1644511149
transform 1 0 111780 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1205
timestamp 1644511149
transform 1 0 111964 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1217
timestamp 1644511149
transform 1 0 113068 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1229
timestamp 1644511149
transform 1 0 114172 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1241
timestamp 1644511149
transform 1 0 115276 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_1253
timestamp 1644511149
transform 1 0 116380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_1259
timestamp 1644511149
transform 1 0 116932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_1261
timestamp 1644511149
transform 1 0 117116 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_1273
timestamp 1644511149
transform 1 0 118220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_237
timestamp 1644511149
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_261
timestamp 1644511149
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_305
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_417
timestamp 1644511149
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1644511149
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_541
timestamp 1644511149
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1644511149
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1644511149
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1644511149
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1644511149
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_629
timestamp 1644511149
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_641
timestamp 1644511149
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_653
timestamp 1644511149
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1644511149
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1644511149
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_673
timestamp 1644511149
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_685
timestamp 1644511149
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_697
timestamp 1644511149
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_709
timestamp 1644511149
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1644511149
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1644511149
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_729
timestamp 1644511149
transform 1 0 68172 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_741
timestamp 1644511149
transform 1 0 69276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_753
timestamp 1644511149
transform 1 0 70380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_765
timestamp 1644511149
transform 1 0 71484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 1644511149
transform 1 0 72588 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 1644511149
transform 1 0 73140 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_785
timestamp 1644511149
transform 1 0 73324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_797
timestamp 1644511149
transform 1 0 74428 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_809
timestamp 1644511149
transform 1 0 75532 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_821
timestamp 1644511149
transform 1 0 76636 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_833
timestamp 1644511149
transform 1 0 77740 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_839
timestamp 1644511149
transform 1 0 78292 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_841
timestamp 1644511149
transform 1 0 78476 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_853
timestamp 1644511149
transform 1 0 79580 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_865
timestamp 1644511149
transform 1 0 80684 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_877
timestamp 1644511149
transform 1 0 81788 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_889
timestamp 1644511149
transform 1 0 82892 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_895
timestamp 1644511149
transform 1 0 83444 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_897
timestamp 1644511149
transform 1 0 83628 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_909
timestamp 1644511149
transform 1 0 84732 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_921
timestamp 1644511149
transform 1 0 85836 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_933
timestamp 1644511149
transform 1 0 86940 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_945
timestamp 1644511149
transform 1 0 88044 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_951
timestamp 1644511149
transform 1 0 88596 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_953
timestamp 1644511149
transform 1 0 88780 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_965
timestamp 1644511149
transform 1 0 89884 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_977
timestamp 1644511149
transform 1 0 90988 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_989
timestamp 1644511149
transform 1 0 92092 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1001
timestamp 1644511149
transform 1 0 93196 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1007
timestamp 1644511149
transform 1 0 93748 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1009
timestamp 1644511149
transform 1 0 93932 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1021
timestamp 1644511149
transform 1 0 95036 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1033
timestamp 1644511149
transform 1 0 96140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1045
timestamp 1644511149
transform 1 0 97244 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1057
timestamp 1644511149
transform 1 0 98348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1063
timestamp 1644511149
transform 1 0 98900 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1065
timestamp 1644511149
transform 1 0 99084 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1077
timestamp 1644511149
transform 1 0 100188 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1089
timestamp 1644511149
transform 1 0 101292 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1101
timestamp 1644511149
transform 1 0 102396 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1113
timestamp 1644511149
transform 1 0 103500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1119
timestamp 1644511149
transform 1 0 104052 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1121
timestamp 1644511149
transform 1 0 104236 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1133
timestamp 1644511149
transform 1 0 105340 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1145
timestamp 1644511149
transform 1 0 106444 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1157
timestamp 1644511149
transform 1 0 107548 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1169
timestamp 1644511149
transform 1 0 108652 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1175
timestamp 1644511149
transform 1 0 109204 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1177
timestamp 1644511149
transform 1 0 109388 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1189
timestamp 1644511149
transform 1 0 110492 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1201
timestamp 1644511149
transform 1 0 111596 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1213
timestamp 1644511149
transform 1 0 112700 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_1225
timestamp 1644511149
transform 1 0 113804 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1231
timestamp 1644511149
transform 1 0 114356 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1233
timestamp 1644511149
transform 1 0 114540 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1245
timestamp 1644511149
transform 1 0 115644 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_1257
timestamp 1644511149
transform 1 0 116748 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_1273
timestamp 1644511149
transform 1 0 118220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_165
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1644511149
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1644511149
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_221
timestamp 1644511149
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_233
timestamp 1644511149
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_321
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_333
timestamp 1644511149
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_345
timestamp 1644511149
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_389
timestamp 1644511149
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1644511149
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1644511149
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_545
timestamp 1644511149
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_557
timestamp 1644511149
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_569
timestamp 1644511149
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1644511149
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1644511149
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_589
timestamp 1644511149
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_601
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_613
timestamp 1644511149
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_625
timestamp 1644511149
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1644511149
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1644511149
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_645
timestamp 1644511149
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_657
timestamp 1644511149
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_669
timestamp 1644511149
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_681
timestamp 1644511149
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1644511149
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1644511149
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_701
timestamp 1644511149
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_713
timestamp 1644511149
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_725
timestamp 1644511149
transform 1 0 67804 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_737
timestamp 1644511149
transform 1 0 68908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_749
timestamp 1644511149
transform 1 0 70012 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_755
timestamp 1644511149
transform 1 0 70564 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_757
timestamp 1644511149
transform 1 0 70748 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_769
timestamp 1644511149
transform 1 0 71852 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_781
timestamp 1644511149
transform 1 0 72956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_793
timestamp 1644511149
transform 1 0 74060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_805
timestamp 1644511149
transform 1 0 75164 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_811
timestamp 1644511149
transform 1 0 75716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_813
timestamp 1644511149
transform 1 0 75900 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_825
timestamp 1644511149
transform 1 0 77004 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_837
timestamp 1644511149
transform 1 0 78108 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_849
timestamp 1644511149
transform 1 0 79212 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_861
timestamp 1644511149
transform 1 0 80316 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_867
timestamp 1644511149
transform 1 0 80868 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_869
timestamp 1644511149
transform 1 0 81052 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_881
timestamp 1644511149
transform 1 0 82156 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_893
timestamp 1644511149
transform 1 0 83260 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_905
timestamp 1644511149
transform 1 0 84364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_917
timestamp 1644511149
transform 1 0 85468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_923
timestamp 1644511149
transform 1 0 86020 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_925
timestamp 1644511149
transform 1 0 86204 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_937
timestamp 1644511149
transform 1 0 87308 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_949
timestamp 1644511149
transform 1 0 88412 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_961
timestamp 1644511149
transform 1 0 89516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_973
timestamp 1644511149
transform 1 0 90620 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_979
timestamp 1644511149
transform 1 0 91172 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_981
timestamp 1644511149
transform 1 0 91356 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_993
timestamp 1644511149
transform 1 0 92460 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1005
timestamp 1644511149
transform 1 0 93564 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1017
timestamp 1644511149
transform 1 0 94668 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1029
timestamp 1644511149
transform 1 0 95772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1035
timestamp 1644511149
transform 1 0 96324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1037
timestamp 1644511149
transform 1 0 96508 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1049
timestamp 1644511149
transform 1 0 97612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1061
timestamp 1644511149
transform 1 0 98716 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1073
timestamp 1644511149
transform 1 0 99820 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1085
timestamp 1644511149
transform 1 0 100924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1091
timestamp 1644511149
transform 1 0 101476 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1093
timestamp 1644511149
transform 1 0 101660 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1105
timestamp 1644511149
transform 1 0 102764 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1117
timestamp 1644511149
transform 1 0 103868 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1129
timestamp 1644511149
transform 1 0 104972 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1141
timestamp 1644511149
transform 1 0 106076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1147
timestamp 1644511149
transform 1 0 106628 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1149
timestamp 1644511149
transform 1 0 106812 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1161
timestamp 1644511149
transform 1 0 107916 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1173
timestamp 1644511149
transform 1 0 109020 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1185
timestamp 1644511149
transform 1 0 110124 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1197
timestamp 1644511149
transform 1 0 111228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1203
timestamp 1644511149
transform 1 0 111780 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1205
timestamp 1644511149
transform 1 0 111964 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1217
timestamp 1644511149
transform 1 0 113068 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1229
timestamp 1644511149
transform 1 0 114172 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_1241
timestamp 1644511149
transform 1 0 115276 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1253
timestamp 1644511149
transform 1 0 116380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1259
timestamp 1644511149
transform 1 0 116932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1261
timestamp 1644511149
transform 1 0 117116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_1273
timestamp 1644511149
transform 1 0 118220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_181
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_193
timestamp 1644511149
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_205
timestamp 1644511149
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1644511149
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_261
timestamp 1644511149
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1644511149
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1644511149
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1644511149
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_417
timestamp 1644511149
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_429
timestamp 1644511149
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1644511149
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1644511149
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1644511149
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_629
timestamp 1644511149
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_641
timestamp 1644511149
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_653
timestamp 1644511149
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1644511149
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1644511149
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_673
timestamp 1644511149
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_685
timestamp 1644511149
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_697
timestamp 1644511149
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_709
timestamp 1644511149
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1644511149
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1644511149
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_729
timestamp 1644511149
transform 1 0 68172 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_741
timestamp 1644511149
transform 1 0 69276 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_753
timestamp 1644511149
transform 1 0 70380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_765
timestamp 1644511149
transform 1 0 71484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_777
timestamp 1644511149
transform 1 0 72588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_783
timestamp 1644511149
transform 1 0 73140 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_785
timestamp 1644511149
transform 1 0 73324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_797
timestamp 1644511149
transform 1 0 74428 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_809
timestamp 1644511149
transform 1 0 75532 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_821
timestamp 1644511149
transform 1 0 76636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_833
timestamp 1644511149
transform 1 0 77740 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_839
timestamp 1644511149
transform 1 0 78292 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_841
timestamp 1644511149
transform 1 0 78476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_853
timestamp 1644511149
transform 1 0 79580 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_865
timestamp 1644511149
transform 1 0 80684 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_877
timestamp 1644511149
transform 1 0 81788 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_889
timestamp 1644511149
transform 1 0 82892 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_895
timestamp 1644511149
transform 1 0 83444 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_897
timestamp 1644511149
transform 1 0 83628 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_909
timestamp 1644511149
transform 1 0 84732 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_921
timestamp 1644511149
transform 1 0 85836 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_933
timestamp 1644511149
transform 1 0 86940 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_945
timestamp 1644511149
transform 1 0 88044 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_951
timestamp 1644511149
transform 1 0 88596 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_953
timestamp 1644511149
transform 1 0 88780 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_965
timestamp 1644511149
transform 1 0 89884 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_977
timestamp 1644511149
transform 1 0 90988 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_989
timestamp 1644511149
transform 1 0 92092 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1001
timestamp 1644511149
transform 1 0 93196 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1007
timestamp 1644511149
transform 1 0 93748 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1009
timestamp 1644511149
transform 1 0 93932 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1021
timestamp 1644511149
transform 1 0 95036 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1033
timestamp 1644511149
transform 1 0 96140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1045
timestamp 1644511149
transform 1 0 97244 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1057
timestamp 1644511149
transform 1 0 98348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1063
timestamp 1644511149
transform 1 0 98900 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1065
timestamp 1644511149
transform 1 0 99084 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1077
timestamp 1644511149
transform 1 0 100188 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1089
timestamp 1644511149
transform 1 0 101292 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1101
timestamp 1644511149
transform 1 0 102396 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1113
timestamp 1644511149
transform 1 0 103500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1119
timestamp 1644511149
transform 1 0 104052 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1121
timestamp 1644511149
transform 1 0 104236 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1133
timestamp 1644511149
transform 1 0 105340 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1145
timestamp 1644511149
transform 1 0 106444 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1157
timestamp 1644511149
transform 1 0 107548 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1169
timestamp 1644511149
transform 1 0 108652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1175
timestamp 1644511149
transform 1 0 109204 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1177
timestamp 1644511149
transform 1 0 109388 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1189
timestamp 1644511149
transform 1 0 110492 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1201
timestamp 1644511149
transform 1 0 111596 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1213
timestamp 1644511149
transform 1 0 112700 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_1225
timestamp 1644511149
transform 1 0 113804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1231
timestamp 1644511149
transform 1 0 114356 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1233
timestamp 1644511149
transform 1 0 114540 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1245
timestamp 1644511149
transform 1 0 115644 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_1257
timestamp 1644511149
transform 1 0 116748 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_1269
timestamp 1644511149
transform 1 0 117852 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_165
timestamp 1644511149
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1644511149
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_265
timestamp 1644511149
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_289
timestamp 1644511149
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1644511149
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_365
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_377
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_389
timestamp 1644511149
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1644511149
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_501
timestamp 1644511149
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_513
timestamp 1644511149
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1644511149
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_545
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_557
timestamp 1644511149
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_569
timestamp 1644511149
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1644511149
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1644511149
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_601
timestamp 1644511149
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_613
timestamp 1644511149
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_625
timestamp 1644511149
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1644511149
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1644511149
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_645
timestamp 1644511149
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_657
timestamp 1644511149
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_669
timestamp 1644511149
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_681
timestamp 1644511149
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1644511149
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1644511149
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_701
timestamp 1644511149
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_713
timestamp 1644511149
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_725
timestamp 1644511149
transform 1 0 67804 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_737
timestamp 1644511149
transform 1 0 68908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_749
timestamp 1644511149
transform 1 0 70012 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_755
timestamp 1644511149
transform 1 0 70564 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_757
timestamp 1644511149
transform 1 0 70748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_769
timestamp 1644511149
transform 1 0 71852 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_781
timestamp 1644511149
transform 1 0 72956 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_793
timestamp 1644511149
transform 1 0 74060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_805
timestamp 1644511149
transform 1 0 75164 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_811
timestamp 1644511149
transform 1 0 75716 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_813
timestamp 1644511149
transform 1 0 75900 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_825
timestamp 1644511149
transform 1 0 77004 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_837
timestamp 1644511149
transform 1 0 78108 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_849
timestamp 1644511149
transform 1 0 79212 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_861
timestamp 1644511149
transform 1 0 80316 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_867
timestamp 1644511149
transform 1 0 80868 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_869
timestamp 1644511149
transform 1 0 81052 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_881
timestamp 1644511149
transform 1 0 82156 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_893
timestamp 1644511149
transform 1 0 83260 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_905
timestamp 1644511149
transform 1 0 84364 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_917
timestamp 1644511149
transform 1 0 85468 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_923
timestamp 1644511149
transform 1 0 86020 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_925
timestamp 1644511149
transform 1 0 86204 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_937
timestamp 1644511149
transform 1 0 87308 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_949
timestamp 1644511149
transform 1 0 88412 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_961
timestamp 1644511149
transform 1 0 89516 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_973
timestamp 1644511149
transform 1 0 90620 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_979
timestamp 1644511149
transform 1 0 91172 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_981
timestamp 1644511149
transform 1 0 91356 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_993
timestamp 1644511149
transform 1 0 92460 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1005
timestamp 1644511149
transform 1 0 93564 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1017
timestamp 1644511149
transform 1 0 94668 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1029
timestamp 1644511149
transform 1 0 95772 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1035
timestamp 1644511149
transform 1 0 96324 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1037
timestamp 1644511149
transform 1 0 96508 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1049
timestamp 1644511149
transform 1 0 97612 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1061
timestamp 1644511149
transform 1 0 98716 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1073
timestamp 1644511149
transform 1 0 99820 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1085
timestamp 1644511149
transform 1 0 100924 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1091
timestamp 1644511149
transform 1 0 101476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1093
timestamp 1644511149
transform 1 0 101660 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1105
timestamp 1644511149
transform 1 0 102764 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1117
timestamp 1644511149
transform 1 0 103868 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1129
timestamp 1644511149
transform 1 0 104972 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1141
timestamp 1644511149
transform 1 0 106076 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1147
timestamp 1644511149
transform 1 0 106628 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1149
timestamp 1644511149
transform 1 0 106812 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1161
timestamp 1644511149
transform 1 0 107916 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1173
timestamp 1644511149
transform 1 0 109020 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1185
timestamp 1644511149
transform 1 0 110124 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1197
timestamp 1644511149
transform 1 0 111228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1203
timestamp 1644511149
transform 1 0 111780 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1205
timestamp 1644511149
transform 1 0 111964 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1217
timestamp 1644511149
transform 1 0 113068 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1229
timestamp 1644511149
transform 1 0 114172 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_1241
timestamp 1644511149
transform 1 0 115276 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_1253
timestamp 1644511149
transform 1 0 116380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1259
timestamp 1644511149
transform 1 0 116932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_1261
timestamp 1644511149
transform 1 0 117116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_1273
timestamp 1644511149
transform 1 0 118220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_205
timestamp 1644511149
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_261
timestamp 1644511149
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1644511149
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_317
timestamp 1644511149
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_349
timestamp 1644511149
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1644511149
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1644511149
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_517
timestamp 1644511149
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_529
timestamp 1644511149
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_541
timestamp 1644511149
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1644511149
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_585
timestamp 1644511149
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_597
timestamp 1644511149
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1644511149
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1644511149
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_629
timestamp 1644511149
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_641
timestamp 1644511149
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_653
timestamp 1644511149
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1644511149
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1644511149
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_673
timestamp 1644511149
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_685
timestamp 1644511149
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_697
timestamp 1644511149
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_709
timestamp 1644511149
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1644511149
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1644511149
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_729
timestamp 1644511149
transform 1 0 68172 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_741
timestamp 1644511149
transform 1 0 69276 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_753
timestamp 1644511149
transform 1 0 70380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_765
timestamp 1644511149
transform 1 0 71484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_777
timestamp 1644511149
transform 1 0 72588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_783
timestamp 1644511149
transform 1 0 73140 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_785
timestamp 1644511149
transform 1 0 73324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_797
timestamp 1644511149
transform 1 0 74428 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_809
timestamp 1644511149
transform 1 0 75532 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_821
timestamp 1644511149
transform 1 0 76636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_833
timestamp 1644511149
transform 1 0 77740 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_839
timestamp 1644511149
transform 1 0 78292 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_841
timestamp 1644511149
transform 1 0 78476 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_853
timestamp 1644511149
transform 1 0 79580 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_865
timestamp 1644511149
transform 1 0 80684 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_877
timestamp 1644511149
transform 1 0 81788 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_889
timestamp 1644511149
transform 1 0 82892 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_895
timestamp 1644511149
transform 1 0 83444 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_897
timestamp 1644511149
transform 1 0 83628 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_909
timestamp 1644511149
transform 1 0 84732 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_921
timestamp 1644511149
transform 1 0 85836 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_933
timestamp 1644511149
transform 1 0 86940 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_945
timestamp 1644511149
transform 1 0 88044 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_951
timestamp 1644511149
transform 1 0 88596 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_953
timestamp 1644511149
transform 1 0 88780 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_965
timestamp 1644511149
transform 1 0 89884 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_977
timestamp 1644511149
transform 1 0 90988 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_989
timestamp 1644511149
transform 1 0 92092 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1001
timestamp 1644511149
transform 1 0 93196 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1007
timestamp 1644511149
transform 1 0 93748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1009
timestamp 1644511149
transform 1 0 93932 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1021
timestamp 1644511149
transform 1 0 95036 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1033
timestamp 1644511149
transform 1 0 96140 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1045
timestamp 1644511149
transform 1 0 97244 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1057
timestamp 1644511149
transform 1 0 98348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1063
timestamp 1644511149
transform 1 0 98900 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1065
timestamp 1644511149
transform 1 0 99084 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1077
timestamp 1644511149
transform 1 0 100188 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1089
timestamp 1644511149
transform 1 0 101292 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1101
timestamp 1644511149
transform 1 0 102396 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1113
timestamp 1644511149
transform 1 0 103500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1119
timestamp 1644511149
transform 1 0 104052 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1121
timestamp 1644511149
transform 1 0 104236 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1133
timestamp 1644511149
transform 1 0 105340 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1145
timestamp 1644511149
transform 1 0 106444 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1157
timestamp 1644511149
transform 1 0 107548 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1169
timestamp 1644511149
transform 1 0 108652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1175
timestamp 1644511149
transform 1 0 109204 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1177
timestamp 1644511149
transform 1 0 109388 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1189
timestamp 1644511149
transform 1 0 110492 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1201
timestamp 1644511149
transform 1 0 111596 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1213
timestamp 1644511149
transform 1 0 112700 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_1225
timestamp 1644511149
transform 1 0 113804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1231
timestamp 1644511149
transform 1 0 114356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1233
timestamp 1644511149
transform 1 0 114540 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1245
timestamp 1644511149
transform 1 0 115644 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_1257
timestamp 1644511149
transform 1 0 116748 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_1269
timestamp 1644511149
transform 1 0 117852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1644511149
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_289
timestamp 1644511149
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1644511149
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_345
timestamp 1644511149
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1644511149
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_401
timestamp 1644511149
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1644511149
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_513
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1644511149
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_557
timestamp 1644511149
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_569
timestamp 1644511149
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1644511149
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1644511149
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_589
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_601
timestamp 1644511149
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_613
timestamp 1644511149
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_625
timestamp 1644511149
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1644511149
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1644511149
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_645
timestamp 1644511149
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_657
timestamp 1644511149
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_669
timestamp 1644511149
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_681
timestamp 1644511149
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1644511149
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1644511149
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_701
timestamp 1644511149
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_713
timestamp 1644511149
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_725
timestamp 1644511149
transform 1 0 67804 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_737
timestamp 1644511149
transform 1 0 68908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_749
timestamp 1644511149
transform 1 0 70012 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_755
timestamp 1644511149
transform 1 0 70564 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_757
timestamp 1644511149
transform 1 0 70748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_769
timestamp 1644511149
transform 1 0 71852 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_781
timestamp 1644511149
transform 1 0 72956 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_793
timestamp 1644511149
transform 1 0 74060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_805
timestamp 1644511149
transform 1 0 75164 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_811
timestamp 1644511149
transform 1 0 75716 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_813
timestamp 1644511149
transform 1 0 75900 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_825
timestamp 1644511149
transform 1 0 77004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_837
timestamp 1644511149
transform 1 0 78108 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_849
timestamp 1644511149
transform 1 0 79212 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_861
timestamp 1644511149
transform 1 0 80316 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_867
timestamp 1644511149
transform 1 0 80868 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_869
timestamp 1644511149
transform 1 0 81052 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_881
timestamp 1644511149
transform 1 0 82156 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_893
timestamp 1644511149
transform 1 0 83260 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_905
timestamp 1644511149
transform 1 0 84364 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_917
timestamp 1644511149
transform 1 0 85468 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_923
timestamp 1644511149
transform 1 0 86020 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_925
timestamp 1644511149
transform 1 0 86204 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_937
timestamp 1644511149
transform 1 0 87308 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_949
timestamp 1644511149
transform 1 0 88412 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_961
timestamp 1644511149
transform 1 0 89516 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_973
timestamp 1644511149
transform 1 0 90620 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_979
timestamp 1644511149
transform 1 0 91172 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_981
timestamp 1644511149
transform 1 0 91356 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_993
timestamp 1644511149
transform 1 0 92460 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1005
timestamp 1644511149
transform 1 0 93564 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1017
timestamp 1644511149
transform 1 0 94668 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1029
timestamp 1644511149
transform 1 0 95772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1035
timestamp 1644511149
transform 1 0 96324 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1037
timestamp 1644511149
transform 1 0 96508 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1049
timestamp 1644511149
transform 1 0 97612 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1061
timestamp 1644511149
transform 1 0 98716 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1073
timestamp 1644511149
transform 1 0 99820 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1085
timestamp 1644511149
transform 1 0 100924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1091
timestamp 1644511149
transform 1 0 101476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1093
timestamp 1644511149
transform 1 0 101660 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1105
timestamp 1644511149
transform 1 0 102764 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1117
timestamp 1644511149
transform 1 0 103868 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1129
timestamp 1644511149
transform 1 0 104972 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1141
timestamp 1644511149
transform 1 0 106076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1147
timestamp 1644511149
transform 1 0 106628 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1149
timestamp 1644511149
transform 1 0 106812 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1161
timestamp 1644511149
transform 1 0 107916 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1173
timestamp 1644511149
transform 1 0 109020 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1185
timestamp 1644511149
transform 1 0 110124 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1197
timestamp 1644511149
transform 1 0 111228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1203
timestamp 1644511149
transform 1 0 111780 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1205
timestamp 1644511149
transform 1 0 111964 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1217
timestamp 1644511149
transform 1 0 113068 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1229
timestamp 1644511149
transform 1 0 114172 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_1241
timestamp 1644511149
transform 1 0 115276 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_1253
timestamp 1644511149
transform 1 0 116380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_1259
timestamp 1644511149
transform 1 0 116932 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_1261
timestamp 1644511149
transform 1 0 117116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_1273
timestamp 1644511149
transform 1 0 118220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1644511149
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_205
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_237
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1644511149
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1644511149
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_349
timestamp 1644511149
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_361
timestamp 1644511149
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_373
timestamp 1644511149
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1644511149
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1644511149
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_561
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_573
timestamp 1644511149
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_585
timestamp 1644511149
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_597
timestamp 1644511149
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1644511149
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1644511149
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_629
timestamp 1644511149
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_641
timestamp 1644511149
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_653
timestamp 1644511149
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1644511149
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1644511149
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_673
timestamp 1644511149
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_685
timestamp 1644511149
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_697
timestamp 1644511149
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_709
timestamp 1644511149
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1644511149
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1644511149
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_729
timestamp 1644511149
transform 1 0 68172 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_741
timestamp 1644511149
transform 1 0 69276 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_753
timestamp 1644511149
transform 1 0 70380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_765
timestamp 1644511149
transform 1 0 71484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_777
timestamp 1644511149
transform 1 0 72588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_783
timestamp 1644511149
transform 1 0 73140 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_785
timestamp 1644511149
transform 1 0 73324 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_797
timestamp 1644511149
transform 1 0 74428 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_809
timestamp 1644511149
transform 1 0 75532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_821
timestamp 1644511149
transform 1 0 76636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_833
timestamp 1644511149
transform 1 0 77740 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_839
timestamp 1644511149
transform 1 0 78292 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_841
timestamp 1644511149
transform 1 0 78476 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_853
timestamp 1644511149
transform 1 0 79580 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_865
timestamp 1644511149
transform 1 0 80684 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_877
timestamp 1644511149
transform 1 0 81788 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_889
timestamp 1644511149
transform 1 0 82892 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_895
timestamp 1644511149
transform 1 0 83444 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_897
timestamp 1644511149
transform 1 0 83628 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_909
timestamp 1644511149
transform 1 0 84732 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_921
timestamp 1644511149
transform 1 0 85836 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_933
timestamp 1644511149
transform 1 0 86940 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_945
timestamp 1644511149
transform 1 0 88044 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_951
timestamp 1644511149
transform 1 0 88596 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_953
timestamp 1644511149
transform 1 0 88780 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_965
timestamp 1644511149
transform 1 0 89884 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_977
timestamp 1644511149
transform 1 0 90988 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_989
timestamp 1644511149
transform 1 0 92092 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1001
timestamp 1644511149
transform 1 0 93196 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1007
timestamp 1644511149
transform 1 0 93748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1009
timestamp 1644511149
transform 1 0 93932 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1021
timestamp 1644511149
transform 1 0 95036 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1033
timestamp 1644511149
transform 1 0 96140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1045
timestamp 1644511149
transform 1 0 97244 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1057
timestamp 1644511149
transform 1 0 98348 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1063
timestamp 1644511149
transform 1 0 98900 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1065
timestamp 1644511149
transform 1 0 99084 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1077
timestamp 1644511149
transform 1 0 100188 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1089
timestamp 1644511149
transform 1 0 101292 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1101
timestamp 1644511149
transform 1 0 102396 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1113
timestamp 1644511149
transform 1 0 103500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1119
timestamp 1644511149
transform 1 0 104052 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1121
timestamp 1644511149
transform 1 0 104236 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1133
timestamp 1644511149
transform 1 0 105340 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1145
timestamp 1644511149
transform 1 0 106444 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1157
timestamp 1644511149
transform 1 0 107548 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1169
timestamp 1644511149
transform 1 0 108652 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1175
timestamp 1644511149
transform 1 0 109204 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1177
timestamp 1644511149
transform 1 0 109388 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1189
timestamp 1644511149
transform 1 0 110492 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1201
timestamp 1644511149
transform 1 0 111596 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1213
timestamp 1644511149
transform 1 0 112700 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_1225
timestamp 1644511149
transform 1 0 113804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1231
timestamp 1644511149
transform 1 0 114356 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1233
timestamp 1644511149
transform 1 0 114540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1245
timestamp 1644511149
transform 1 0 115644 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_1257
timestamp 1644511149
transform 1 0 116748 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_1273
timestamp 1644511149
transform 1 0 118220 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_153
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_221
timestamp 1644511149
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_233
timestamp 1644511149
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_277
timestamp 1644511149
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_321
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_333
timestamp 1644511149
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_345
timestamp 1644511149
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_401
timestamp 1644511149
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1644511149
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1644511149
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1644511149
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_545
timestamp 1644511149
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_557
timestamp 1644511149
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_569
timestamp 1644511149
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1644511149
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1644511149
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_589
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_625
timestamp 1644511149
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1644511149
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1644511149
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_645
timestamp 1644511149
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_657
timestamp 1644511149
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_669
timestamp 1644511149
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_681
timestamp 1644511149
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1644511149
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1644511149
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_701
timestamp 1644511149
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_713
timestamp 1644511149
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_725
timestamp 1644511149
transform 1 0 67804 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_737
timestamp 1644511149
transform 1 0 68908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_749
timestamp 1644511149
transform 1 0 70012 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_755
timestamp 1644511149
transform 1 0 70564 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_757
timestamp 1644511149
transform 1 0 70748 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_769
timestamp 1644511149
transform 1 0 71852 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_781
timestamp 1644511149
transform 1 0 72956 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_793
timestamp 1644511149
transform 1 0 74060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_805
timestamp 1644511149
transform 1 0 75164 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_811
timestamp 1644511149
transform 1 0 75716 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_813
timestamp 1644511149
transform 1 0 75900 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_825
timestamp 1644511149
transform 1 0 77004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_837
timestamp 1644511149
transform 1 0 78108 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_849
timestamp 1644511149
transform 1 0 79212 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_861
timestamp 1644511149
transform 1 0 80316 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_867
timestamp 1644511149
transform 1 0 80868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_869
timestamp 1644511149
transform 1 0 81052 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_881
timestamp 1644511149
transform 1 0 82156 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_893
timestamp 1644511149
transform 1 0 83260 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_905
timestamp 1644511149
transform 1 0 84364 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_917
timestamp 1644511149
transform 1 0 85468 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_923
timestamp 1644511149
transform 1 0 86020 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_925
timestamp 1644511149
transform 1 0 86204 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_937
timestamp 1644511149
transform 1 0 87308 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_949
timestamp 1644511149
transform 1 0 88412 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_961
timestamp 1644511149
transform 1 0 89516 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_973
timestamp 1644511149
transform 1 0 90620 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_979
timestamp 1644511149
transform 1 0 91172 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_981
timestamp 1644511149
transform 1 0 91356 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_993
timestamp 1644511149
transform 1 0 92460 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1005
timestamp 1644511149
transform 1 0 93564 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1017
timestamp 1644511149
transform 1 0 94668 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1029
timestamp 1644511149
transform 1 0 95772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1035
timestamp 1644511149
transform 1 0 96324 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1037
timestamp 1644511149
transform 1 0 96508 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1049
timestamp 1644511149
transform 1 0 97612 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1061
timestamp 1644511149
transform 1 0 98716 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1073
timestamp 1644511149
transform 1 0 99820 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1085
timestamp 1644511149
transform 1 0 100924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1091
timestamp 1644511149
transform 1 0 101476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1093
timestamp 1644511149
transform 1 0 101660 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1105
timestamp 1644511149
transform 1 0 102764 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1117
timestamp 1644511149
transform 1 0 103868 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1129
timestamp 1644511149
transform 1 0 104972 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1141
timestamp 1644511149
transform 1 0 106076 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1147
timestamp 1644511149
transform 1 0 106628 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1149
timestamp 1644511149
transform 1 0 106812 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1161
timestamp 1644511149
transform 1 0 107916 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1173
timestamp 1644511149
transform 1 0 109020 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1185
timestamp 1644511149
transform 1 0 110124 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1197
timestamp 1644511149
transform 1 0 111228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1203
timestamp 1644511149
transform 1 0 111780 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1205
timestamp 1644511149
transform 1 0 111964 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1217
timestamp 1644511149
transform 1 0 113068 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1229
timestamp 1644511149
transform 1 0 114172 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1241
timestamp 1644511149
transform 1 0 115276 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_1253
timestamp 1644511149
transform 1 0 116380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1259
timestamp 1644511149
transform 1 0 116932 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_1261
timestamp 1644511149
transform 1 0 117116 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_1273
timestamp 1644511149
transform 1 0 118220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1644511149
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1644511149
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_261
timestamp 1644511149
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1644511149
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1644511149
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1644511149
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1644511149
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_361
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_373
timestamp 1644511149
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1644511149
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_517
timestamp 1644511149
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_529
timestamp 1644511149
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_541
timestamp 1644511149
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1644511149
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1644511149
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_585
timestamp 1644511149
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_597
timestamp 1644511149
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1644511149
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1644511149
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_629
timestamp 1644511149
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_641
timestamp 1644511149
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_653
timestamp 1644511149
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1644511149
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1644511149
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_673
timestamp 1644511149
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_685
timestamp 1644511149
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_697
timestamp 1644511149
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_709
timestamp 1644511149
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1644511149
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1644511149
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_729
timestamp 1644511149
transform 1 0 68172 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_741
timestamp 1644511149
transform 1 0 69276 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_753
timestamp 1644511149
transform 1 0 70380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_765
timestamp 1644511149
transform 1 0 71484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_777
timestamp 1644511149
transform 1 0 72588 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_783
timestamp 1644511149
transform 1 0 73140 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_785
timestamp 1644511149
transform 1 0 73324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_797
timestamp 1644511149
transform 1 0 74428 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_809
timestamp 1644511149
transform 1 0 75532 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_821
timestamp 1644511149
transform 1 0 76636 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_833
timestamp 1644511149
transform 1 0 77740 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_839
timestamp 1644511149
transform 1 0 78292 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_841
timestamp 1644511149
transform 1 0 78476 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_853
timestamp 1644511149
transform 1 0 79580 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_865
timestamp 1644511149
transform 1 0 80684 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_877
timestamp 1644511149
transform 1 0 81788 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_889
timestamp 1644511149
transform 1 0 82892 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_895
timestamp 1644511149
transform 1 0 83444 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_897
timestamp 1644511149
transform 1 0 83628 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_909
timestamp 1644511149
transform 1 0 84732 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_921
timestamp 1644511149
transform 1 0 85836 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_933
timestamp 1644511149
transform 1 0 86940 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_945
timestamp 1644511149
transform 1 0 88044 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_951
timestamp 1644511149
transform 1 0 88596 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_953
timestamp 1644511149
transform 1 0 88780 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_965
timestamp 1644511149
transform 1 0 89884 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_977
timestamp 1644511149
transform 1 0 90988 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_989
timestamp 1644511149
transform 1 0 92092 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1001
timestamp 1644511149
transform 1 0 93196 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1007
timestamp 1644511149
transform 1 0 93748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1009
timestamp 1644511149
transform 1 0 93932 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1021
timestamp 1644511149
transform 1 0 95036 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1033
timestamp 1644511149
transform 1 0 96140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1045
timestamp 1644511149
transform 1 0 97244 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1057
timestamp 1644511149
transform 1 0 98348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1063
timestamp 1644511149
transform 1 0 98900 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1065
timestamp 1644511149
transform 1 0 99084 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1077
timestamp 1644511149
transform 1 0 100188 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1089
timestamp 1644511149
transform 1 0 101292 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1101
timestamp 1644511149
transform 1 0 102396 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1113
timestamp 1644511149
transform 1 0 103500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1119
timestamp 1644511149
transform 1 0 104052 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1121
timestamp 1644511149
transform 1 0 104236 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1133
timestamp 1644511149
transform 1 0 105340 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1145
timestamp 1644511149
transform 1 0 106444 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1157
timestamp 1644511149
transform 1 0 107548 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1169
timestamp 1644511149
transform 1 0 108652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1175
timestamp 1644511149
transform 1 0 109204 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1177
timestamp 1644511149
transform 1 0 109388 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1189
timestamp 1644511149
transform 1 0 110492 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1201
timestamp 1644511149
transform 1 0 111596 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1213
timestamp 1644511149
transform 1 0 112700 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_1225
timestamp 1644511149
transform 1 0 113804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1231
timestamp 1644511149
transform 1 0 114356 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1233
timestamp 1644511149
transform 1 0 114540 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1245
timestamp 1644511149
transform 1 0 115644 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_1257
timestamp 1644511149
transform 1 0 116748 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_1273
timestamp 1644511149
transform 1 0 118220 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_165
timestamp 1644511149
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_177
timestamp 1644511149
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_221
timestamp 1644511149
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_233
timestamp 1644511149
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_277
timestamp 1644511149
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1644511149
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1644511149
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_333
timestamp 1644511149
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_345
timestamp 1644511149
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1644511149
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_389
timestamp 1644511149
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_401
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1644511149
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1644511149
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_513
timestamp 1644511149
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1644511149
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1644511149
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_557
timestamp 1644511149
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_569
timestamp 1644511149
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1644511149
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1644511149
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_589
timestamp 1644511149
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_601
timestamp 1644511149
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_625
timestamp 1644511149
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1644511149
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1644511149
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_645
timestamp 1644511149
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_657
timestamp 1644511149
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_669
timestamp 1644511149
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_681
timestamp 1644511149
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1644511149
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1644511149
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_701
timestamp 1644511149
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_713
timestamp 1644511149
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_725
timestamp 1644511149
transform 1 0 67804 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_737
timestamp 1644511149
transform 1 0 68908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_749
timestamp 1644511149
transform 1 0 70012 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_755
timestamp 1644511149
transform 1 0 70564 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_757
timestamp 1644511149
transform 1 0 70748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_769
timestamp 1644511149
transform 1 0 71852 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_781
timestamp 1644511149
transform 1 0 72956 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_793
timestamp 1644511149
transform 1 0 74060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_805
timestamp 1644511149
transform 1 0 75164 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_811
timestamp 1644511149
transform 1 0 75716 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_813
timestamp 1644511149
transform 1 0 75900 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_825
timestamp 1644511149
transform 1 0 77004 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_837
timestamp 1644511149
transform 1 0 78108 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_849
timestamp 1644511149
transform 1 0 79212 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_861
timestamp 1644511149
transform 1 0 80316 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_867
timestamp 1644511149
transform 1 0 80868 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_869
timestamp 1644511149
transform 1 0 81052 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_881
timestamp 1644511149
transform 1 0 82156 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_893
timestamp 1644511149
transform 1 0 83260 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_905
timestamp 1644511149
transform 1 0 84364 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_917
timestamp 1644511149
transform 1 0 85468 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_923
timestamp 1644511149
transform 1 0 86020 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_925
timestamp 1644511149
transform 1 0 86204 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_937
timestamp 1644511149
transform 1 0 87308 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_949
timestamp 1644511149
transform 1 0 88412 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_961
timestamp 1644511149
transform 1 0 89516 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_973
timestamp 1644511149
transform 1 0 90620 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_979
timestamp 1644511149
transform 1 0 91172 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_981
timestamp 1644511149
transform 1 0 91356 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_993
timestamp 1644511149
transform 1 0 92460 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1005
timestamp 1644511149
transform 1 0 93564 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1017
timestamp 1644511149
transform 1 0 94668 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1029
timestamp 1644511149
transform 1 0 95772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1035
timestamp 1644511149
transform 1 0 96324 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1037
timestamp 1644511149
transform 1 0 96508 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1049
timestamp 1644511149
transform 1 0 97612 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1061
timestamp 1644511149
transform 1 0 98716 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1073
timestamp 1644511149
transform 1 0 99820 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1085
timestamp 1644511149
transform 1 0 100924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1091
timestamp 1644511149
transform 1 0 101476 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1093
timestamp 1644511149
transform 1 0 101660 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1105
timestamp 1644511149
transform 1 0 102764 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1117
timestamp 1644511149
transform 1 0 103868 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1129
timestamp 1644511149
transform 1 0 104972 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1141
timestamp 1644511149
transform 1 0 106076 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1147
timestamp 1644511149
transform 1 0 106628 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1149
timestamp 1644511149
transform 1 0 106812 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1161
timestamp 1644511149
transform 1 0 107916 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1173
timestamp 1644511149
transform 1 0 109020 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1185
timestamp 1644511149
transform 1 0 110124 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1197
timestamp 1644511149
transform 1 0 111228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1203
timestamp 1644511149
transform 1 0 111780 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1205
timestamp 1644511149
transform 1 0 111964 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1217
timestamp 1644511149
transform 1 0 113068 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1229
timestamp 1644511149
transform 1 0 114172 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1241
timestamp 1644511149
transform 1 0 115276 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_1253
timestamp 1644511149
transform 1 0 116380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_1259
timestamp 1644511149
transform 1 0 116932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_1261
timestamp 1644511149
transform 1 0 117116 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_1273
timestamp 1644511149
transform 1 0 118220 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1644511149
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_205
timestamp 1644511149
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_237
timestamp 1644511149
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_261
timestamp 1644511149
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_305
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_317
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1644511149
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_361
timestamp 1644511149
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_373
timestamp 1644511149
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1644511149
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_517
timestamp 1644511149
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_529
timestamp 1644511149
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_541
timestamp 1644511149
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1644511149
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_561
timestamp 1644511149
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_573
timestamp 1644511149
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_585
timestamp 1644511149
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_597
timestamp 1644511149
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1644511149
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1644511149
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_629
timestamp 1644511149
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_641
timestamp 1644511149
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_653
timestamp 1644511149
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1644511149
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1644511149
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_673
timestamp 1644511149
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_685
timestamp 1644511149
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_697
timestamp 1644511149
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_709
timestamp 1644511149
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 1644511149
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 1644511149
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_729
timestamp 1644511149
transform 1 0 68172 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_741
timestamp 1644511149
transform 1 0 69276 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_753
timestamp 1644511149
transform 1 0 70380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_765
timestamp 1644511149
transform 1 0 71484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_777
timestamp 1644511149
transform 1 0 72588 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_783
timestamp 1644511149
transform 1 0 73140 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_785
timestamp 1644511149
transform 1 0 73324 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_797
timestamp 1644511149
transform 1 0 74428 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_809
timestamp 1644511149
transform 1 0 75532 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_821
timestamp 1644511149
transform 1 0 76636 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_833
timestamp 1644511149
transform 1 0 77740 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_839
timestamp 1644511149
transform 1 0 78292 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_841
timestamp 1644511149
transform 1 0 78476 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_853
timestamp 1644511149
transform 1 0 79580 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_865
timestamp 1644511149
transform 1 0 80684 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_877
timestamp 1644511149
transform 1 0 81788 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_889
timestamp 1644511149
transform 1 0 82892 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_895
timestamp 1644511149
transform 1 0 83444 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_897
timestamp 1644511149
transform 1 0 83628 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_909
timestamp 1644511149
transform 1 0 84732 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_921
timestamp 1644511149
transform 1 0 85836 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_933
timestamp 1644511149
transform 1 0 86940 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_945
timestamp 1644511149
transform 1 0 88044 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_951
timestamp 1644511149
transform 1 0 88596 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_953
timestamp 1644511149
transform 1 0 88780 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_965
timestamp 1644511149
transform 1 0 89884 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_977
timestamp 1644511149
transform 1 0 90988 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_989
timestamp 1644511149
transform 1 0 92092 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1001
timestamp 1644511149
transform 1 0 93196 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1007
timestamp 1644511149
transform 1 0 93748 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1009
timestamp 1644511149
transform 1 0 93932 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1021
timestamp 1644511149
transform 1 0 95036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1033
timestamp 1644511149
transform 1 0 96140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1045
timestamp 1644511149
transform 1 0 97244 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1057
timestamp 1644511149
transform 1 0 98348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1063
timestamp 1644511149
transform 1 0 98900 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1065
timestamp 1644511149
transform 1 0 99084 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1077
timestamp 1644511149
transform 1 0 100188 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1089
timestamp 1644511149
transform 1 0 101292 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1101
timestamp 1644511149
transform 1 0 102396 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1113
timestamp 1644511149
transform 1 0 103500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1119
timestamp 1644511149
transform 1 0 104052 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1121
timestamp 1644511149
transform 1 0 104236 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1133
timestamp 1644511149
transform 1 0 105340 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1145
timestamp 1644511149
transform 1 0 106444 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1157
timestamp 1644511149
transform 1 0 107548 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1169
timestamp 1644511149
transform 1 0 108652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1175
timestamp 1644511149
transform 1 0 109204 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1177
timestamp 1644511149
transform 1 0 109388 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1189
timestamp 1644511149
transform 1 0 110492 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1201
timestamp 1644511149
transform 1 0 111596 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1213
timestamp 1644511149
transform 1 0 112700 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_1225
timestamp 1644511149
transform 1 0 113804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1231
timestamp 1644511149
transform 1 0 114356 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1233
timestamp 1644511149
transform 1 0 114540 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1245
timestamp 1644511149
transform 1 0 115644 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_1257
timestamp 1644511149
transform 1 0 116748 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_1273
timestamp 1644511149
transform 1 0 118220 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1644511149
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_333
timestamp 1644511149
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_345
timestamp 1644511149
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1644511149
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_377
timestamp 1644511149
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_389
timestamp 1644511149
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1644511149
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_501
timestamp 1644511149
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_513
timestamp 1644511149
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1644511149
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_625
timestamp 1644511149
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1644511149
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1644511149
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_645
timestamp 1644511149
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_657
timestamp 1644511149
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_669
timestamp 1644511149
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_681
timestamp 1644511149
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1644511149
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1644511149
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_701
timestamp 1644511149
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_713
timestamp 1644511149
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_725
timestamp 1644511149
transform 1 0 67804 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_737
timestamp 1644511149
transform 1 0 68908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_749
timestamp 1644511149
transform 1 0 70012 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_755
timestamp 1644511149
transform 1 0 70564 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_757
timestamp 1644511149
transform 1 0 70748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_769
timestamp 1644511149
transform 1 0 71852 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_781
timestamp 1644511149
transform 1 0 72956 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_793
timestamp 1644511149
transform 1 0 74060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_805
timestamp 1644511149
transform 1 0 75164 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_811
timestamp 1644511149
transform 1 0 75716 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_813
timestamp 1644511149
transform 1 0 75900 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_825
timestamp 1644511149
transform 1 0 77004 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_837
timestamp 1644511149
transform 1 0 78108 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_849
timestamp 1644511149
transform 1 0 79212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_861
timestamp 1644511149
transform 1 0 80316 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_867
timestamp 1644511149
transform 1 0 80868 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_869
timestamp 1644511149
transform 1 0 81052 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_881
timestamp 1644511149
transform 1 0 82156 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_893
timestamp 1644511149
transform 1 0 83260 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_905
timestamp 1644511149
transform 1 0 84364 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_917
timestamp 1644511149
transform 1 0 85468 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_923
timestamp 1644511149
transform 1 0 86020 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_925
timestamp 1644511149
transform 1 0 86204 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_937
timestamp 1644511149
transform 1 0 87308 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_949
timestamp 1644511149
transform 1 0 88412 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_961
timestamp 1644511149
transform 1 0 89516 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_973
timestamp 1644511149
transform 1 0 90620 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_979
timestamp 1644511149
transform 1 0 91172 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_981
timestamp 1644511149
transform 1 0 91356 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_993
timestamp 1644511149
transform 1 0 92460 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1005
timestamp 1644511149
transform 1 0 93564 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1017
timestamp 1644511149
transform 1 0 94668 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1029
timestamp 1644511149
transform 1 0 95772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1035
timestamp 1644511149
transform 1 0 96324 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1037
timestamp 1644511149
transform 1 0 96508 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1049
timestamp 1644511149
transform 1 0 97612 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1061
timestamp 1644511149
transform 1 0 98716 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1073
timestamp 1644511149
transform 1 0 99820 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1085
timestamp 1644511149
transform 1 0 100924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1091
timestamp 1644511149
transform 1 0 101476 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1093
timestamp 1644511149
transform 1 0 101660 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1105
timestamp 1644511149
transform 1 0 102764 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1117
timestamp 1644511149
transform 1 0 103868 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1129
timestamp 1644511149
transform 1 0 104972 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1141
timestamp 1644511149
transform 1 0 106076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1147
timestamp 1644511149
transform 1 0 106628 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1149
timestamp 1644511149
transform 1 0 106812 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1161
timestamp 1644511149
transform 1 0 107916 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1173
timestamp 1644511149
transform 1 0 109020 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1185
timestamp 1644511149
transform 1 0 110124 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1197
timestamp 1644511149
transform 1 0 111228 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1203
timestamp 1644511149
transform 1 0 111780 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1205
timestamp 1644511149
transform 1 0 111964 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1217
timestamp 1644511149
transform 1 0 113068 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1229
timestamp 1644511149
transform 1 0 114172 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1241
timestamp 1644511149
transform 1 0 115276 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_1253
timestamp 1644511149
transform 1 0 116380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1259
timestamp 1644511149
transform 1 0 116932 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_1261
timestamp 1644511149
transform 1 0 117116 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_1273
timestamp 1644511149
transform 1 0 118220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1644511149
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1644511149
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_517
timestamp 1644511149
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_529
timestamp 1644511149
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_541
timestamp 1644511149
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1644511149
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1644511149
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_561
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_573
timestamp 1644511149
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_585
timestamp 1644511149
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_597
timestamp 1644511149
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1644511149
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1644511149
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_617
timestamp 1644511149
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_629
timestamp 1644511149
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_641
timestamp 1644511149
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_653
timestamp 1644511149
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1644511149
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1644511149
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_673
timestamp 1644511149
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_685
timestamp 1644511149
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_697
timestamp 1644511149
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_709
timestamp 1644511149
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1644511149
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1644511149
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_729
timestamp 1644511149
transform 1 0 68172 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_741
timestamp 1644511149
transform 1 0 69276 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_753
timestamp 1644511149
transform 1 0 70380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_765
timestamp 1644511149
transform 1 0 71484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_777
timestamp 1644511149
transform 1 0 72588 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_783
timestamp 1644511149
transform 1 0 73140 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_785
timestamp 1644511149
transform 1 0 73324 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_797
timestamp 1644511149
transform 1 0 74428 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_809
timestamp 1644511149
transform 1 0 75532 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_821
timestamp 1644511149
transform 1 0 76636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_833
timestamp 1644511149
transform 1 0 77740 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_839
timestamp 1644511149
transform 1 0 78292 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_841
timestamp 1644511149
transform 1 0 78476 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_853
timestamp 1644511149
transform 1 0 79580 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_865
timestamp 1644511149
transform 1 0 80684 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_877
timestamp 1644511149
transform 1 0 81788 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_889
timestamp 1644511149
transform 1 0 82892 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_895
timestamp 1644511149
transform 1 0 83444 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_897
timestamp 1644511149
transform 1 0 83628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_909
timestamp 1644511149
transform 1 0 84732 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_921
timestamp 1644511149
transform 1 0 85836 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_933
timestamp 1644511149
transform 1 0 86940 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_945
timestamp 1644511149
transform 1 0 88044 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_951
timestamp 1644511149
transform 1 0 88596 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_953
timestamp 1644511149
transform 1 0 88780 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_965
timestamp 1644511149
transform 1 0 89884 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_977
timestamp 1644511149
transform 1 0 90988 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_989
timestamp 1644511149
transform 1 0 92092 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1001
timestamp 1644511149
transform 1 0 93196 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1007
timestamp 1644511149
transform 1 0 93748 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1009
timestamp 1644511149
transform 1 0 93932 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1021
timestamp 1644511149
transform 1 0 95036 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1033
timestamp 1644511149
transform 1 0 96140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1045
timestamp 1644511149
transform 1 0 97244 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1057
timestamp 1644511149
transform 1 0 98348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1063
timestamp 1644511149
transform 1 0 98900 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1065
timestamp 1644511149
transform 1 0 99084 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1077
timestamp 1644511149
transform 1 0 100188 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1089
timestamp 1644511149
transform 1 0 101292 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1101
timestamp 1644511149
transform 1 0 102396 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1113
timestamp 1644511149
transform 1 0 103500 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1119
timestamp 1644511149
transform 1 0 104052 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1121
timestamp 1644511149
transform 1 0 104236 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1133
timestamp 1644511149
transform 1 0 105340 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1145
timestamp 1644511149
transform 1 0 106444 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1157
timestamp 1644511149
transform 1 0 107548 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1169
timestamp 1644511149
transform 1 0 108652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1175
timestamp 1644511149
transform 1 0 109204 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1177
timestamp 1644511149
transform 1 0 109388 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1189
timestamp 1644511149
transform 1 0 110492 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1201
timestamp 1644511149
transform 1 0 111596 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1213
timestamp 1644511149
transform 1 0 112700 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_1225
timestamp 1644511149
transform 1 0 113804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1231
timestamp 1644511149
transform 1 0 114356 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1233
timestamp 1644511149
transform 1 0 114540 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1245
timestamp 1644511149
transform 1 0 115644 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_1257
timestamp 1644511149
transform 1 0 116748 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_1273
timestamp 1644511149
transform 1 0 118220 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_265
timestamp 1644511149
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1644511149
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_333
timestamp 1644511149
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_345
timestamp 1644511149
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1644511149
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1644511149
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_501
timestamp 1644511149
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_513
timestamp 1644511149
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1644511149
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1644511149
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_545
timestamp 1644511149
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_557
timestamp 1644511149
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_569
timestamp 1644511149
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1644511149
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1644511149
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_625
timestamp 1644511149
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1644511149
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1644511149
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_645
timestamp 1644511149
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_657
timestamp 1644511149
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_669
timestamp 1644511149
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_681
timestamp 1644511149
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1644511149
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1644511149
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_701
timestamp 1644511149
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_713
timestamp 1644511149
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_725
timestamp 1644511149
transform 1 0 67804 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_737
timestamp 1644511149
transform 1 0 68908 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_749
timestamp 1644511149
transform 1 0 70012 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_755
timestamp 1644511149
transform 1 0 70564 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_757
timestamp 1644511149
transform 1 0 70748 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_769
timestamp 1644511149
transform 1 0 71852 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_781
timestamp 1644511149
transform 1 0 72956 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_793
timestamp 1644511149
transform 1 0 74060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_805
timestamp 1644511149
transform 1 0 75164 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_811
timestamp 1644511149
transform 1 0 75716 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_813
timestamp 1644511149
transform 1 0 75900 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_825
timestamp 1644511149
transform 1 0 77004 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_837
timestamp 1644511149
transform 1 0 78108 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_849
timestamp 1644511149
transform 1 0 79212 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_861
timestamp 1644511149
transform 1 0 80316 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_867
timestamp 1644511149
transform 1 0 80868 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_869
timestamp 1644511149
transform 1 0 81052 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_881
timestamp 1644511149
transform 1 0 82156 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_893
timestamp 1644511149
transform 1 0 83260 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_905
timestamp 1644511149
transform 1 0 84364 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_917
timestamp 1644511149
transform 1 0 85468 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_923
timestamp 1644511149
transform 1 0 86020 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_925
timestamp 1644511149
transform 1 0 86204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_937
timestamp 1644511149
transform 1 0 87308 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_949
timestamp 1644511149
transform 1 0 88412 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_961
timestamp 1644511149
transform 1 0 89516 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_973
timestamp 1644511149
transform 1 0 90620 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_979
timestamp 1644511149
transform 1 0 91172 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_981
timestamp 1644511149
transform 1 0 91356 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_993
timestamp 1644511149
transform 1 0 92460 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1005
timestamp 1644511149
transform 1 0 93564 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1017
timestamp 1644511149
transform 1 0 94668 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1029
timestamp 1644511149
transform 1 0 95772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1035
timestamp 1644511149
transform 1 0 96324 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1037
timestamp 1644511149
transform 1 0 96508 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1049
timestamp 1644511149
transform 1 0 97612 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1061
timestamp 1644511149
transform 1 0 98716 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1073
timestamp 1644511149
transform 1 0 99820 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1085
timestamp 1644511149
transform 1 0 100924 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1091
timestamp 1644511149
transform 1 0 101476 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1093
timestamp 1644511149
transform 1 0 101660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1105
timestamp 1644511149
transform 1 0 102764 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1117
timestamp 1644511149
transform 1 0 103868 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1129
timestamp 1644511149
transform 1 0 104972 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1141
timestamp 1644511149
transform 1 0 106076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1147
timestamp 1644511149
transform 1 0 106628 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1149
timestamp 1644511149
transform 1 0 106812 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1161
timestamp 1644511149
transform 1 0 107916 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1173
timestamp 1644511149
transform 1 0 109020 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1185
timestamp 1644511149
transform 1 0 110124 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1197
timestamp 1644511149
transform 1 0 111228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1203
timestamp 1644511149
transform 1 0 111780 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1205
timestamp 1644511149
transform 1 0 111964 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1217
timestamp 1644511149
transform 1 0 113068 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1229
timestamp 1644511149
transform 1 0 114172 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_1241
timestamp 1644511149
transform 1 0 115276 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_1253
timestamp 1644511149
transform 1 0 116380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1259
timestamp 1644511149
transform 1 0 116932 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_1261
timestamp 1644511149
transform 1 0 117116 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_1273
timestamp 1644511149
transform 1 0 118220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1644511149
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_305
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_317
timestamp 1644511149
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1644511149
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1644511149
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_361
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1644511149
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1644511149
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1644511149
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_517
timestamp 1644511149
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_529
timestamp 1644511149
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_541
timestamp 1644511149
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1644511149
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_561
timestamp 1644511149
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_573
timestamp 1644511149
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_585
timestamp 1644511149
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_597
timestamp 1644511149
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1644511149
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1644511149
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_629
timestamp 1644511149
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_641
timestamp 1644511149
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_653
timestamp 1644511149
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1644511149
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1644511149
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_673
timestamp 1644511149
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_685
timestamp 1644511149
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_697
timestamp 1644511149
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_709
timestamp 1644511149
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1644511149
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1644511149
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_729
timestamp 1644511149
transform 1 0 68172 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_741
timestamp 1644511149
transform 1 0 69276 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_753
timestamp 1644511149
transform 1 0 70380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_765
timestamp 1644511149
transform 1 0 71484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_777
timestamp 1644511149
transform 1 0 72588 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_783
timestamp 1644511149
transform 1 0 73140 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_785
timestamp 1644511149
transform 1 0 73324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_797
timestamp 1644511149
transform 1 0 74428 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_809
timestamp 1644511149
transform 1 0 75532 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_821
timestamp 1644511149
transform 1 0 76636 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_833
timestamp 1644511149
transform 1 0 77740 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_839
timestamp 1644511149
transform 1 0 78292 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_841
timestamp 1644511149
transform 1 0 78476 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_853
timestamp 1644511149
transform 1 0 79580 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_865
timestamp 1644511149
transform 1 0 80684 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_877
timestamp 1644511149
transform 1 0 81788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_889
timestamp 1644511149
transform 1 0 82892 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_895
timestamp 1644511149
transform 1 0 83444 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_897
timestamp 1644511149
transform 1 0 83628 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_909
timestamp 1644511149
transform 1 0 84732 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_921
timestamp 1644511149
transform 1 0 85836 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_933
timestamp 1644511149
transform 1 0 86940 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_945
timestamp 1644511149
transform 1 0 88044 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_951
timestamp 1644511149
transform 1 0 88596 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_953
timestamp 1644511149
transform 1 0 88780 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_965
timestamp 1644511149
transform 1 0 89884 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_977
timestamp 1644511149
transform 1 0 90988 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_989
timestamp 1644511149
transform 1 0 92092 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1001
timestamp 1644511149
transform 1 0 93196 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1007
timestamp 1644511149
transform 1 0 93748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1009
timestamp 1644511149
transform 1 0 93932 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1021
timestamp 1644511149
transform 1 0 95036 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1033
timestamp 1644511149
transform 1 0 96140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1045
timestamp 1644511149
transform 1 0 97244 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1057
timestamp 1644511149
transform 1 0 98348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1063
timestamp 1644511149
transform 1 0 98900 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1065
timestamp 1644511149
transform 1 0 99084 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1077
timestamp 1644511149
transform 1 0 100188 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1089
timestamp 1644511149
transform 1 0 101292 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1101
timestamp 1644511149
transform 1 0 102396 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1113
timestamp 1644511149
transform 1 0 103500 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1119
timestamp 1644511149
transform 1 0 104052 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1121
timestamp 1644511149
transform 1 0 104236 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1133
timestamp 1644511149
transform 1 0 105340 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1145
timestamp 1644511149
transform 1 0 106444 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1157
timestamp 1644511149
transform 1 0 107548 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1169
timestamp 1644511149
transform 1 0 108652 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1175
timestamp 1644511149
transform 1 0 109204 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1177
timestamp 1644511149
transform 1 0 109388 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1189
timestamp 1644511149
transform 1 0 110492 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1201
timestamp 1644511149
transform 1 0 111596 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1213
timestamp 1644511149
transform 1 0 112700 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_1225
timestamp 1644511149
transform 1 0 113804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1231
timestamp 1644511149
transform 1 0 114356 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1233
timestamp 1644511149
transform 1 0 114540 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1245
timestamp 1644511149
transform 1 0 115644 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1257
timestamp 1644511149
transform 1 0 116748 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1269
timestamp 1644511149
transform 1 0 117852 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_221
timestamp 1644511149
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_233
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_265
timestamp 1644511149
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_289
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_513
timestamp 1644511149
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_533
timestamp 1644511149
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_545
timestamp 1644511149
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_557
timestamp 1644511149
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_569
timestamp 1644511149
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1644511149
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_625
timestamp 1644511149
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1644511149
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1644511149
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_645
timestamp 1644511149
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_657
timestamp 1644511149
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_669
timestamp 1644511149
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_681
timestamp 1644511149
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1644511149
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1644511149
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_701
timestamp 1644511149
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_713
timestamp 1644511149
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_725
timestamp 1644511149
transform 1 0 67804 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_737
timestamp 1644511149
transform 1 0 68908 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_749
timestamp 1644511149
transform 1 0 70012 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_755
timestamp 1644511149
transform 1 0 70564 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_757
timestamp 1644511149
transform 1 0 70748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_769
timestamp 1644511149
transform 1 0 71852 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_781
timestamp 1644511149
transform 1 0 72956 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_793
timestamp 1644511149
transform 1 0 74060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_805
timestamp 1644511149
transform 1 0 75164 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_811
timestamp 1644511149
transform 1 0 75716 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_813
timestamp 1644511149
transform 1 0 75900 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_825
timestamp 1644511149
transform 1 0 77004 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_837
timestamp 1644511149
transform 1 0 78108 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_849
timestamp 1644511149
transform 1 0 79212 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_861
timestamp 1644511149
transform 1 0 80316 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_867
timestamp 1644511149
transform 1 0 80868 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_869
timestamp 1644511149
transform 1 0 81052 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_881
timestamp 1644511149
transform 1 0 82156 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_893
timestamp 1644511149
transform 1 0 83260 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_905
timestamp 1644511149
transform 1 0 84364 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_917
timestamp 1644511149
transform 1 0 85468 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_923
timestamp 1644511149
transform 1 0 86020 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_925
timestamp 1644511149
transform 1 0 86204 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_937
timestamp 1644511149
transform 1 0 87308 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_949
timestamp 1644511149
transform 1 0 88412 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_961
timestamp 1644511149
transform 1 0 89516 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_973
timestamp 1644511149
transform 1 0 90620 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_979
timestamp 1644511149
transform 1 0 91172 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_981
timestamp 1644511149
transform 1 0 91356 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_993
timestamp 1644511149
transform 1 0 92460 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1005
timestamp 1644511149
transform 1 0 93564 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1017
timestamp 1644511149
transform 1 0 94668 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1029
timestamp 1644511149
transform 1 0 95772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1035
timestamp 1644511149
transform 1 0 96324 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1037
timestamp 1644511149
transform 1 0 96508 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1049
timestamp 1644511149
transform 1 0 97612 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1061
timestamp 1644511149
transform 1 0 98716 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1073
timestamp 1644511149
transform 1 0 99820 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1085
timestamp 1644511149
transform 1 0 100924 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1091
timestamp 1644511149
transform 1 0 101476 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1093
timestamp 1644511149
transform 1 0 101660 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1105
timestamp 1644511149
transform 1 0 102764 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1117
timestamp 1644511149
transform 1 0 103868 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1129
timestamp 1644511149
transform 1 0 104972 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1141
timestamp 1644511149
transform 1 0 106076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1147
timestamp 1644511149
transform 1 0 106628 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1149
timestamp 1644511149
transform 1 0 106812 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1161
timestamp 1644511149
transform 1 0 107916 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1173
timestamp 1644511149
transform 1 0 109020 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1185
timestamp 1644511149
transform 1 0 110124 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1197
timestamp 1644511149
transform 1 0 111228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1203
timestamp 1644511149
transform 1 0 111780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1205
timestamp 1644511149
transform 1 0 111964 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1217
timestamp 1644511149
transform 1 0 113068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1229
timestamp 1644511149
transform 1 0 114172 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1241
timestamp 1644511149
transform 1 0 115276 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_1253
timestamp 1644511149
transform 1 0 116380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1259
timestamp 1644511149
transform 1 0 116932 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_1261
timestamp 1644511149
transform 1 0 117116 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1273
timestamp 1644511149
transform 1 0 118220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1644511149
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_305
timestamp 1644511149
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_529
timestamp 1644511149
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_541
timestamp 1644511149
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1644511149
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1644511149
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_629
timestamp 1644511149
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_641
timestamp 1644511149
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_653
timestamp 1644511149
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1644511149
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1644511149
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_673
timestamp 1644511149
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_685
timestamp 1644511149
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_697
timestamp 1644511149
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_709
timestamp 1644511149
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1644511149
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1644511149
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_729
timestamp 1644511149
transform 1 0 68172 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_741
timestamp 1644511149
transform 1 0 69276 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_753
timestamp 1644511149
transform 1 0 70380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_765
timestamp 1644511149
transform 1 0 71484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_777
timestamp 1644511149
transform 1 0 72588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_783
timestamp 1644511149
transform 1 0 73140 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_785
timestamp 1644511149
transform 1 0 73324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_797
timestamp 1644511149
transform 1 0 74428 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_809
timestamp 1644511149
transform 1 0 75532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_821
timestamp 1644511149
transform 1 0 76636 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_833
timestamp 1644511149
transform 1 0 77740 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_839
timestamp 1644511149
transform 1 0 78292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_841
timestamp 1644511149
transform 1 0 78476 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_853
timestamp 1644511149
transform 1 0 79580 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_865
timestamp 1644511149
transform 1 0 80684 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_877
timestamp 1644511149
transform 1 0 81788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_889
timestamp 1644511149
transform 1 0 82892 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_895
timestamp 1644511149
transform 1 0 83444 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_897
timestamp 1644511149
transform 1 0 83628 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_909
timestamp 1644511149
transform 1 0 84732 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_921
timestamp 1644511149
transform 1 0 85836 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_933
timestamp 1644511149
transform 1 0 86940 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_945
timestamp 1644511149
transform 1 0 88044 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_951
timestamp 1644511149
transform 1 0 88596 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_953
timestamp 1644511149
transform 1 0 88780 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_965
timestamp 1644511149
transform 1 0 89884 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_977
timestamp 1644511149
transform 1 0 90988 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_989
timestamp 1644511149
transform 1 0 92092 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1001
timestamp 1644511149
transform 1 0 93196 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1007
timestamp 1644511149
transform 1 0 93748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1009
timestamp 1644511149
transform 1 0 93932 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1021
timestamp 1644511149
transform 1 0 95036 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1033
timestamp 1644511149
transform 1 0 96140 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1045
timestamp 1644511149
transform 1 0 97244 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1057
timestamp 1644511149
transform 1 0 98348 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1063
timestamp 1644511149
transform 1 0 98900 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1065
timestamp 1644511149
transform 1 0 99084 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1077
timestamp 1644511149
transform 1 0 100188 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1089
timestamp 1644511149
transform 1 0 101292 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1101
timestamp 1644511149
transform 1 0 102396 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1113
timestamp 1644511149
transform 1 0 103500 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1119
timestamp 1644511149
transform 1 0 104052 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1121
timestamp 1644511149
transform 1 0 104236 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1133
timestamp 1644511149
transform 1 0 105340 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1145
timestamp 1644511149
transform 1 0 106444 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1157
timestamp 1644511149
transform 1 0 107548 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1169
timestamp 1644511149
transform 1 0 108652 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1175
timestamp 1644511149
transform 1 0 109204 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1177
timestamp 1644511149
transform 1 0 109388 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1189
timestamp 1644511149
transform 1 0 110492 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1201
timestamp 1644511149
transform 1 0 111596 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1213
timestamp 1644511149
transform 1 0 112700 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_1225
timestamp 1644511149
transform 1 0 113804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1231
timestamp 1644511149
transform 1 0 114356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1233
timestamp 1644511149
transform 1 0 114540 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1245
timestamp 1644511149
transform 1 0 115644 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1257
timestamp 1644511149
transform 1 0 116748 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1269
timestamp 1644511149
transform 1 0 117852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_289
timestamp 1644511149
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1644511149
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1644511149
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_513
timestamp 1644511149
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1644511149
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_625
timestamp 1644511149
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1644511149
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1644511149
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_645
timestamp 1644511149
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_657
timestamp 1644511149
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_669
timestamp 1644511149
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_681
timestamp 1644511149
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1644511149
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1644511149
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_701
timestamp 1644511149
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_713
timestamp 1644511149
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_725
timestamp 1644511149
transform 1 0 67804 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_737
timestamp 1644511149
transform 1 0 68908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_749
timestamp 1644511149
transform 1 0 70012 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_755
timestamp 1644511149
transform 1 0 70564 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_757
timestamp 1644511149
transform 1 0 70748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_769
timestamp 1644511149
transform 1 0 71852 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_781
timestamp 1644511149
transform 1 0 72956 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_793
timestamp 1644511149
transform 1 0 74060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_805
timestamp 1644511149
transform 1 0 75164 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_811
timestamp 1644511149
transform 1 0 75716 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_813
timestamp 1644511149
transform 1 0 75900 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_825
timestamp 1644511149
transform 1 0 77004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_837
timestamp 1644511149
transform 1 0 78108 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_849
timestamp 1644511149
transform 1 0 79212 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_861
timestamp 1644511149
transform 1 0 80316 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_867
timestamp 1644511149
transform 1 0 80868 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_869
timestamp 1644511149
transform 1 0 81052 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_881
timestamp 1644511149
transform 1 0 82156 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_893
timestamp 1644511149
transform 1 0 83260 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_905
timestamp 1644511149
transform 1 0 84364 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_917
timestamp 1644511149
transform 1 0 85468 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_923
timestamp 1644511149
transform 1 0 86020 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_925
timestamp 1644511149
transform 1 0 86204 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_937
timestamp 1644511149
transform 1 0 87308 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_949
timestamp 1644511149
transform 1 0 88412 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_961
timestamp 1644511149
transform 1 0 89516 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_973
timestamp 1644511149
transform 1 0 90620 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_979
timestamp 1644511149
transform 1 0 91172 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_981
timestamp 1644511149
transform 1 0 91356 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_993
timestamp 1644511149
transform 1 0 92460 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1005
timestamp 1644511149
transform 1 0 93564 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1017
timestamp 1644511149
transform 1 0 94668 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1029
timestamp 1644511149
transform 1 0 95772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1035
timestamp 1644511149
transform 1 0 96324 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1037
timestamp 1644511149
transform 1 0 96508 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1049
timestamp 1644511149
transform 1 0 97612 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1061
timestamp 1644511149
transform 1 0 98716 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1073
timestamp 1644511149
transform 1 0 99820 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1085
timestamp 1644511149
transform 1 0 100924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1091
timestamp 1644511149
transform 1 0 101476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1093
timestamp 1644511149
transform 1 0 101660 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1105
timestamp 1644511149
transform 1 0 102764 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1117
timestamp 1644511149
transform 1 0 103868 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1129
timestamp 1644511149
transform 1 0 104972 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1141
timestamp 1644511149
transform 1 0 106076 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1147
timestamp 1644511149
transform 1 0 106628 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1149
timestamp 1644511149
transform 1 0 106812 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1161
timestamp 1644511149
transform 1 0 107916 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1173
timestamp 1644511149
transform 1 0 109020 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1185
timestamp 1644511149
transform 1 0 110124 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1197
timestamp 1644511149
transform 1 0 111228 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1203
timestamp 1644511149
transform 1 0 111780 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1205
timestamp 1644511149
transform 1 0 111964 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1217
timestamp 1644511149
transform 1 0 113068 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1229
timestamp 1644511149
transform 1 0 114172 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1241
timestamp 1644511149
transform 1 0 115276 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1253
timestamp 1644511149
transform 1 0 116380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1259
timestamp 1644511149
transform 1 0 116932 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1261
timestamp 1644511149
transform 1 0 117116 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_1273
timestamp 1644511149
transform 1 0 118220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_261
timestamp 1644511149
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1644511149
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1644511149
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_317
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1644511149
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_505
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_517
timestamp 1644511149
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_529
timestamp 1644511149
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_541
timestamp 1644511149
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1644511149
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1644511149
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1644511149
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1644511149
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_617
timestamp 1644511149
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_629
timestamp 1644511149
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_641
timestamp 1644511149
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_653
timestamp 1644511149
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1644511149
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1644511149
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_673
timestamp 1644511149
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_685
timestamp 1644511149
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_697
timestamp 1644511149
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_709
timestamp 1644511149
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1644511149
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1644511149
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_729
timestamp 1644511149
transform 1 0 68172 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_741
timestamp 1644511149
transform 1 0 69276 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_753
timestamp 1644511149
transform 1 0 70380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_765
timestamp 1644511149
transform 1 0 71484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_777
timestamp 1644511149
transform 1 0 72588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_783
timestamp 1644511149
transform 1 0 73140 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_785
timestamp 1644511149
transform 1 0 73324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_797
timestamp 1644511149
transform 1 0 74428 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_809
timestamp 1644511149
transform 1 0 75532 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_821
timestamp 1644511149
transform 1 0 76636 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_833
timestamp 1644511149
transform 1 0 77740 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_839
timestamp 1644511149
transform 1 0 78292 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_841
timestamp 1644511149
transform 1 0 78476 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_853
timestamp 1644511149
transform 1 0 79580 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_865
timestamp 1644511149
transform 1 0 80684 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_877
timestamp 1644511149
transform 1 0 81788 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_889
timestamp 1644511149
transform 1 0 82892 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_895
timestamp 1644511149
transform 1 0 83444 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_897
timestamp 1644511149
transform 1 0 83628 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_909
timestamp 1644511149
transform 1 0 84732 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_921
timestamp 1644511149
transform 1 0 85836 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_933
timestamp 1644511149
transform 1 0 86940 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_945
timestamp 1644511149
transform 1 0 88044 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_951
timestamp 1644511149
transform 1 0 88596 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_953
timestamp 1644511149
transform 1 0 88780 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_965
timestamp 1644511149
transform 1 0 89884 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_977
timestamp 1644511149
transform 1 0 90988 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_989
timestamp 1644511149
transform 1 0 92092 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1001
timestamp 1644511149
transform 1 0 93196 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1007
timestamp 1644511149
transform 1 0 93748 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1009
timestamp 1644511149
transform 1 0 93932 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1021
timestamp 1644511149
transform 1 0 95036 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1033
timestamp 1644511149
transform 1 0 96140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1045
timestamp 1644511149
transform 1 0 97244 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1057
timestamp 1644511149
transform 1 0 98348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1063
timestamp 1644511149
transform 1 0 98900 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1065
timestamp 1644511149
transform 1 0 99084 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1077
timestamp 1644511149
transform 1 0 100188 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1089
timestamp 1644511149
transform 1 0 101292 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1101
timestamp 1644511149
transform 1 0 102396 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1113
timestamp 1644511149
transform 1 0 103500 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1119
timestamp 1644511149
transform 1 0 104052 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1121
timestamp 1644511149
transform 1 0 104236 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1133
timestamp 1644511149
transform 1 0 105340 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1145
timestamp 1644511149
transform 1 0 106444 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1157
timestamp 1644511149
transform 1 0 107548 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1169
timestamp 1644511149
transform 1 0 108652 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1175
timestamp 1644511149
transform 1 0 109204 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1177
timestamp 1644511149
transform 1 0 109388 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1189
timestamp 1644511149
transform 1 0 110492 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1201
timestamp 1644511149
transform 1 0 111596 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1213
timestamp 1644511149
transform 1 0 112700 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_1225
timestamp 1644511149
transform 1 0 113804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1231
timestamp 1644511149
transform 1 0 114356 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1233
timestamp 1644511149
transform 1 0 114540 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1245
timestamp 1644511149
transform 1 0 115644 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1257
timestamp 1644511149
transform 1 0 116748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1265
timestamp 1644511149
transform 1 0 117484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1273
timestamp 1644511149
transform 1 0 118220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1644511149
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1644511149
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1644511149
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_181
timestamp 1644511149
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1644511149
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_237
timestamp 1644511149
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1644511149
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1644511149
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_293
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1644511149
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_321
timestamp 1644511149
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1644511149
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1644511149
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_393
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_405
timestamp 1644511149
transform 1 0 38364 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1644511149
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_449
timestamp 1644511149
transform 1 0 42412 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_461
timestamp 1644511149
transform 1 0 43516 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_473
timestamp 1644511149
transform 1 0 44620 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_501
timestamp 1644511149
transform 1 0 47196 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_505
timestamp 1644511149
transform 1 0 47564 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_517
timestamp 1644511149
transform 1 0 48668 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_529
timestamp 1644511149
transform 1 0 49772 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_545
timestamp 1644511149
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_557
timestamp 1644511149
transform 1 0 52348 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_561
timestamp 1644511149
transform 1 0 52716 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_573
timestamp 1644511149
transform 1 0 53820 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_585
timestamp 1644511149
transform 1 0 54924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_601
timestamp 1644511149
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_613
timestamp 1644511149
transform 1 0 57500 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_617
timestamp 1644511149
transform 1 0 57868 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_629
timestamp 1644511149
transform 1 0 58972 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_641
timestamp 1644511149
transform 1 0 60076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_645
timestamp 1644511149
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_657
timestamp 1644511149
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_669
timestamp 1644511149
transform 1 0 62652 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_673
timestamp 1644511149
transform 1 0 63020 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_685
timestamp 1644511149
transform 1 0 64124 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_697
timestamp 1644511149
transform 1 0 65228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_701
timestamp 1644511149
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_713
timestamp 1644511149
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_725
timestamp 1644511149
transform 1 0 67804 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_729
timestamp 1644511149
transform 1 0 68172 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_741
timestamp 1644511149
transform 1 0 69276 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_753
timestamp 1644511149
transform 1 0 70380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_757
timestamp 1644511149
transform 1 0 70748 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_769
timestamp 1644511149
transform 1 0 71852 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_781
timestamp 1644511149
transform 1 0 72956 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_785
timestamp 1644511149
transform 1 0 73324 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_797
timestamp 1644511149
transform 1 0 74428 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_809
timestamp 1644511149
transform 1 0 75532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_813
timestamp 1644511149
transform 1 0 75900 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_825
timestamp 1644511149
transform 1 0 77004 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_837
timestamp 1644511149
transform 1 0 78108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_841
timestamp 1644511149
transform 1 0 78476 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_853
timestamp 1644511149
transform 1 0 79580 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_865
timestamp 1644511149
transform 1 0 80684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_869
timestamp 1644511149
transform 1 0 81052 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_881
timestamp 1644511149
transform 1 0 82156 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_893
timestamp 1644511149
transform 1 0 83260 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_897
timestamp 1644511149
transform 1 0 83628 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_909
timestamp 1644511149
transform 1 0 84732 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_921
timestamp 1644511149
transform 1 0 85836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_925
timestamp 1644511149
transform 1 0 86204 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_937
timestamp 1644511149
transform 1 0 87308 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_949
timestamp 1644511149
transform 1 0 88412 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_953
timestamp 1644511149
transform 1 0 88780 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_965
timestamp 1644511149
transform 1 0 89884 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_977
timestamp 1644511149
transform 1 0 90988 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_981
timestamp 1644511149
transform 1 0 91356 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_993
timestamp 1644511149
transform 1 0 92460 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1005
timestamp 1644511149
transform 1 0 93564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1009
timestamp 1644511149
transform 1 0 93932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1021
timestamp 1644511149
transform 1 0 95036 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1033
timestamp 1644511149
transform 1 0 96140 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1037
timestamp 1644511149
transform 1 0 96508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1049
timestamp 1644511149
transform 1 0 97612 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1061
timestamp 1644511149
transform 1 0 98716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1065
timestamp 1644511149
transform 1 0 99084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1077
timestamp 1644511149
transform 1 0 100188 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1089
timestamp 1644511149
transform 1 0 101292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1093
timestamp 1644511149
transform 1 0 101660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1105
timestamp 1644511149
transform 1 0 102764 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1117
timestamp 1644511149
transform 1 0 103868 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1121
timestamp 1644511149
transform 1 0 104236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1133
timestamp 1644511149
transform 1 0 105340 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1145
timestamp 1644511149
transform 1 0 106444 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1149
timestamp 1644511149
transform 1 0 106812 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1161
timestamp 1644511149
transform 1 0 107916 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1173
timestamp 1644511149
transform 1 0 109020 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1177
timestamp 1644511149
transform 1 0 109388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1189
timestamp 1644511149
transform 1 0 110492 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1201
timestamp 1644511149
transform 1 0 111596 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1205
timestamp 1644511149
transform 1 0 111964 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1217
timestamp 1644511149
transform 1 0 113068 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1229
timestamp 1644511149
transform 1 0 114172 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1233
timestamp 1644511149
transform 1 0 114540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1245
timestamp 1644511149
transform 1 0 115644 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1257
timestamp 1644511149
transform 1 0 116748 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1265
timestamp 1644511149
transform 1 0 117484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_1273
timestamp 1644511149
transform 1 0 118220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 118864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 118864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 118864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 118864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 118864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 118864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 118864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 118864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 118864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 118864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 118864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 118864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 118864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 118864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 118864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 118864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 118864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 118864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 118864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 118864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 118864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 118864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 118864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 118864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 118864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 118864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 118864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 118864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 118864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 118864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 118864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 118864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 118864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 118864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 118864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 118864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 118864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 118864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 118864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 118864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 118864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 118864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 118864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 118864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 118864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 118864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 118864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 118864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 118864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 118864 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 118864 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 118864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 118864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 118864 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 118864 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 118864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 118864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 118864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 118864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 118864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 118864 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 118864 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 118864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 118864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 118864 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 80960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 83536 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 86112 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 88688 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 91264 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 93840 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 96416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 98992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 101568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 104144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 106720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 109296 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 111872 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 114448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 117024 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 83536 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 88688 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 93840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 98992 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 104144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 109296 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 114448 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 80960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 86112 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 91264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 96416 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 101568 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 106720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 111872 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 117024 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 83536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 88688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 93840 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 98992 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 104144 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 109296 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 114448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 80960 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 86112 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 91264 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 96416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 101568 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 106720 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 111872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 117024 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 83536 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 88688 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 93840 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 98992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 104144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 109296 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 114448 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 80960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 86112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 91264 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 96416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 101568 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 106720 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 111872 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 117024 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 83536 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 88688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 93840 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 98992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 104144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 109296 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 114448 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 80960 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 86112 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 91264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 96416 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 101568 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 106720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 111872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 117024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 83536 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 88688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 93840 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 98992 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 104144 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 109296 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 114448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 80960 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 86112 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 91264 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 96416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 101568 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 106720 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 111872 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 117024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 83536 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 88688 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 93840 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 98992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 104144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 109296 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 114448 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 80960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 86112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 91264 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 96416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 101568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 106720 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 111872 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 117024 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 83536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 88688 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 93840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 98992 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 104144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 109296 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 114448 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 80960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 86112 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 91264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 96416 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 101568 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 106720 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 111872 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 117024 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 83536 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 88688 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 93840 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 98992 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 104144 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 109296 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 114448 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 80960 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 86112 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 91264 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 96416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 101568 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 106720 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 111872 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 117024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 83536 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 88688 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 93840 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 98992 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 104144 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 109296 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 114448 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 80960 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 86112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 91264 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 96416 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 101568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 106720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 111872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 117024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 83536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 88688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 93840 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 98992 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 104144 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 109296 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 114448 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 80960 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 86112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 91264 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 96416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 101568 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 106720 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 111872 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 117024 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 83536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 88688 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 93840 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 98992 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 104144 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 109296 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 114448 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 80960 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 86112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 91264 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 96416 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 101568 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 106720 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 111872 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 117024 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 83536 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 88688 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 93840 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 98992 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 104144 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 109296 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 114448 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 80960 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 86112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 91264 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 96416 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 101568 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 106720 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 111872 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 117024 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 83536 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 88688 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 93840 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 98992 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 104144 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 109296 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 114448 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 80960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 86112 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 91264 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 96416 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 101568 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 106720 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 111872 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 117024 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 83536 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 88688 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 93840 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 98992 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 104144 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 109296 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 114448 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 70656 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 75808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 80960 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 86112 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 91264 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 96416 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 101568 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 106720 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 111872 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 117024 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 73232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 78384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 83536 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 88688 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 93840 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 98992 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 104144 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 109296 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 114448 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 70656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 75808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 80960 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 86112 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 91264 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 96416 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 101568 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 106720 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 111872 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 117024 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 73232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 78384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 83536 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 88688 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 93840 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 98992 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 104144 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 109296 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 114448 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 70656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 75808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 80960 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 86112 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 91264 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 96416 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 101568 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 106720 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 111872 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 117024 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 73232 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 78384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 83536 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 88688 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 93840 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 98992 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 104144 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 109296 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 114448 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 70656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 75808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 80960 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 86112 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 91264 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 96416 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 101568 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 106720 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 111872 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 117024 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 73232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 78384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 83536 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 88688 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 93840 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 98992 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 104144 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 109296 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 114448 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1644511149
transform 1 0 70656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1644511149
transform 1 0 75808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1644511149
transform 1 0 80960 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1644511149
transform 1 0 86112 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1644511149
transform 1 0 91264 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1644511149
transform 1 0 96416 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1644511149
transform 1 0 101568 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1644511149
transform 1 0 106720 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1644511149
transform 1 0 111872 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1644511149
transform 1 0 117024 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1644511149
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1644511149
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1644511149
transform 1 0 73232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1644511149
transform 1 0 78384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1644511149
transform 1 0 83536 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1644511149
transform 1 0 88688 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1644511149
transform 1 0 93840 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1644511149
transform 1 0 98992 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1644511149
transform 1 0 104144 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1644511149
transform 1 0 109296 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1644511149
transform 1 0 114448 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1644511149
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1644511149
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1644511149
transform 1 0 70656 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1644511149
transform 1 0 75808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1644511149
transform 1 0 80960 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1644511149
transform 1 0 86112 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1644511149
transform 1 0 91264 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1644511149
transform 1 0 96416 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1644511149
transform 1 0 101568 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1644511149
transform 1 0 106720 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1644511149
transform 1 0 111872 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1644511149
transform 1 0 117024 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1644511149
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1644511149
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1644511149
transform 1 0 73232 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1644511149
transform 1 0 78384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1644511149
transform 1 0 83536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1644511149
transform 1 0 88688 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1644511149
transform 1 0 93840 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1644511149
transform 1 0 98992 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1644511149
transform 1 0 104144 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1644511149
transform 1 0 109296 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1644511149
transform 1 0 114448 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1644511149
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1644511149
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1644511149
transform 1 0 70656 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1644511149
transform 1 0 75808 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1644511149
transform 1 0 80960 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1644511149
transform 1 0 86112 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1644511149
transform 1 0 91264 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1644511149
transform 1 0 96416 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1644511149
transform 1 0 101568 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1644511149
transform 1 0 106720 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1644511149
transform 1 0 111872 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1644511149
transform 1 0 117024 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1644511149
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1644511149
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1644511149
transform 1 0 73232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1644511149
transform 1 0 78384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1644511149
transform 1 0 83536 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1644511149
transform 1 0 88688 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1644511149
transform 1 0 93840 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1644511149
transform 1 0 98992 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1644511149
transform 1 0 104144 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1644511149
transform 1 0 109296 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1644511149
transform 1 0 114448 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1644511149
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1644511149
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1644511149
transform 1 0 70656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1644511149
transform 1 0 75808 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1644511149
transform 1 0 80960 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1644511149
transform 1 0 86112 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1644511149
transform 1 0 91264 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1644511149
transform 1 0 96416 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1644511149
transform 1 0 101568 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1644511149
transform 1 0 106720 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1644511149
transform 1 0 111872 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1644511149
transform 1 0 117024 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1644511149
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1644511149
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1644511149
transform 1 0 73232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1644511149
transform 1 0 78384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1644511149
transform 1 0 83536 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1644511149
transform 1 0 88688 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1644511149
transform 1 0 93840 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1644511149
transform 1 0 98992 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1644511149
transform 1 0 104144 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1644511149
transform 1 0 109296 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1644511149
transform 1 0 114448 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1644511149
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1644511149
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1644511149
transform 1 0 70656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1644511149
transform 1 0 75808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1644511149
transform 1 0 80960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1644511149
transform 1 0 86112 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1644511149
transform 1 0 91264 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1644511149
transform 1 0 96416 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1644511149
transform 1 0 101568 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1644511149
transform 1 0 106720 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1644511149
transform 1 0 111872 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1644511149
transform 1 0 117024 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1644511149
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1644511149
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1644511149
transform 1 0 73232 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1644511149
transform 1 0 78384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1644511149
transform 1 0 83536 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1644511149
transform 1 0 88688 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1644511149
transform 1 0 93840 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1644511149
transform 1 0 98992 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1644511149
transform 1 0 104144 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1644511149
transform 1 0 109296 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1644511149
transform 1 0 114448 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1644511149
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1644511149
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1644511149
transform 1 0 70656 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1644511149
transform 1 0 75808 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1644511149
transform 1 0 80960 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1644511149
transform 1 0 86112 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1644511149
transform 1 0 91264 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1644511149
transform 1 0 96416 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1644511149
transform 1 0 101568 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1644511149
transform 1 0 106720 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1644511149
transform 1 0 111872 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1644511149
transform 1 0 117024 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1644511149
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1644511149
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1644511149
transform 1 0 73232 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1644511149
transform 1 0 78384 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1644511149
transform 1 0 83536 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1644511149
transform 1 0 88688 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1644511149
transform 1 0 93840 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1644511149
transform 1 0 98992 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1644511149
transform 1 0 104144 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1644511149
transform 1 0 109296 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1644511149
transform 1 0 114448 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1644511149
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1644511149
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1644511149
transform 1 0 70656 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1644511149
transform 1 0 75808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1644511149
transform 1 0 80960 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1644511149
transform 1 0 86112 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1644511149
transform 1 0 91264 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1644511149
transform 1 0 96416 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1644511149
transform 1 0 101568 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1644511149
transform 1 0 106720 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1644511149
transform 1 0 111872 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1644511149
transform 1 0 117024 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1644511149
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1644511149
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1644511149
transform 1 0 73232 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1644511149
transform 1 0 78384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1644511149
transform 1 0 83536 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1644511149
transform 1 0 88688 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1644511149
transform 1 0 93840 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1644511149
transform 1 0 98992 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1644511149
transform 1 0 104144 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1644511149
transform 1 0 109296 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1644511149
transform 1 0 114448 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1644511149
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1644511149
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1644511149
transform 1 0 70656 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1644511149
transform 1 0 75808 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1644511149
transform 1 0 80960 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1644511149
transform 1 0 86112 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1644511149
transform 1 0 91264 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1644511149
transform 1 0 96416 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1644511149
transform 1 0 101568 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1644511149
transform 1 0 106720 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1644511149
transform 1 0 111872 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1644511149
transform 1 0 117024 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1644511149
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1644511149
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1644511149
transform 1 0 73232 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1644511149
transform 1 0 78384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1644511149
transform 1 0 83536 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1644511149
transform 1 0 88688 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1644511149
transform 1 0 93840 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1644511149
transform 1 0 98992 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1644511149
transform 1 0 104144 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1644511149
transform 1 0 109296 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1644511149
transform 1 0 114448 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1644511149
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1644511149
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1644511149
transform 1 0 70656 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1644511149
transform 1 0 75808 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1644511149
transform 1 0 80960 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1644511149
transform 1 0 86112 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1644511149
transform 1 0 91264 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1644511149
transform 1 0 96416 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1644511149
transform 1 0 101568 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1644511149
transform 1 0 106720 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1644511149
transform 1 0 111872 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1644511149
transform 1 0 117024 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1644511149
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1644511149
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1644511149
transform 1 0 73232 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1644511149
transform 1 0 78384 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1644511149
transform 1 0 83536 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1644511149
transform 1 0 88688 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1644511149
transform 1 0 93840 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1644511149
transform 1 0 98992 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1644511149
transform 1 0 104144 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1644511149
transform 1 0 109296 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1644511149
transform 1 0 114448 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1644511149
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1644511149
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1644511149
transform 1 0 70656 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1644511149
transform 1 0 75808 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1644511149
transform 1 0 80960 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1644511149
transform 1 0 86112 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1644511149
transform 1 0 91264 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1644511149
transform 1 0 96416 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1644511149
transform 1 0 101568 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1644511149
transform 1 0 106720 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1644511149
transform 1 0 111872 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1644511149
transform 1 0 117024 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1644511149
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1644511149
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1644511149
transform 1 0 73232 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1644511149
transform 1 0 78384 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1644511149
transform 1 0 83536 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1644511149
transform 1 0 88688 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1644511149
transform 1 0 93840 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1644511149
transform 1 0 98992 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1644511149
transform 1 0 104144 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1644511149
transform 1 0 109296 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1644511149
transform 1 0 114448 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1644511149
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1644511149
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1644511149
transform 1 0 70656 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1644511149
transform 1 0 75808 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1644511149
transform 1 0 80960 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1644511149
transform 1 0 86112 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1644511149
transform 1 0 91264 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1644511149
transform 1 0 96416 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1644511149
transform 1 0 101568 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1644511149
transform 1 0 106720 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1644511149
transform 1 0 111872 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1644511149
transform 1 0 117024 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1644511149
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1644511149
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1644511149
transform 1 0 73232 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1644511149
transform 1 0 78384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1644511149
transform 1 0 83536 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1644511149
transform 1 0 88688 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1644511149
transform 1 0 93840 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1644511149
transform 1 0 98992 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1644511149
transform 1 0 104144 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1644511149
transform 1 0 109296 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1644511149
transform 1 0 114448 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1644511149
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1644511149
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1644511149
transform 1 0 70656 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1644511149
transform 1 0 75808 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1644511149
transform 1 0 80960 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1644511149
transform 1 0 86112 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1644511149
transform 1 0 91264 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1644511149
transform 1 0 96416 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1644511149
transform 1 0 101568 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1644511149
transform 1 0 106720 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1644511149
transform 1 0 111872 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1644511149
transform 1 0 117024 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1644511149
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1644511149
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1644511149
transform 1 0 73232 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1644511149
transform 1 0 78384 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1644511149
transform 1 0 83536 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1644511149
transform 1 0 88688 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1644511149
transform 1 0 93840 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1644511149
transform 1 0 98992 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1644511149
transform 1 0 104144 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1644511149
transform 1 0 109296 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1644511149
transform 1 0 114448 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1644511149
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1644511149
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1644511149
transform 1 0 70656 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1644511149
transform 1 0 75808 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1644511149
transform 1 0 80960 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1644511149
transform 1 0 86112 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1644511149
transform 1 0 91264 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1644511149
transform 1 0 96416 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1644511149
transform 1 0 101568 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1644511149
transform 1 0 106720 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1644511149
transform 1 0 111872 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1644511149
transform 1 0 117024 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1644511149
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1644511149
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1644511149
transform 1 0 73232 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1644511149
transform 1 0 78384 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1644511149
transform 1 0 83536 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1644511149
transform 1 0 88688 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1644511149
transform 1 0 93840 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1644511149
transform 1 0 98992 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1644511149
transform 1 0 104144 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1644511149
transform 1 0 109296 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1644511149
transform 1 0 114448 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1644511149
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1644511149
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1644511149
transform 1 0 70656 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1644511149
transform 1 0 75808 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1644511149
transform 1 0 80960 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1644511149
transform 1 0 86112 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1644511149
transform 1 0 91264 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1644511149
transform 1 0 96416 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1644511149
transform 1 0 101568 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1644511149
transform 1 0 106720 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1644511149
transform 1 0 111872 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1644511149
transform 1 0 117024 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1644511149
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1644511149
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1644511149
transform 1 0 73232 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1644511149
transform 1 0 78384 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1644511149
transform 1 0 83536 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1644511149
transform 1 0 88688 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1644511149
transform 1 0 93840 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1644511149
transform 1 0 98992 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1644511149
transform 1 0 104144 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1644511149
transform 1 0 109296 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1644511149
transform 1 0 114448 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1644511149
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1644511149
transform 1 0 52624 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1644511149
transform 1 0 57776 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1644511149
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1644511149
transform 1 0 62928 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1644511149
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1644511149
transform 1 0 68080 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1644511149
transform 1 0 70656 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1644511149
transform 1 0 73232 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1644511149
transform 1 0 75808 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1644511149
transform 1 0 78384 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1644511149
transform 1 0 80960 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1644511149
transform 1 0 83536 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1644511149
transform 1 0 86112 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1644511149
transform 1 0 88688 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1644511149
transform 1 0 91264 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1644511149
transform 1 0 93840 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1644511149
transform 1 0 96416 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1644511149
transform 1 0 98992 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1644511149
transform 1 0 101568 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1644511149
transform 1 0 104144 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1644511149
transform 1 0 106720 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1644511149
transform 1 0 109296 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1644511149
transform 1 0 111872 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1644511149
transform 1 0 114448 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1644511149
transform 1 0 117024 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _039_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 100280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _040_
timestamp 1644511149
transform 1 0 108560 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _041_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 105064 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _042_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 105800 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _043_
timestamp 1644511149
transform 1 0 105616 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _044_
timestamp 1644511149
transform 1 0 106812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _045_
timestamp 1644511149
transform 1 0 107272 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _046_
timestamp 1644511149
transform 1 0 108284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _047_
timestamp 1644511149
transform 1 0 109388 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _048_
timestamp 1644511149
transform 1 0 110584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _049_
timestamp 1644511149
transform 1 0 109388 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _050_
timestamp 1644511149
transform 1 0 111688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _051_
timestamp 1644511149
transform 1 0 112424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _052_
timestamp 1644511149
transform 1 0 111964 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _053_
timestamp 1644511149
transform 1 0 115092 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _054_
timestamp 1644511149
transform 1 0 113252 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _055_
timestamp 1644511149
transform 1 0 115828 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _056_
timestamp 1644511149
transform 1 0 114908 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1644511149
transform 1 0 116564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _058_
timestamp 1644511149
transform 1 0 115828 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1644511149
transform 1 0 116196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _060_
timestamp 1644511149
transform 1 0 115736 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1644511149
transform 1 0 114724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1644511149
transform 1 0 98256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _063_
timestamp 1644511149
transform 1 0 99084 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _064_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 98716 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _065_
timestamp 1644511149
transform 1 0 74612 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1644511149
transform 1 0 75900 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _067_
timestamp 1644511149
transform 1 0 75900 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _068_
timestamp 1644511149
transform 1 0 76452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _069_
timestamp 1644511149
transform 1 0 77188 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _070_
timestamp 1644511149
transform 1 0 78476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _071_
timestamp 1644511149
transform 1 0 78660 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _072_
timestamp 1644511149
transform 1 0 79396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1644511149
transform 1 0 87400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 1644511149
transform 1 0 81052 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _075_
timestamp 1644511149
transform 1 0 81512 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp 1644511149
transform 1 0 82616 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _077_
timestamp 1644511149
transform 1 0 82432 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _078_
timestamp 1644511149
transform 1 0 83628 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _079_
timestamp 1644511149
transform 1 0 83628 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _080_
timestamp 1644511149
transform 1 0 84824 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _081_
timestamp 1644511149
transform 1 0 85008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _082_
timestamp 1644511149
transform 1 0 86204 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _083_
timestamp 1644511149
transform 1 0 86480 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _084_
timestamp 1644511149
transform 1 0 88780 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _085_
timestamp 1644511149
transform 1 0 87492 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1644511149
transform 1 0 88780 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _087_
timestamp 1644511149
transform 1 0 88780 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1644511149
transform 1 0 89240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _089_
timestamp 1644511149
transform 1 0 90068 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1644511149
transform 1 0 90804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _091_
timestamp 1644511149
transform 1 0 91540 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1644511149
transform 1 0 92184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _093_
timestamp 1644511149
transform 1 0 92184 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1644511149
transform 1 0 92920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _095_
timestamp 1644511149
transform 1 0 97520 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _096_
timestamp 1644511149
transform 1 0 95036 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1644511149
transform 1 0 95772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _098_
timestamp 1644511149
transform 1 0 96508 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1644511149
transform 1 0 96508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _100_
timestamp 1644511149
transform 1 0 97704 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1644511149
transform 1 0 97888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _102_
timestamp 1644511149
transform 1 0 99084 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1644511149
transform 1 0 99636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _104_
timestamp 1644511149
transform 1 0 100280 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1644511149
transform 1 0 100372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _106_
timestamp 1644511149
transform 1 0 101660 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1644511149
transform 1 0 102212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _108_
timestamp 1644511149
transform 1 0 102856 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1644511149
transform 1 0 104236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _110_
timestamp 1644511149
transform 1 0 60904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _111_
timestamp 1644511149
transform 1 0 63020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _112_
timestamp 1644511149
transform 1 0 63940 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _113_
timestamp 1644511149
transform 1 0 65596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _114_
timestamp 1644511149
transform 1 0 66608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _115_
timestamp 1644511149
transform 1 0 68172 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _116_
timestamp 1644511149
transform 1 0 69460 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _117_
timestamp 1644511149
transform 1 0 70932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _118_
timestamp 1644511149
transform 1 0 72312 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _119_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 61456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1644511149
transform 1 0 62928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1644511149
transform 1 0 64676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1644511149
transform 1 0 65780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1644511149
transform 1 0 67160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1644511149
transform 1 0 68632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1644511149
transform 1 0 70012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1644511149
transform 1 0 71484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1644511149
transform 1 0 73324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _128_
timestamp 1644511149
transform 1 0 59432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1644511149
transform 1 0 60076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 1644511149
transform 1 0 117668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 117668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1644511149
transform 1 0 117668 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 1644511149
transform 1 0 117668 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input5
timestamp 1644511149
transform 1 0 117668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1644511149
transform 1 0 117668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1644511149
transform 1 0 117668 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1644511149
transform 1 0 117668 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 1644511149
transform 1 0 117668 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1644511149
transform 1 0 117668 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input11 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 116472 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input12
timestamp 1644511149
transform 1 0 14996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input13
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 1644511149
transform 1 0 30728 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input16
timestamp 1644511149
transform 1 0 33580 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1644511149
transform 1 0 35052 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input18
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input20
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input21
timestamp 1644511149
transform 1 0 40756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input22
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1644511149
transform 1 0 46368 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input27
timestamp 1644511149
transform 1 0 47840 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input28
timestamp 1644511149
transform 1 0 49128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input29
timestamp 1644511149
transform 1 0 50692 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input30
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input31
timestamp 1644511149
transform 1 0 53636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input32
timestamp 1644511149
transform 1 0 55292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 1644511149
transform 1 0 56396 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input34
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input35
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 1644511149
transform 1 0 59248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input37
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input39
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input41
timestamp 1644511149
transform 1 0 25300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input42
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input43
timestamp 1644511149
transform 1 0 27876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1644511149
transform 1 0 74980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1644511149
transform 1 0 89516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1644511149
transform 1 0 90712 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1644511149
transform 1 0 91540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1644511149
transform 1 0 93932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 94944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 96508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform 1 0 97796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1644511149
transform 1 0 101016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1644511149
transform 1 0 100648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1644511149
transform 1 0 102948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1644511149
transform 1 0 76360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 104236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1644511149
transform 1 0 104788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1644511149
transform 1 0 106812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1644511149
transform 1 0 107640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1644511149
transform 1 0 110584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1644511149
transform 1 0 111044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform 1 0 112056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1644511149
transform 1 0 113528 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1644511149
transform 1 0 114908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1644511149
transform 1 0 117024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1644511149
transform 1 0 77740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1644511149
transform 1 0 117760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 117300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1644511149
transform 1 0 79856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1644511149
transform 1 0 80684 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1644511149
transform 1 0 82064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1644511149
transform 1 0 83536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1644511149
transform 1 0 84916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1644511149
transform 1 0 86388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1644511149
transform 1 0 87768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 6440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform 1 0 62100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 63572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 64860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 66240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform 1 0 69092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform 1 0 70656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 72128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform 1 0 73508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform 1 0 60720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform 1 0 117852 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1644511149
transform 1 0 117852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1644511149
transform 1 0 117852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1644511149
transform 1 0 117852 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1644511149
transform 1 0 117852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1644511149
transform 1 0 117852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1644511149
transform 1 0 117852 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1644511149
transform 1 0 117852 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1644511149
transform 1 0 117852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1644511149
transform 1 0 117852 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1644511149
transform 1 0 117852 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1644511149
transform 1 0 117852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1644511149
transform 1 0 117852 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1644511149
transform 1 0 117852 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1644511149
transform 1 0 117852 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1644511149
transform 1 0 117852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1644511149
transform 1 0 117852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1644511149
transform 1 0 117852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1644511149
transform 1 0 117852 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1644511149
transform 1 0 117852 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1644511149
transform 1 0 117852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1644511149
transform 1 0 117852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1644511149
transform 1 0 117852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1644511149
transform 1 0 117116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1644511149
transform 1 0 117116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1644511149
transform 1 0 117852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1644511149
transform 1 0 117852 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1644511149
transform 1 0 117852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1644511149
transform 1 0 117852 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1644511149
transform 1 0 117852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1644511149
transform 1 0 117852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1644511149
transform 1 0 117852 0 -1 19584
box -38 -48 406 592
<< labels >>
rlabel metal3 s 119200 1232 120000 1352 6 addr[0]
port 0 nsew signal input
rlabel metal3 s 119200 2184 120000 2304 6 addr[1]
port 1 nsew signal input
rlabel metal3 s 119200 3136 120000 3256 6 addr[2]
port 2 nsew signal input
rlabel metal3 s 119200 4088 120000 4208 6 addr[3]
port 3 nsew signal input
rlabel metal3 s 119200 5040 120000 5160 6 addr[4]
port 4 nsew signal input
rlabel metal3 s 119200 5992 120000 6112 6 addr[5]
port 5 nsew signal input
rlabel metal3 s 119200 6808 120000 6928 6 addr[6]
port 6 nsew signal input
rlabel metal3 s 119200 7760 120000 7880 6 addr[7]
port 7 nsew signal input
rlabel metal3 s 119200 8712 120000 8832 6 addr[8]
port 8 nsew signal input
rlabel metal3 s 119200 9664 120000 9784 6 addr[9]
port 9 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 addr_mem0[0]
port 10 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 addr_mem0[1]
port 11 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 addr_mem0[2]
port 12 nsew signal tristate
rlabel metal2 s 6366 0 6422 800 6 addr_mem0[3]
port 13 nsew signal tristate
rlabel metal2 s 7746 0 7802 800 6 addr_mem0[4]
port 14 nsew signal tristate
rlabel metal2 s 9218 0 9274 800 6 addr_mem0[5]
port 15 nsew signal tristate
rlabel metal2 s 10598 0 10654 800 6 addr_mem0[6]
port 16 nsew signal tristate
rlabel metal2 s 12070 0 12126 800 6 addr_mem0[7]
port 17 nsew signal tristate
rlabel metal2 s 13450 0 13506 800 6 addr_mem0[8]
port 18 nsew signal tristate
rlabel metal2 s 62026 0 62082 800 6 addr_mem1[0]
port 19 nsew signal tristate
rlabel metal2 s 63498 0 63554 800 6 addr_mem1[1]
port 20 nsew signal tristate
rlabel metal2 s 64878 0 64934 800 6 addr_mem1[2]
port 21 nsew signal tristate
rlabel metal2 s 66350 0 66406 800 6 addr_mem1[3]
port 22 nsew signal tristate
rlabel metal2 s 67730 0 67786 800 6 addr_mem1[4]
port 23 nsew signal tristate
rlabel metal2 s 69202 0 69258 800 6 addr_mem1[5]
port 24 nsew signal tristate
rlabel metal2 s 70582 0 70638 800 6 addr_mem1[6]
port 25 nsew signal tristate
rlabel metal2 s 72054 0 72110 800 6 addr_mem1[7]
port 26 nsew signal tristate
rlabel metal2 s 73434 0 73490 800 6 addr_mem1[8]
port 27 nsew signal tristate
rlabel metal3 s 119200 416 120000 536 6 csb
port 28 nsew signal input
rlabel metal2 s 662 0 718 800 6 csb_mem0
port 29 nsew signal tristate
rlabel metal2 s 60646 0 60702 800 6 csb_mem1
port 30 nsew signal tristate
rlabel metal3 s 119200 10616 120000 10736 6 dout[0]
port 31 nsew signal tristate
rlabel metal3 s 119200 19864 120000 19984 6 dout[10]
port 32 nsew signal tristate
rlabel metal3 s 119200 20816 120000 20936 6 dout[11]
port 33 nsew signal tristate
rlabel metal3 s 119200 21768 120000 21888 6 dout[12]
port 34 nsew signal tristate
rlabel metal3 s 119200 22720 120000 22840 6 dout[13]
port 35 nsew signal tristate
rlabel metal3 s 119200 23536 120000 23656 6 dout[14]
port 36 nsew signal tristate
rlabel metal3 s 119200 24488 120000 24608 6 dout[15]
port 37 nsew signal tristate
rlabel metal3 s 119200 25440 120000 25560 6 dout[16]
port 38 nsew signal tristate
rlabel metal3 s 119200 26392 120000 26512 6 dout[17]
port 39 nsew signal tristate
rlabel metal3 s 119200 27344 120000 27464 6 dout[18]
port 40 nsew signal tristate
rlabel metal3 s 119200 28296 120000 28416 6 dout[19]
port 41 nsew signal tristate
rlabel metal3 s 119200 11568 120000 11688 6 dout[1]
port 42 nsew signal tristate
rlabel metal3 s 119200 29112 120000 29232 6 dout[20]
port 43 nsew signal tristate
rlabel metal3 s 119200 30064 120000 30184 6 dout[21]
port 44 nsew signal tristate
rlabel metal3 s 119200 31016 120000 31136 6 dout[22]
port 45 nsew signal tristate
rlabel metal3 s 119200 31968 120000 32088 6 dout[23]
port 46 nsew signal tristate
rlabel metal3 s 119200 32920 120000 33040 6 dout[24]
port 47 nsew signal tristate
rlabel metal3 s 119200 33872 120000 33992 6 dout[25]
port 48 nsew signal tristate
rlabel metal3 s 119200 34688 120000 34808 6 dout[26]
port 49 nsew signal tristate
rlabel metal3 s 119200 35640 120000 35760 6 dout[27]
port 50 nsew signal tristate
rlabel metal3 s 119200 36592 120000 36712 6 dout[28]
port 51 nsew signal tristate
rlabel metal3 s 119200 37544 120000 37664 6 dout[29]
port 52 nsew signal tristate
rlabel metal3 s 119200 12384 120000 12504 6 dout[2]
port 53 nsew signal tristate
rlabel metal3 s 119200 38496 120000 38616 6 dout[30]
port 54 nsew signal tristate
rlabel metal3 s 119200 39448 120000 39568 6 dout[31]
port 55 nsew signal tristate
rlabel metal3 s 119200 13336 120000 13456 6 dout[3]
port 56 nsew signal tristate
rlabel metal3 s 119200 14288 120000 14408 6 dout[4]
port 57 nsew signal tristate
rlabel metal3 s 119200 15240 120000 15360 6 dout[5]
port 58 nsew signal tristate
rlabel metal3 s 119200 16192 120000 16312 6 dout[6]
port 59 nsew signal tristate
rlabel metal3 s 119200 17144 120000 17264 6 dout[7]
port 60 nsew signal tristate
rlabel metal3 s 119200 17960 120000 18080 6 dout[8]
port 61 nsew signal tristate
rlabel metal3 s 119200 18912 120000 19032 6 dout[9]
port 62 nsew signal tristate
rlabel metal2 s 14922 0 14978 800 6 dout_mem0[0]
port 63 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 dout_mem0[10]
port 64 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 dout_mem0[11]
port 65 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 dout_mem0[12]
port 66 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 dout_mem0[13]
port 67 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 dout_mem0[14]
port 68 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 dout_mem0[15]
port 69 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 dout_mem0[16]
port 70 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 dout_mem0[17]
port 71 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 dout_mem0[18]
port 72 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 dout_mem0[19]
port 73 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 dout_mem0[1]
port 74 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 dout_mem0[20]
port 75 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 dout_mem0[21]
port 76 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 dout_mem0[22]
port 77 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 dout_mem0[23]
port 78 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 dout_mem0[24]
port 79 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 dout_mem0[25]
port 80 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 dout_mem0[26]
port 81 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 dout_mem0[27]
port 82 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 dout_mem0[28]
port 83 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 dout_mem0[29]
port 84 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 dout_mem0[2]
port 85 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 dout_mem0[30]
port 86 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 dout_mem0[31]
port 87 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 dout_mem0[3]
port 88 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 dout_mem0[4]
port 89 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 dout_mem0[5]
port 90 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 dout_mem0[6]
port 91 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 dout_mem0[7]
port 92 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 dout_mem0[8]
port 93 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 dout_mem0[9]
port 94 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 dout_mem1[0]
port 95 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 dout_mem1[10]
port 96 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 dout_mem1[11]
port 97 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 dout_mem1[12]
port 98 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 dout_mem1[13]
port 99 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 dout_mem1[14]
port 100 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 dout_mem1[15]
port 101 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 dout_mem1[16]
port 102 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 dout_mem1[17]
port 103 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 dout_mem1[18]
port 104 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 dout_mem1[19]
port 105 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 dout_mem1[1]
port 106 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 dout_mem1[20]
port 107 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 dout_mem1[21]
port 108 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 dout_mem1[22]
port 109 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 dout_mem1[23]
port 110 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 dout_mem1[24]
port 111 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 dout_mem1[25]
port 112 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 dout_mem1[26]
port 113 nsew signal input
rlabel metal2 s 113454 0 113510 800 6 dout_mem1[27]
port 114 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 dout_mem1[28]
port 115 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 dout_mem1[29]
port 116 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 dout_mem1[2]
port 117 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 dout_mem1[30]
port 118 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 dout_mem1[31]
port 119 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 dout_mem1[3]
port 120 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 dout_mem1[4]
port 121 nsew signal input
rlabel metal2 s 81990 0 82046 800 6 dout_mem1[5]
port 122 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 dout_mem1[6]
port 123 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 dout_mem1[7]
port 124 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 dout_mem1[8]
port 125 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 dout_mem1[9]
port 126 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 127 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 127 nsew power input
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 127 nsew power input
rlabel metal4 s 96368 2128 96688 37584 6 vccd1
port 127 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 128 nsew ground input
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 128 nsew ground input
rlabel metal4 s 81008 2128 81328 37584 6 vssd1
port 128 nsew ground input
rlabel metal4 s 111728 2128 112048 37584 6 vssd1
port 128 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 120000 40000
<< end >>
