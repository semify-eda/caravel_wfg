* NGSPICE file created from wfg_top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

.subckt wfg_top addr1[0] addr1[1] addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7]
+ addr1[8] addr1[9] csb1 dout1[0] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14]
+ dout1[15] dout1[16] dout1[17] dout1[18] dout1[19] dout1[1] dout1[20] dout1[21] dout1[22]
+ dout1[23] dout1[24] dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[2] dout1[30]
+ dout1[31] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7] dout1[8] dout1[9] io_oeb[0]
+ io_oeb[10] io_oeb[1] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_wbs_ack io_wbs_adr[0] io_wbs_adr[10] io_wbs_adr[11] io_wbs_adr[12]
+ io_wbs_adr[13] io_wbs_adr[14] io_wbs_adr[15] io_wbs_adr[16] io_wbs_adr[17] io_wbs_adr[18]
+ io_wbs_adr[19] io_wbs_adr[1] io_wbs_adr[20] io_wbs_adr[21] io_wbs_adr[22] io_wbs_adr[23]
+ io_wbs_adr[24] io_wbs_adr[25] io_wbs_adr[26] io_wbs_adr[27] io_wbs_adr[28] io_wbs_adr[29]
+ io_wbs_adr[2] io_wbs_adr[30] io_wbs_adr[31] io_wbs_adr[3] io_wbs_adr[4] io_wbs_adr[5]
+ io_wbs_adr[6] io_wbs_adr[7] io_wbs_adr[8] io_wbs_adr[9] io_wbs_clk io_wbs_cyc io_wbs_datrd[0]
+ io_wbs_datrd[10] io_wbs_datrd[11] io_wbs_datrd[12] io_wbs_datrd[13] io_wbs_datrd[14]
+ io_wbs_datrd[15] io_wbs_datrd[16] io_wbs_datrd[17] io_wbs_datrd[18] io_wbs_datrd[19]
+ io_wbs_datrd[1] io_wbs_datrd[20] io_wbs_datrd[21] io_wbs_datrd[22] io_wbs_datrd[23]
+ io_wbs_datrd[24] io_wbs_datrd[25] io_wbs_datrd[26] io_wbs_datrd[27] io_wbs_datrd[28]
+ io_wbs_datrd[29] io_wbs_datrd[2] io_wbs_datrd[30] io_wbs_datrd[31] io_wbs_datrd[3]
+ io_wbs_datrd[4] io_wbs_datrd[5] io_wbs_datrd[6] io_wbs_datrd[7] io_wbs_datrd[8]
+ io_wbs_datrd[9] io_wbs_datwr[0] io_wbs_datwr[10] io_wbs_datwr[11] io_wbs_datwr[12]
+ io_wbs_datwr[13] io_wbs_datwr[14] io_wbs_datwr[15] io_wbs_datwr[16] io_wbs_datwr[17]
+ io_wbs_datwr[18] io_wbs_datwr[19] io_wbs_datwr[1] io_wbs_datwr[20] io_wbs_datwr[21]
+ io_wbs_datwr[22] io_wbs_datwr[23] io_wbs_datwr[24] io_wbs_datwr[25] io_wbs_datwr[26]
+ io_wbs_datwr[27] io_wbs_datwr[28] io_wbs_datwr[29] io_wbs_datwr[2] io_wbs_datwr[30]
+ io_wbs_datwr[31] io_wbs_datwr[3] io_wbs_datwr[4] io_wbs_datwr[5] io_wbs_datwr[6]
+ io_wbs_datwr[7] io_wbs_datwr[8] io_wbs_datwr[9] io_wbs_rst io_wbs_stb io_wbs_we
+ vccd1 vssd1 wfg_drive_pat_dout_o[0] wfg_drive_pat_dout_o[10] wfg_drive_pat_dout_o[11]
+ wfg_drive_pat_dout_o[12] wfg_drive_pat_dout_o[13] wfg_drive_pat_dout_o[14] wfg_drive_pat_dout_o[15]
+ wfg_drive_pat_dout_o[16] wfg_drive_pat_dout_o[17] wfg_drive_pat_dout_o[18] wfg_drive_pat_dout_o[19]
+ wfg_drive_pat_dout_o[1] wfg_drive_pat_dout_o[20] wfg_drive_pat_dout_o[21] wfg_drive_pat_dout_o[22]
+ wfg_drive_pat_dout_o[23] wfg_drive_pat_dout_o[24] wfg_drive_pat_dout_o[25] wfg_drive_pat_dout_o[26]
+ wfg_drive_pat_dout_o[27] wfg_drive_pat_dout_o[28] wfg_drive_pat_dout_o[29] wfg_drive_pat_dout_o[2]
+ wfg_drive_pat_dout_o[30] wfg_drive_pat_dout_o[31] wfg_drive_pat_dout_o[3] wfg_drive_pat_dout_o[4]
+ wfg_drive_pat_dout_o[5] wfg_drive_pat_dout_o[6] wfg_drive_pat_dout_o[7] wfg_drive_pat_dout_o[8]
+ wfg_drive_pat_dout_o[9] wfg_drive_spi_cs_no wfg_drive_spi_sclk_o wfg_drive_spi_sdo_o
XFILLER_95_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06883_ _06880_/Y _13778_/Q _13775_/Q _06881_/Y _06882_/Y vssd1 vssd1 vccd1 vccd1
+ _06883_/X sky130_fd_sc_hd__a221o_1
X_09671_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09673_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08622_ _08622_/A _08893_/A vssd1 vssd1 vccd1 vccd1 _08626_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08553_ _14017_/Q vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__buf_2
XFILLER_39_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07504_ hold29/X _14185_/Q _07506_/S vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__mux2_1
X_08484_ _08484_/A _08713_/A vssd1 vssd1 vccd1 vccd1 _08543_/A sky130_fd_sc_hd__or2_1
XFILLER_51_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07435_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07435_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_io_wbs_clk clkbuf_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_io_wbs_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07366_ _14215_/Q _14217_/Q _07387_/S vssd1 vssd1 vccd1 vccd1 _07366_/X sky130_fd_sc_hd__mux2_1
X_09105_ _09102_/X _09103_/Y _09071_/X _09023_/B vssd1 vssd1 vccd1 vccd1 _09106_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_56_io_wbs_clk clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14440_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07297_ _07519_/A vssd1 vssd1 vccd1 vccd1 _14192_/D sky130_fd_sc_hd__clkbuf_2
X_09036_ _08964_/Y _08965_/X _09034_/X _09035_/Y vssd1 vssd1 vccd1 vccd1 _10631_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_50_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07222__A0 _14087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09938_ _09938_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__xnor2_1
XFILLER_77_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09869_ _09869_/A _09869_/B vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__xor2_4
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11900_ _11902_/B vssd1 vssd1 vccd1 vccd1 _11900_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13525__A _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12880_ _14140_/Q _12872_/X _12878_/X _12879_/X vssd1 vssd1 vccd1 vccd1 _14140_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _14000_/Q _11797_/A _11830_/X _14119_/Q vssd1 vssd1 vccd1 vccd1 _11831_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ input59/X _11767_/B _11766_/B input60/X vssd1 vssd1 vccd1 vccd1 _12426_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12821__A2 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _12664_/X _14397_/Q _13511_/S vssd1 vssd1 vccd1 vccd1 _13502_/B sky130_fd_sc_hd__mux2_1
X_10713_ _10713_/A vssd1 vssd1 vccd1 vccd1 _10765_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _13770_/Q _11719_/B vssd1 vssd1 vccd1 vccd1 _11730_/B sky130_fd_sc_hd__or2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input92_A io_wbs_datwr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ _13444_/A _13432_/B vssd1 vssd1 vccd1 vccd1 _13433_/A sky130_fd_sc_hd__and2_1
XFILLER_13_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10644_ _10644_/A _10644_/B _10644_/C vssd1 vssd1 vccd1 vccd1 _10644_/X sky130_fd_sc_hd__and3_1
XFILLER_107_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _13375_/A _13363_/B vssd1 vssd1 vccd1 vccd1 _13364_/A sky130_fd_sc_hd__and2_1
X_10575_ _09664_/X _10574_/X _09655_/B vssd1 vssd1 vccd1 vccd1 _10576_/C sky130_fd_sc_hd__a21o_1
XFILLER_10_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ _12316_/A vssd1 vssd1 vccd1 vccd1 _12314_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13294_ _13315_/A vssd1 vssd1 vccd1 vccd1 _13294_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output179_A _14169_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12245_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07213__A0 _14274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12176_ _13202_/A _13203_/B vssd1 vssd1 vccd1 vccd1 _13359_/A sky130_fd_sc_hd__or2_4
XFILLER_110_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07764__A1 _14149_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _11127_/A _11127_/B _11127_/C vssd1 vssd1 vccd1 vccd1 _11127_/X sky130_fd_sc_hd__and3_1
XFILLER_7_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11058_ _11058_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11059_/B sky130_fd_sc_hd__or2_1
XANTENNA__09913__A _10271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10009_ _10009_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _10048_/B sky130_fd_sc_hd__xnor2_2
XFILLER_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07433__A _07460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_17_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14369__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07220_ _07220_/A vssd1 vssd1 vccd1 vccd1 _14272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07151_ _07240_/A vssd1 vssd1 vccd1 vccd1 _07259_/S sky130_fd_sc_hd__buf_2
XFILLER_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07082_ _07051_/X _07081_/X _14363_/Q vssd1 vssd1 vccd1 vccd1 _07083_/S sky130_fd_sc_hd__o21a_1
XFILLER_105_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07984_ _08012_/A _08573_/B _09241_/D _09234_/B vssd1 vssd1 vccd1 vccd1 _07985_/B
+ sky130_fd_sc_hd__and4_1
X_09723_ _09723_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _09724_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09823__A _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06935_ _14430_/Q _06942_/B _14462_/Q vssd1 vssd1 vccd1 vccd1 _06935_/X sky130_fd_sc_hd__and3b_1
XFILLER_80_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12500__A1 _10547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12500__B2 _14055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09654_ _09663_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _10596_/A sky130_fd_sc_hd__xnor2_1
XFILLER_103_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06866_ _14399_/Q _13778_/Q vssd1 vssd1 vccd1 vccd1 _06866_/X sky130_fd_sc_hd__xor2_1
X_08605_ _09053_/B _08982_/B _08983_/C _08978_/A vssd1 vssd1 vccd1 vccd1 _08605_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07343__A _14103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09585_ _09629_/A _09585_/B vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__xor2_1
XFILLER_103_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08536_ _08537_/A _08566_/B _08537_/C vssd1 vssd1 vccd1 vccd1 _08538_/A sky130_fd_sc_hd__a21oi_1
XFILLER_36_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08467_ _08828_/A vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07418_ _14090_/Q _07404_/X _07406_/X _13890_/Q _07417_/X vssd1 vssd1 vccd1 vccd1
+ _07418_/X sky130_fd_sc_hd__a221o_1
XANTENNA__13213__C1 _13053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08398_ _09690_/A _08403_/B vssd1 vssd1 vccd1 vccd1 _09729_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07349_ _07376_/A vssd1 vssd1 vccd1 vccd1 _07349_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10360_ _10360_/A _10360_/B _10360_/C vssd1 vssd1 vccd1 vccd1 _10361_/B sky130_fd_sc_hd__nor3_1
XFILLER_3_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09019_ _09098_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__xnor2_2
X_10291_ _09984_/A _10289_/Y _10290_/Y vssd1 vssd1 vccd1 vccd1 _10292_/B sky130_fd_sc_hd__o21a_1
XFILLER_88_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08621__B _08783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12030_ _12044_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12031_/A sky130_fd_sc_hd__and2_1
XFILLER_88_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08943__B1 _10171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13981_ _13982_/CLK _13981_/D _12408_/Y vssd1 vssd1 vccd1 vccd1 _13981_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12932_ _12932_/A _12940_/B vssd1 vssd1 vccd1 vccd1 _12932_/X sky130_fd_sc_hd__or2_1
XFILLER_19_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08349__A _14023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _14134_/Q _12857_/X _12862_/X _12817_/X vssd1 vssd1 vccd1 vccd1 _14134_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _14237_/Q _13037_/A _11800_/X _14113_/Q vssd1 vssd1 vccd1 vccd1 _11814_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _14155_/Q _12783_/X _12774_/A _14131_/Q vssd1 vssd1 vccd1 vccd1 _12794_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11153__S1 _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11745_ hold12/X vssd1 vssd1 vccd1 vccd1 _11745_/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_clkbuf_leaf_8_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14464_ _14464_/CLK _14464_/D vssd1 vssd1 vccd1 vccd1 _14464_/Q sky130_fd_sc_hd__dfxtp_1
X_11676_ _11659_/B _11679_/B _11675_/X _13779_/Q _11680_/D vssd1 vssd1 vccd1 vccd1
+ _13779_/D sky130_fd_sc_hd__o221a_1
XANTENNA__12558__A1 _09762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11222__B _11294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13415_ _13415_/A vssd1 vssd1 vccd1 vccd1 _14371_/D sky130_fd_sc_hd__clkbuf_1
X_10627_ _10627_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10627_/X sky130_fd_sc_hd__xor2_1
XFILLER_70_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14395_ _14440_/CLK _14395_/D vssd1 vssd1 vccd1 vccd1 _14395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13346_ _14432_/Q _13327_/X _13345_/X _13341_/X vssd1 vssd1 vccd1 vccd1 _13346_/X
+ sky130_fd_sc_hd__a211o_1
X_10558_ _10566_/A _10566_/B vssd1 vssd1 vccd1 vccd1 _10558_/X sky130_fd_sc_hd__or2_1
XFILLER_6_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ _14416_/Q _13199_/X _13275_/X _13276_/X vssd1 vssd1 vccd1 vccd1 _13277_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_29_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10489_ _10489_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10491_/C sky130_fd_sc_hd__xnor2_1
XFILLER_97_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12228_ _12209_/X _12229_/S _12227_/Y vssd1 vssd1 vccd1 vccd1 _13838_/D sky130_fd_sc_hd__o21a_1
XFILLER_97_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12159_ input91/X vssd1 vssd1 vccd1 vccd1 _12911_/A sky130_fd_sc_hd__buf_6
XFILLER_29_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13286__A2 _13236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _09074_/B _09286_/X _09369_/X vssd1 vssd1 vccd1 vccd1 _09371_/B sky130_fd_sc_hd__a21bo_1
XFILLER_91_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12797__A1 _14156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08321_ _08322_/B _08322_/C _08322_/A vssd1 vssd1 vccd1 vccd1 _08380_/A sky130_fd_sc_hd__a21o_2
XANTENNA__12797__B2 _14132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__A2 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08252_ _09999_/A _08252_/B _09088_/A vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__and3_1
XFILLER_21_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07203_ _07203_/A vssd1 vssd1 vccd1 vccd1 _07258_/S sky130_fd_sc_hd__buf_2
X_08183_ _09134_/A vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14198_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07134_ _14423_/Q _07134_/B _14455_/Q vssd1 vssd1 vccd1 vccd1 _07134_/X sky130_fd_sc_hd__and3b_1
XFILLER_106_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07065_ _14260_/Q _07046_/X _07064_/X _14356_/Q vssd1 vssd1 vccd1 vccd1 _07065_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07338__A _14227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07967_ _08004_/B _07968_/B _07969_/B vssd1 vssd1 vccd1 vccd1 _08024_/B sky130_fd_sc_hd__or3_1
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06896__B _07085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09706_ _09672_/X _09674_/X _09704_/X _09705_/Y vssd1 vssd1 vccd1 vccd1 _09706_/Y
+ sky130_fd_sc_hd__a211oi_2
X_06918_ _14432_/Q _06942_/B _14464_/Q vssd1 vssd1 vccd1 vccd1 _06918_/X sky130_fd_sc_hd__and3b_1
XFILLER_68_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07898_ _07897_/X _13976_/Q _07912_/S vssd1 vssd1 vccd1 vccd1 _07899_/A sky130_fd_sc_hd__mux2_1
XFILLER_83_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09637_ _09634_/Y _09635_/Y _09638_/A _09636_/Y vssd1 vssd1 vccd1 vccd1 _09638_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ _09565_/X _09566_/Y _09540_/A _09540_/Y vssd1 vssd1 vccd1 vccd1 _09586_/C
+ sky130_fd_sc_hd__o211ai_2
X_08519_ _08980_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08530_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12419__A _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ _09499_/A _09499_/B vssd1 vssd1 vccd1 vccd1 _09540_/B sky130_fd_sc_hd__xor2_1
XFILLER_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11530_ _11525_/A _11529_/Y _11464_/X vssd1 vssd1 vccd1 vccd1 _11530_/X sky130_fd_sc_hd__a21o_1
XFILLER_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11461_ _11534_/S vssd1 vssd1 vccd1 vccd1 _11461_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12853__S _12853_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09405__A1 _09641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13200_ _13206_/A _13200_/B vssd1 vssd1 vccd1 vccd1 _13637_/A sky130_fd_sc_hd__and2_2
X_10412_ _10412_/A _10412_/B vssd1 vssd1 vccd1 vccd1 _10418_/A sky130_fd_sc_hd__nand2_1
X_14180_ _14256_/CLK _14180_/D _12966_/Y vssd1 vssd1 vccd1 vccd1 _14180_/Q sky130_fd_sc_hd__dfrtp_1
X_11392_ _11392_/A vssd1 vssd1 vccd1 vccd1 _11392_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08632__A _08632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13131_ _13134_/A vssd1 vssd1 vccd1 vccd1 _13131_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10343_ _10314_/A _10314_/B _10342_/Y vssd1 vssd1 vccd1 vccd1 _10345_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12154__A _12906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A io_wbs_adr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13062_ _13062_/A _13079_/B vssd1 vssd1 vccd1 vccd1 _13076_/S sky130_fd_sc_hd__or2_4
X_10274_ _10274_/A _10274_/B _10272_/X vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__or3b_1
XFILLER_3_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12013_ _12013_/A vssd1 vssd1 vccd1 vccd1 _13786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13964_ _14031_/CLK _13964_/D _12388_/Y vssd1 vssd1 vccd1 vccd1 _13964_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12915_ _12928_/A vssd1 vssd1 vccd1 vccd1 _12915_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13895_ _13897_/CLK _13895_/D _12302_/Y vssd1 vssd1 vccd1 vccd1 _13895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12846_ _12645_/X _14130_/Q _12846_/S vssd1 vssd1 vccd1 vccd1 _12847_/B sky130_fd_sc_hd__mux2_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _14134_/Q _12776_/X _12760_/X vssd1 vssd1 vccd1 vccd1 _12777_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07104__C1 _14360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _13768_/Q _11714_/X _11716_/X _11727_/X vssd1 vssd1 vccd1 vccd1 _13768_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13728__A0 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _14449_/CLK _14447_/D vssd1 vssd1 vccd1 vccd1 _14447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11659_ _11659_/A _11659_/B vssd1 vssd1 vccd1 vccd1 _11669_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14378_ _14467_/CLK _14378_/D vssd1 vssd1 vccd1 vccd1 _14378_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08542__A _08571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ _14380_/Q _13328_/X _13315_/X _14460_/Q vssd1 vssd1 vccd1 vccd1 _13329_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09076__C _09076_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08870_ _08897_/A _08897_/B vssd1 vssd1 vccd1 vccd1 _08872_/B sky130_fd_sc_hd__and2_1
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07821_ _14032_/Q _13978_/Q vssd1 vssd1 vccd1 vccd1 _07848_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09092__B _09153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07752_ _07674_/Y _07723_/X _07724_/X vssd1 vssd1 vccd1 vccd1 _07752_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_38_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07683_ _14134_/Q vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__inv_2
XFILLER_93_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09422_ _09114_/Y _09115_/X _09032_/X _09040_/Y vssd1 vssd1 vccd1 vccd1 _10632_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_52_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07621__A _14132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09353_ _09313_/B _09313_/C _09313_/A vssd1 vssd1 vccd1 vccd1 _09354_/C sky130_fd_sc_hd__a21bo_1
X_08304_ _14023_/Q vssd1 vssd1 vccd1 vccd1 _09424_/A sky130_fd_sc_hd__clkbuf_2
X_09284_ _09284_/A _09284_/B _09284_/C vssd1 vssd1 vccd1 vccd1 _09291_/A sky130_fd_sc_hd__nand3_1
XFILLER_100_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ _08274_/A _08234_/B _08234_/C vssd1 vssd1 vccd1 vccd1 _08235_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08166_ _08167_/B _08167_/C _08243_/A vssd1 vssd1 vccd1 vccd1 _08168_/A sky130_fd_sc_hd__a21oi_1
XFILLER_118_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07117_ _14467_/Q _14291_/Q vssd1 vssd1 vccd1 vccd1 _07117_/Y sky130_fd_sc_hd__nand2_1
X_08097_ _08789_/A _08097_/B vssd1 vssd1 vccd1 vccd1 _09459_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08071__B1 _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07048_ _07087_/A vssd1 vssd1 vccd1 vccd1 _07048_/X sky130_fd_sc_hd__buf_2
XFILLER_47_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12702__A _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06909__C1 _14358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__A1 _08571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08999_ _08622_/A _08893_/A _08625_/B _08623_/X vssd1 vssd1 vccd1 vccd1 _09005_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06924__A2 _06873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10961_ _10722_/B _10944_/X _10960_/X _10729_/A vssd1 vssd1 vccd1 vccd1 _10961_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11130__B1 _10851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12700_ _12700_/A vssd1 vssd1 vccd1 vccd1 _14059_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13533__A _13539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13680_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13695_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10892_ _13931_/Q _10891_/X _10897_/S vssd1 vssd1 vccd1 vccd1 _10893_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12631_ _12635_/A _12631_/B vssd1 vssd1 vccd1 vccd1 _12632_/A sky130_fd_sc_hd__and2_1
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12630__A0 _12515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12562_ _12561_/X _09762_/A _12562_/S vssd1 vssd1 vccd1 vccd1 _12563_/B sky130_fd_sc_hd__mux2_1
XFILLER_54_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ _14411_/CLK _14301_/D _13168_/Y vssd1 vssd1 vccd1 vccd1 _14301_/Q sky130_fd_sc_hd__dfrtp_4
X_11513_ _11513_/A vssd1 vssd1 vccd1 vccd1 _11513_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12493_ _09762_/B _12486_/X _12476_/X _14053_/Q vssd1 vssd1 vccd1 vccd1 _12493_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14232_ _14441_/CLK _14232_/D vssd1 vssd1 vccd1 vccd1 _14232_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11444_ _11302_/A _11082_/A _11446_/S vssd1 vssd1 vccd1 vccd1 _11466_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14163_ _14163_/CLK _14163_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_2
X_11375_ _13853_/Q _11377_/B vssd1 vssd1 vccd1 vccd1 _11375_/X sky130_fd_sc_hd__or2_1
XFILLER_113_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13114_ _13114_/A vssd1 vssd1 vccd1 vccd1 _14258_/D sky130_fd_sc_hd__clkinv_2
XFILLER_113_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ _10326_/A _10373_/B vssd1 vssd1 vccd1 vccd1 _10598_/C sky130_fd_sc_hd__xor2_1
X_14094_ _14102_/CLK _14094_/D _12743_/Y vssd1 vssd1 vccd1 vccd1 _14094_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_output161_A _14316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ hold23/A _13036_/S _13042_/Y hold26/A _13032_/A vssd1 vssd1 vccd1 vccd1 _13045_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10257_ _10383_/A _10119_/B _10118_/B _10118_/A vssd1 vssd1 vccd1 vccd1 _10259_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12612__A _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09193__A _09402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ _10188_/A _10188_/B vssd1 vssd1 vccd1 vccd1 _10190_/A sky130_fd_sc_hd__xor2_1
XFILLER_61_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13947_ _13947_/CLK _13947_/D _12366_/Y vssd1 vssd1 vccd1 vccd1 _13947_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11121__B1 _11100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ _14198_/CLK _13878_/D _12281_/Y vssd1 vssd1 vccd1 vccd1 _13878_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12829_ _12827_/X _14125_/Q _12853_/S vssd1 vssd1 vccd1 vccd1 _12830_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12059__A _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12621__A0 _12942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09093__A2 _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08020_ _08131_/A _08020_/B _08078_/B vssd1 vssd1 vccd1 vccd1 _08078_/C sky130_fd_sc_hd__nor3_1
XANTENNA__09368__A _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08272__A _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ _10271_/A _10045_/A vssd1 vssd1 vccd1 vccd1 _09973_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08922_ _08953_/A _08953_/B vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08356__A1 _09153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__B2 _08623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08853_ _08850_/X _08883_/A _08840_/X _08811_/Y vssd1 vssd1 vccd1 vccd1 _08858_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_112_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07804_ _10648_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _10727_/B sky130_fd_sc_hd__nand2_1
X_08784_ _08842_/A _08937_/C _10156_/A _08716_/A vssd1 vssd1 vccd1 vccd1 _08803_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_38_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ _14069_/Q _07733_/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07736_/A sky130_fd_sc_hd__mux2_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07666_ _07666_/A _07642_/Y vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__or2b_1
XFILLER_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09405_ _09641_/A _09404_/C _09404_/B vssd1 vssd1 vccd1 vccd1 _09405_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07597_ _07597_/A vssd1 vssd1 vccd1 vccd1 _14085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09336_ _09336_/A _09408_/B vssd1 vssd1 vccd1 vccd1 _09345_/B sky130_fd_sc_hd__xor2_1
XFILLER_90_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10623__C1 _09788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _09267_/A _09267_/B vssd1 vssd1 vccd1 vccd1 _10621_/A sky130_fd_sc_hd__nor2_4
X_08218_ _08218_/A _08218_/B vssd1 vssd1 vccd1 vccd1 _08219_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08182__A _14009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09198_ _09198_/A _09198_/B _09198_/C vssd1 vssd1 vccd1 vccd1 _09198_/Y sky130_fd_sc_hd__nand3_1
XFILLER_14_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08149_ _09999_/A vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__buf_4
XFILLER_49_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11160_ _10771_/Y _11159_/X _11145_/X _10744_/A vssd1 vssd1 vccd1 vccd1 _11160_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10111_ _10111_/A _10111_/B vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13528__A _13634_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11091_ _11142_/B _10701_/X _11090_/Y _10826_/X vssd1 vssd1 vccd1 vccd1 _13927_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10042_ _10354_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _10042_/X sky130_fd_sc_hd__and2_1
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA__11048__A _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14102__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13801_ _14348_/CLK _13801_/D vssd1 vssd1 vccd1 vccd1 _13801_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11990__B _11990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input18_A dout1[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11103__B1 _11100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ input57/X input56/X _11993_/C input54/X vssd1 vssd1 vccd1 vccd1 _12952_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_90_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13732_ input85/X _14463_/Q _13738_/S vssd1 vssd1 vccd1 vccd1 _13733_/B sky130_fd_sc_hd__mux2_1
X_10944_ _13896_/Q _13897_/Q _10944_/S vssd1 vssd1 vccd1 vccd1 _10944_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08357__A _14020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07261__A _14165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13663_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13678_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10875_ _13976_/Q _10874_/Y _10875_/S vssd1 vssd1 vccd1 vccd1 _10875_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _12938_/A _14037_/Q _12621_/S vssd1 vssd1 vccd1 vccd1 _12615_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09075__A2 _09811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ _13607_/A _13594_/B vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__and2_1
XFILLER_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12545_ _12551_/A _12545_/B vssd1 vssd1 vccd1 vccd1 _12546_/A sky130_fd_sc_hd__and2_1
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09188__A _09188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12476_ _12476_/A vssd1 vssd1 vccd1 vccd1 _12476_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08092__A _14009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11230__B _11288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ _14215_/CLK _14215_/D _13009_/Y vssd1 vssd1 vccd1 vccd1 _14215_/Q sky130_fd_sc_hd__dfrtp_1
X_11427_ _11502_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10127__A _10127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14146_ _14149_/CLK _14146_/D vssd1 vssd1 vccd1 vccd1 _14146_/Q sky130_fd_sc_hd__dfxtp_2
X_11358_ _13857_/Q _11536_/B vssd1 vssd1 vccd1 vccd1 _11358_/X sky130_fd_sc_hd__and2_1
XFILLER_99_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _10338_/A _10338_/B vssd1 vssd1 vccd1 vccd1 _10310_/B sky130_fd_sc_hd__xor2_1
XFILLER_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14077_ _14283_/CLK _14077_/D _12721_/Y vssd1 vssd1 vccd1 vccd1 _14077_/Q sky130_fd_sc_hd__dfrtp_4
X_11289_ _11327_/A _11289_/B vssd1 vssd1 vccd1 vccd1 _11330_/A sky130_fd_sc_hd__or2_1
XFILLER_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12342__A _12348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _13028_/A vssd1 vssd1 vccd1 vccd1 _13028_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07520_ _14177_/Q _07520_/B vssd1 vssd1 vccd1 vccd1 _07520_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08267__A _08403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08510__A1 _08823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08510__B2 _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07451_ _07425_/X _07449_/X _07450_/X _07435_/X _14201_/Q vssd1 vssd1 vccd1 vccd1
+ _14201_/D sky130_fd_sc_hd__a32o_1
XFILLER_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07382_ _14096_/Q _07363_/X vssd1 vssd1 vccd1 vccd1 _07382_/X sky130_fd_sc_hd__or2b_1
X_09121_ _09191_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _09192_/B sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_46_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14354_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__12517__A _12517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09052_ _08468_/B _08132_/D _09793_/A _08925_/A vssd1 vssd1 vccd1 vccd1 _09054_/A
+ sky130_fd_sc_hd__a22oi_2
X_08003_ _08003_/A _08003_/B vssd1 vssd1 vccd1 vccd1 _08005_/A sky130_fd_sc_hd__xnor2_2
XFILLER_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08577__A1 _08716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09954_ _09954_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09954_/X sky130_fd_sc_hd__or2_1
XANTENNA__12252__A _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08905_ _08905_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _08906_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_24_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09885_ _09905_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09885_/X sky130_fd_sc_hd__and2_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08941_/A _08836_/B vssd1 vssd1 vccd1 vccd1 _08848_/A sky130_fd_sc_hd__nand2_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08767_ _08905_/A _08767_/B vssd1 vssd1 vccd1 vccd1 _08770_/A sky130_fd_sc_hd__nand2_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _14072_/Q _07717_/X _07730_/S vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__mux2_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _08791_/A _09457_/B _09866_/A _09199_/D vssd1 vssd1 vccd1 vccd1 _08745_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_26_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08177__A _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07649_ _14074_/Q _07656_/A vssd1 vssd1 vccd1 vccd1 _07706_/A sky130_fd_sc_hd__xnor2_2
XFILLER_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ _13948_/Q vssd1 vssd1 vccd1 vccd1 _10954_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08905__A _08905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09319_ _09319_/A _09319_/B vssd1 vssd1 vccd1 vccd1 _09321_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12061__A1 _13799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ _09663_/A _09663_/B _10597_/B vssd1 vssd1 vccd1 vccd1 _10592_/B sky130_fd_sc_hd__a21oi_1
X_12330_ _12348_/A vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__buf_2
XFILLER_103_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ _12385_/A vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_108_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14000_ _14396_/CLK _14000_/D vssd1 vssd1 vccd1 vccd1 _14000_/Q sky130_fd_sc_hd__dfxtp_1
X_11212_ _11216_/B _11217_/A _11216_/A vssd1 vssd1 vccd1 vccd1 _11213_/B sky130_fd_sc_hd__o21a_1
X_12192_ _12192_/A _13037_/B _13037_/C vssd1 vssd1 vccd1 vccd1 _12202_/C sky130_fd_sc_hd__and3_1
XFILLER_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11143_ _11143_/A vssd1 vssd1 vccd1 vccd1 _11143_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11074_ _11102_/B _11074_/B vssd1 vssd1 vccd1 vccd1 _11104_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10025_ _10110_/B _10110_/A vssd1 vssd1 vccd1 vccd1 _10025_/X sky130_fd_sc_hd__or2b_1
XFILLER_62_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11976_ _11976_/A vssd1 vssd1 vccd1 vccd1 _11976_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08087__A _14011_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13715_ input80/X _14458_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13716_/B sky130_fd_sc_hd__mux2_1
X_10927_ _10713_/A _10926_/X _10916_/X vssd1 vssd1 vccd1 vccd1 _10927_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13646_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10858_ _10858_/A _10858_/B _10858_/C vssd1 vssd1 vccd1 vccd1 _10858_/X sky130_fd_sc_hd__and3_1
XANTENNA__08815__A _09188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _13590_/A _13577_/B vssd1 vssd1 vccd1 vccd1 _13578_/A sky130_fd_sc_hd__and2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _10889_/B _10789_/B vssd1 vssd1 vccd1 vccd1 _10894_/C sky130_fd_sc_hd__or2_1
X_12528_ _12534_/A _12528_/B vssd1 vssd1 vccd1 vccd1 _12529_/A sky130_fd_sc_hd__and2_1
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12459_ _13993_/Q _12422_/X _12456_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _13993_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_67_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09756__B1 _09755_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14129_ _14152_/CLK _14129_/D vssd1 vssd1 vccd1 vccd1 _14129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06951_ _06934_/X _06950_/X _14380_/Q vssd1 vssd1 vccd1 vccd1 _06952_/S sky130_fd_sc_hd__o21a_1
XANTENNA__06990__B1 hold33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09670_ _09591_/A _09670_/B vssd1 vssd1 vccd1 vccd1 _09671_/B sky130_fd_sc_hd__and2b_1
XFILLER_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06882_ _14389_/Q _06865_/Y _13775_/Q _06881_/Y vssd1 vssd1 vccd1 vccd1 _06882_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_39_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08621_ _08621_/A _08783_/A vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08552_ _08716_/B _08899_/A vssd1 vssd1 vccd1 vccd1 _08559_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07503_ _07503_/A vssd1 vssd1 vccd1 vccd1 _14186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08483_ _08484_/A _08479_/Y _09491_/A _08863_/D vssd1 vssd1 vccd1 vccd1 _08713_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_51_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07434_ _14087_/Q _07432_/X _07433_/X _13887_/Q _07417_/X vssd1 vssd1 vccd1 vccd1
+ _07434_/X sky130_fd_sc_hd__a221o_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07365_ _07482_/S vssd1 vssd1 vccd1 vccd1 _07387_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__12247__A _12251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09104_ _09071_/X _09023_/B _09102_/X _09103_/Y vssd1 vssd1 vccd1 vccd1 _09106_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_109_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07296_ _07296_/A vssd1 vssd1 vccd1 vccd1 _14227_/D sky130_fd_sc_hd__clkbuf_1
X_09035_ _09032_/X _09033_/Y _08688_/A _08966_/X vssd1 vssd1 vccd1 vccd1 _09035_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_108_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08460__A _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09937_ _09937_/A vssd1 vssd1 vccd1 vccd1 _10003_/A sky130_fd_sc_hd__inv_2
XFILLER_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09868_ _10126_/B _10083_/A vssd1 vssd1 vccd1 vccd1 _09872_/A sky130_fd_sc_hd__nor2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08819_ _08798_/A _08797_/A _08797_/B vssd1 vssd1 vccd1 vccd1 _08837_/B sky130_fd_sc_hd__o21ba_1
XFILLER_100_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09799_ _09799_/A vssd1 vssd1 vccd1 vccd1 _10280_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _12768_/A vssd1 vssd1 vccd1 vccd1 _11830_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12806__B1 _12804_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ input61/X _11774_/B _11774_/C vssd1 vssd1 vccd1 vccd1 _11766_/B sky130_fd_sc_hd__nor3_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13500_/A vssd1 vssd1 vccd1 vccd1 _14396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _11164_/S vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13541__A _13592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _13769_/Q _11692_/B vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__or2_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ input78/X _14376_/Q _13443_/S vssd1 vssd1 vccd1 vccd1 _13432_/B sky130_fd_sc_hd__mux2_1
X_10643_ _10631_/A _09037_/X _10642_/X vssd1 vssd1 vccd1 vccd1 _10644_/C sky130_fd_sc_hd__o21ai_4
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12157__A _12909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11061__A _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input85_A io_wbs_datwr[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13362_ _12827_/X _14356_/Q _13374_/S vssd1 vssd1 vccd1 vccd1 _13363_/B sky130_fd_sc_hd__mux2_1
X_10574_ _10596_/B _10596_/C _10592_/A _10596_/A vssd1 vssd1 vccd1 vccd1 _10574_/X
+ sky130_fd_sc_hd__a211o_1
X_12313_ _12316_/A vssd1 vssd1 vccd1 vccd1 _12313_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11996__A _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07461__A1 _14082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13293_ _14339_/Q _13289_/X _13292_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _14339_/D
+ sky130_fd_sc_hd__o211a_1
X_12244_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12244_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14440__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07213__A1 _07212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ _12933_/A vssd1 vssd1 vccd1 vccd1 _13343_/A sky130_fd_sc_hd__buf_4
XFILLER_64_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11126_ _11054_/A _11110_/X _11124_/X _11125_/Y vssd1 vssd1 vccd1 vccd1 _13915_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11057_ _11122_/B _11125_/B _11122_/A vssd1 vssd1 vccd1 vccd1 _11120_/C sky130_fd_sc_hd__o21ai_1
XFILLER_27_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10008_ _10007_/Y _09848_/X _09847_/X vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__a21oi_1
XFILLER_114_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11959_ _11959_/A vssd1 vssd1 vccd1 vccd1 _11959_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08545__A _14018_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13629_ _13644_/A _13629_/B vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__and2_1
XANTENNA__12025__B2 _13830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12067__A _12536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07150_ _07150_/A _14259_/D vssd1 vssd1 vccd1 vccd1 _07240_/A sky130_fd_sc_hd__and2_2
XFILLER_69_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07081_ _14411_/Q _07098_/B _14443_/Q vssd1 vssd1 vccd1 vccd1 _07081_/X sky130_fd_sc_hd__and3b_1
XFILLER_69_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07983_ _13872_/Q vssd1 vssd1 vccd1 vccd1 _09234_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10034__B _10090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09722_ _09723_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _09724_/A sky130_fd_sc_hd__or2_2
XANTENNA__11839__A1 _14338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06934_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06934_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08704__A1 _09241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08704__B2 _09241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _09411_/B _09411_/C _09411_/A vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__a21bo_4
XFILLER_83_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06865_ _13776_/Q vssd1 vssd1 vccd1 vccd1 _06865_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08604_ _09053_/A _09053_/B _08983_/C vssd1 vssd1 vccd1 vccd1 _08604_/X sky130_fd_sc_hd__and3_1
XFILLER_83_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09584_ _09584_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09585_/B sky130_fd_sc_hd__xnor2_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08535_ _08470_/A _08469_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08537_/C sky130_fd_sc_hd__o21ba_1
XFILLER_24_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13361__A _13467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08466_ _14011_/Q vssd1 vssd1 vccd1 vccd1 _08828_/A sky130_fd_sc_hd__buf_2
XFILLER_51_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07417_ _07471_/A vssd1 vssd1 vccd1 vccd1 _07417_/X sky130_fd_sc_hd__clkbuf_2
X_08397_ _09673_/A _08402_/B vssd1 vssd1 vccd1 vccd1 _08403_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07348_ _07348_/A vssd1 vssd1 vccd1 vccd1 _07348_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07279_ _07280_/A _07307_/B _07307_/C vssd1 vssd1 vccd1 vccd1 _07312_/B sky130_fd_sc_hd__nor3_1
X_09018_ _09088_/A _10092_/A _09017_/X vssd1 vssd1 vccd1 vccd1 _09098_/B sky130_fd_sc_hd__o21a_1
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10290_ _10290_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _10290_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08190__A _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10225__A _10279_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08943__A1 _08937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__B2 _08946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13536__A _13539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13980_ _14102_/CLK _13980_/D _12407_/Y vssd1 vssd1 vccd1 vccd1 _13980_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12931_ _14159_/Q _12928_/X _12930_/X _12920_/X vssd1 vssd1 vccd1 vccd1 _14159_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11056__A _11056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12862_ _12906_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__or2_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ _14328_/Q _11808_/X _11811_/X _11812_/X vssd1 vssd1 vccd1 vccd1 _11813_/X
+ sky130_fd_sc_hd__a211o_4
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12793_ _14113_/Q _12782_/X _12790_/X _12792_/X _12216_/X vssd1 vssd1 vccd1 vccd1
+ _14113_/D sky130_fd_sc_hd__o221a_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09656__C1 _10632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11740_/B _11714_/A _11716_/A _11743_/X vssd1 vssd1 vccd1 vccd1 _13763_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14463_ _14464_/CLK _14463_/D vssd1 vssd1 vccd1 vccd1 _14463_/Q sky130_fd_sc_hd__dfxtp_1
X_11675_ _11675_/A _11682_/C vssd1 vssd1 vccd1 vccd1 _11675_/X sky130_fd_sc_hd__and2_1
XANTENNA__12007__B2 _13825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13414_ _13426_/A _13414_/B vssd1 vssd1 vccd1 vccd1 _13415_/A sky130_fd_sc_hd__and2_1
X_10626_ _10626_/A _10626_/B vssd1 vssd1 vccd1 vccd1 _10626_/Y sky130_fd_sc_hd__nor2_1
X_14394_ _14440_/CLK _14394_/D vssd1 vssd1 vccd1 vccd1 _14394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13345_ _14384_/Q _13328_/X _13336_/X _14464_/Q vssd1 vssd1 vccd1 vccd1 _13345_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07434__A1 _14087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557_ _10557_/A _10557_/B _10557_/C vssd1 vssd1 vccd1 vccd1 _10566_/A sky130_fd_sc_hd__and3_1
XANTENNA__13830__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13276_ _14368_/Q _13236_/X _13210_/X vssd1 vssd1 vccd1 vccd1 _13276_/X sky130_fd_sc_hd__a21o_1
X_10488_ _09766_/A _09969_/A _09969_/B _09998_/A vssd1 vssd1 vccd1 vccd1 _10489_/B
+ sky130_fd_sc_hd__a22o_1
X_12227_ _07146_/B _12229_/S _11935_/A vssd1 vssd1 vccd1 vccd1 _12227_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07198__A0 _14278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12158_ _13825_/Q _12146_/X _12157_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _13825_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13980__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _11007_/B _10701_/X _11107_/X _11108_/Y vssd1 vssd1 vccd1 vccd1 _13921_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13446__A _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12089_ _13062_/A vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__buf_4
XFILLER_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07444__A _07471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13691__A0 _12688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12494__A1 _14037_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13443__A0 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08320_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__xnor2_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08251_ _08251_/A _08312_/A vssd1 vssd1 vccd1 vccd1 _09088_/A sky130_fd_sc_hd__nand2_4
XFILLER_21_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07202_ _07202_/A vssd1 vssd1 vccd1 vccd1 _14277_/D sky130_fd_sc_hd__clkbuf_1
X_08182_ _14009_/Q vssd1 vssd1 vccd1 vccd1 _09134_/A sky130_fd_sc_hd__buf_2
XFILLER_119_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07133_ _14279_/Q _06968_/A _07132_/X _14375_/Q vssd1 vssd1 vccd1 vccd1 _07133_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09818__B _09818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07064_ _14404_/Q _07063_/Y _07048_/X vssd1 vssd1 vccd1 vccd1 _07064_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07189__A0 _14281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09834__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12260__A _13153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07966_ _07966_/A _08315_/A vssd1 vssd1 vccd1 vccd1 _07969_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09705_ _09702_/X _09703_/Y _09692_/A _09692_/Y vssd1 vssd1 vccd1 vccd1 _09705_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_114_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06917_ _14288_/Q _06873_/X _06916_/X _14384_/Q vssd1 vssd1 vccd1 vccd1 _06917_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07897_ _07897_/A _07897_/B vssd1 vssd1 vccd1 vccd1 _07897_/X sky130_fd_sc_hd__xor2_1
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09350__A1 _08791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _09527_/X _09632_/Y _09631_/A _09631_/Y vssd1 vssd1 vccd1 vccd1 _09636_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__09350__B2 _08791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13434__A0 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ _09540_/A _09540_/Y _09565_/X _09566_/Y vssd1 vssd1 vccd1 vccd1 _09586_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_71_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08518_ _08517_/A _08517_/C _08517_/B vssd1 vssd1 vccd1 vccd1 _08531_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09498_ _09496_/X _09498_/B vssd1 vssd1 vccd1 vccd1 _09499_/B sky130_fd_sc_hd__and2b_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08449_ _09233_/A _08449_/B _08449_/C _09011_/B vssd1 vssd1 vccd1 vccd1 _08503_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ _11513_/A vssd1 vssd1 vccd1 vccd1 _11460_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ _10411_/A _10459_/B vssd1 vssd1 vccd1 vccd1 _10412_/B sky130_fd_sc_hd__or2b_1
X_11391_ _13883_/Q _11379_/X _11383_/X _11390_/X vssd1 vssd1 vccd1 vccd1 _13883_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08632__B _09001_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13130_ _13134_/A vssd1 vssd1 vccd1 vccd1 _13130_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10342_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10342_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _12904_/A _12210_/X _13079_/B _13060_/X _12008_/A vssd1 vssd1 vccd1 vccd1
+ _14240_/D sky130_fd_sc_hd__o311a_1
X_10273_ _10274_/A _10274_/B _10272_/X vssd1 vssd1 vccd1 vccd1 _10273_/X sky130_fd_sc_hd__o21ba_1
X_12012_ _12026_/A _12012_/B vssd1 vssd1 vccd1 vccd1 _12013_/A sky130_fd_sc_hd__and2_1
XANTENNA_input48_A io_wbs_adr[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12170__A _12919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14359__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13963_ _13963_/CLK _13963_/D _12387_/Y vssd1 vssd1 vccd1 vccd1 _13963_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12914_ _14153_/Q _12901_/X _12913_/X _12907_/X vssd1 vssd1 vccd1 vccd1 _14153_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13894_ _13897_/CLK _13894_/D _12301_/Y vssd1 vssd1 vccd1 vccd1 _13894_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12845_ _12845_/A vssd1 vssd1 vccd1 vccd1 _14129_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12228__A1 _12209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13425__A0 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08807__B _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__A _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__A2 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12776_/A vssd1 vssd1 vccd1 vccd1 _12776_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11727_ _11692_/B _11726_/Y _11718_/X _13828_/Q vssd1 vssd1 vccd1 vccd1 _11727_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_30_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11658_ _13779_/Q _11675_/A vssd1 vssd1 vccd1 vccd1 _11659_/B sky130_fd_sc_hd__nand2_1
X_14446_ _14449_/CLK _14446_/D vssd1 vssd1 vccd1 vccd1 _14446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08823__A _08823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07407__A1 _14092_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10609_ _10032_/A _10032_/B _10608_/X vssd1 vssd1 vccd1 vccd1 _10610_/B sky130_fd_sc_hd__o21ai_1
X_14377_ _14457_/CLK _14377_/D vssd1 vssd1 vccd1 vccd1 _14377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11589_ _13856_/Q _11655_/B vssd1 vssd1 vccd1 vccd1 _11589_/X sky130_fd_sc_hd__and2_1
XANTENNA__08542__B _08783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13328_ _13328_/A vssd1 vssd1 vccd1 vccd1 _13328_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13259_ _14364_/Q _13208_/X _13257_/X _13258_/X vssd1 vssd1 vccd1 vccd1 _13259_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ _14033_/Q _13979_/Q vssd1 vssd1 vccd1 vccd1 _07885_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07591__A0 _14087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_29_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07751_ _14153_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07751_/X sky130_fd_sc_hd__and2_1
XANTENNA__13664__A0 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12467__A1 _14030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07682_ _07685_/B _07682_/B vssd1 vssd1 vccd1 vccd1 _07763_/A sky130_fd_sc_hd__nand2_1
XFILLER_53_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12188__A_N _12211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09421_ _10621_/A _10627_/B _09421_/C _10613_/C vssd1 vssd1 vccd1 vccd1 _09421_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13416__A0 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _09351_/A _09351_/C _09351_/B vssd1 vssd1 vccd1 vccd1 _09354_/B sky130_fd_sc_hd__o21ai_1
XFILLER_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08303_ _08002_/A _08684_/A _07966_/A _07963_/Y vssd1 vssd1 vccd1 vccd1 _08315_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_100_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09283_ _09202_/B _09202_/C _09202_/A vssd1 vssd1 vccd1 vccd1 _09284_/C sky130_fd_sc_hd__a21bo_1
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08234_ _08274_/A _08234_/B _08234_/C vssd1 vssd1 vccd1 vccd1 _08274_/B sky130_fd_sc_hd__nor3_2
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09829__A _10435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08733__A _08905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12927__C1 _12920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08165_ _08298_/A vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07116_ _07116_/A vssd1 vssd1 vccd1 vccd1 _14295_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07349__A _07376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08096_ _14012_/Q vssd1 vssd1 vccd1 vccd1 _08789_/A sky130_fd_sc_hd__clkbuf_2
X_07047_ _14447_/Q _14271_/Q vssd1 vssd1 vccd1 vccd1 _07047_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08374__A2 _08980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08998_ _08998_/A _08998_/B vssd1 vssd1 vccd1 vccd1 _09007_/A sky130_fd_sc_hd__nand2_1
XFILLER_75_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07949_ _08004_/A _07944_/Y _08135_/A _09793_/A vssd1 vssd1 vccd1 vccd1 _08004_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10960_ _13898_/Q _13899_/Q _10960_/S vssd1 vssd1 vccd1 vccd1 _10960_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11130__A1 _11119_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11130__B2 _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09619_ _09721_/B _09617_/Y _09575_/X _09622_/A vssd1 vssd1 vccd1 vccd1 _09666_/A
+ sky130_fd_sc_hd__a211oi_1
X_10891_ _10836_/S _10884_/C _10889_/X _10890_/X vssd1 vssd1 vccd1 vccd1 _10891_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12630_ _12515_/X _14041_/Q _12642_/S vssd1 vssd1 vccd1 vccd1 _12631_/B sky130_fd_sc_hd__mux2_1
XFILLER_93_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12561_ input71/X vssd1 vssd1 vccd1 vccd1 _12561_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_31_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ _11506_/A _11511_/Y _11472_/X vssd1 vssd1 vccd1 vccd1 _11512_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14300_ _14367_/CLK _14300_/D _13167_/Y vssd1 vssd1 vccd1 vccd1 _14300_/Q sky130_fd_sc_hd__dfrtp_4
X_12492_ _14001_/Q _12481_/X _12491_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _14001_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14231_ _14244_/CLK _14231_/D _13030_/Y vssd1 vssd1 vccd1 vccd1 _14231_/Q sky130_fd_sc_hd__dfrtp_2
X_11443_ _11471_/A _11471_/B vssd1 vssd1 vccd1 vccd1 _11466_/A sky130_fd_sc_hd__nand2_1
X_14162_ _14163_/CLK _14162_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_2
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11374_ _13890_/Q _11363_/X _11370_/X _11373_/X vssd1 vssd1 vccd1 vccd1 _13890_/D
+ sky130_fd_sc_hd__a22o_1
X_13113_ _14258_/Q _13113_/B _12185_/A vssd1 vssd1 vccd1 vccd1 _13114_/A sky130_fd_sc_hd__or3b_1
X_10325_ _10346_/A _09995_/B _09994_/A vssd1 vssd1 vccd1 vccd1 _10373_/B sky130_fd_sc_hd__a21o_1
X_14093_ _14102_/CLK _14093_/D _12742_/Y vssd1 vssd1 vccd1 vccd1 _14093_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14181__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13044_ _14233_/Q _13041_/X _13043_/X _13039_/X vssd1 vssd1 vccd1 vccd1 _14233_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ _10395_/A _10256_/B vssd1 vssd1 vccd1 vccd1 _10259_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13749__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output154_A _14310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10187_ _10151_/X _10169_/Y _10185_/Y _10186_/Y vssd1 vssd1 vccd1 vccd1 _10187_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12449__A1 _08891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09314__A1 _08867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13946_ _13946_/CLK _13946_/D _12365_/Y vssd1 vssd1 vccd1 vccd1 _13946_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11121__A1 _11119_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11121__B2 _11058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07722__A hold1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13877_ _14028_/CLK _13877_/D _12279_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_90_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11244__A _11244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ _12828_/A _12828_/B _12828_/C _13200_/B vssd1 vssd1 vccd1 vccd1 _12853_/S
+ sky130_fd_sc_hd__or4b_4
XFILLER_37_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12621__A1 _14039_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12768_/A _13037_/B _13037_/C vssd1 vssd1 vccd1 vccd1 _12809_/A sky130_fd_sc_hd__nand3_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_36_io_wbs_clk clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14304_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_72_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08553__A _14017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14429_ _14465_/CLK _14429_/D vssd1 vssd1 vccd1 vccd1 _14429_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09368__B _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09970_ _09970_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__xnor2_2
X_08921_ _08921_/A _08921_/B vssd1 vssd1 vccd1 vccd1 _08953_/B sky130_fd_sc_hd__or2_1
XFILLER_83_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09002__B1 _09091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08852_ _08858_/B vssd1 vssd1 vccd1 vccd1 _08852_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07803_ _11164_/S _10676_/A _10670_/B vssd1 vssd1 vccd1 vccd1 _07804_/B sky130_fd_sc_hd__and3_2
XFILLER_57_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08783_ _08783_/A vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__buf_2
XFILLER_84_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07734_ _07765_/S vssd1 vssd1 vccd1 vccd1 _07761_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_75_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14158_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07665_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07665_/Y sky130_fd_sc_hd__nand2_2
XFILLER_26_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09404_ _09641_/A _09404_/B _09404_/C vssd1 vssd1 vccd1 vccd1 _09404_/X sky130_fd_sc_hd__and3_2
XFILLER_77_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07596_ _14085_/Q input32/X _07604_/S vssd1 vssd1 vccd1 vccd1 _07597_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09335_ _09335_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09408_/B sky130_fd_sc_hd__xnor2_1
X_09266_ _09262_/X _09264_/Y _09187_/X _09190_/Y vssd1 vssd1 vccd1 vccd1 _09267_/B
+ sky130_fd_sc_hd__o211a_2
X_08217_ _08217_/A _08217_/B _08217_/C vssd1 vssd1 vccd1 vccd1 _08218_/B sky130_fd_sc_hd__nand3_1
X_09197_ _09629_/A _09341_/B vssd1 vssd1 vccd1 vccd1 _09274_/A sky130_fd_sc_hd__xor2_2
XFILLER_101_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08148_ _10000_/A vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08079_ _08167_/B _08079_/B vssd1 vssd1 vccd1 vccd1 _08163_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10110_ _10110_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10111_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07807__A _14007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11090_ _11090_/A _11090_/B vssd1 vssd1 vccd1 vccd1 _11090_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09544__A1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _10354_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _10073_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09544__B2 _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10233__A _10271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13800_ _14400_/CLK _13800_/D vssd1 vssd1 vccd1 vccd1 _13800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11992_ input99/X input53/X vssd1 vssd1 vccd1 vccd1 _11993_/C sky130_fd_sc_hd__nand2_1
XFILLER_99_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11103__B2 _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10943_ _10936_/B _10933_/X _13949_/Q vssd1 vssd1 vccd1 vccd1 _10943_/X sky130_fd_sc_hd__mux2_2
X_13731_ _13731_/A vssd1 vssd1 vccd1 vccd1 _13745_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13662_ _13662_/A vssd1 vssd1 vccd1 vccd1 _14442_/D sky130_fd_sc_hd__clkbuf_1
X_10874_ _10874_/A _10874_/B vssd1 vssd1 vccd1 vccd1 _10874_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12613_ _12613_/A vssd1 vssd1 vccd1 vccd1 _14036_/D sky130_fd_sc_hd__clkbuf_1
X_13593_ input76/X _14423_/Q _13593_/S vssd1 vssd1 vccd1 vccd1 _13594_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12544_ _12926_/A _08632_/A _12555_/S vssd1 vssd1 vccd1 vccd1 _12545_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09480__B1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08373__A _09824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09188__B _09188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12475_ _13997_/Q _12460_/X _12474_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _13997_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08092__B _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ _11426_/A vssd1 vssd1 vccd1 vccd1 _11502_/B sky130_fd_sc_hd__inv_2
X_14214_ _14217_/CLK _14214_/D _13008_/Y vssd1 vssd1 vccd1 vccd1 _14214_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14145_ _14149_/CLK _14145_/D vssd1 vssd1 vccd1 vccd1 _14145_/Q sky130_fd_sc_hd__dfxtp_2
X_11357_ _14057_/Q _13969_/Q vssd1 vssd1 vccd1 vccd1 _11536_/B sky130_fd_sc_hd__or2_2
XANTENNA__10842__S _10875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ _10284_/A _10284_/B _10307_/X vssd1 vssd1 vccd1 vccd1 _10338_/B sky130_fd_sc_hd__a21oi_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14076_ _14283_/CLK _14076_/D _12720_/Y vssd1 vssd1 vccd1 vccd1 _14076_/Q sky130_fd_sc_hd__dfrtp_4
X_11288_ _11288_/A _11288_/B vssd1 vssd1 vccd1 vccd1 _11289_/B sky130_fd_sc_hd__nor2_1
XFILLER_98_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _13028_/A vssd1 vssd1 vccd1 vccd1 _13027_/Y sky130_fd_sc_hd__inv_2
X_10239_ _10151_/X _10169_/Y _10187_/X vssd1 vssd1 vccd1 vccd1 _10239_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11878__C1 _11874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07546__A0 _14107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08548__A _08824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07452__A _07452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13929_ _13987_/CLK _13929_/D _12344_/Y vssd1 vssd1 vccd1 vccd1 _13929_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07450_ _14084_/Q _07432_/X _07433_/X _13884_/Q _07444_/X vssd1 vssd1 vccd1 vccd1
+ _07450_/X sky130_fd_sc_hd__a221o_1
XFILLER_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07381_ _14214_/Q _07373_/X _07375_/X _07380_/X vssd1 vssd1 vccd1 vccd1 _14214_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09120_ _09054_/A _09056_/B _09054_/B vssd1 vssd1 vccd1 vccd1 _09191_/B sky130_fd_sc_hd__o21ba_1
XFILLER_31_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10605__B1 _10597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09379__A _13870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11802__C1 _11801_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09051_ _09007_/A _09007_/C _09007_/B vssd1 vssd1 vccd1 vccd1 _09067_/A sky130_fd_sc_hd__a21bo_1
X_14476__188 vssd1 vssd1 vccd1 vccd1 _14476__188/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XANTENNA__10318__A _10393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08002_ _08002_/A _08132_/D vssd1 vssd1 vccd1 vccd1 _08003_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13629__A _13644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09953_ _09954_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__xnor2_1
XFILLER_106_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08904_ _08904_/A _08904_/B vssd1 vssd1 vccd1 vccd1 _08911_/A sky130_fd_sc_hd__xnor2_1
XFILLER_112_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09884_ _09884_/A _13860_/Q vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__or2_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12530__A0 _12917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09842__A _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08835_ _08837_/B _08844_/B vssd1 vssd1 vccd1 vccd1 _08839_/A sky130_fd_sc_hd__or2b_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10988__A _11092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08766_ _08764_/A _08764_/C _08805_/C vssd1 vssd1 vccd1 vccd1 _08771_/B sky130_fd_sc_hd__o21ai_1
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08458__A _09132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ _07716_/Y hold14/X _07723_/A vssd1 vssd1 vccd1 vccd1 _07717_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _09865_/A vssd1 vssd1 vccd1 vccd1 _09866_/A sky130_fd_sc_hd__buf_2
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07081__B _07098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07648_ _14073_/Q _07716_/A vssd1 vssd1 vccd1 vccd1 _07656_/A sky130_fd_sc_hd__and2_1
XFILLER_0_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07579_ _07579_/A vssd1 vssd1 vccd1 vccd1 _14093_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12597__A0 _12924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08905__B _10215_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09318_ _08208_/C _08091_/A _09317_/Y vssd1 vssd1 vccd1 vccd1 _09319_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12061__A2 _12059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10590_ _10596_/B _10596_/C _10596_/A vssd1 vssd1 vccd1 vccd1 _10597_/B sky130_fd_sc_hd__a21oi_1
XFILLER_103_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09249_ _09248_/A _09248_/C _09248_/B vssd1 vssd1 vccd1 vccd1 _09249_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12260_ _13153_/A vssd1 vssd1 vccd1 vccd1 _12385_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11211_ _11300_/A vssd1 vssd1 vccd1 vccd1 _11214_/A sky130_fd_sc_hd__clkinv_2
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13539__A _13539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ _13194_/C vssd1 vssd1 vccd1 vccd1 _13037_/C sky130_fd_sc_hd__clkbuf_2
X_11142_ _11142_/A _11142_/B vssd1 vssd1 vccd1 vccd1 _11143_/A sky130_fd_sc_hd__or2_2
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11073_ _11002_/B _11073_/B vssd1 vssd1 vccd1 vccd1 _11074_/B sky130_fd_sc_hd__and2b_1
XFILLER_95_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10024_ _10110_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10024_/X sky130_fd_sc_hd__and2b_1
XFILLER_27_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input30_A dout1[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11875__A2 _11872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13274__A _13637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__A _14017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11975_ _11976_/A vssd1 vssd1 vccd1 vccd1 _11975_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08087__B _08796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13714_ _13731_/A vssd1 vssd1 vccd1 vccd1 _13729_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10926_ _13907_/Q _13908_/Q _13909_/Q _13910_/Q _10944_/S _10946_/A vssd1 vssd1 vccd1
+ vccd1 _10926_/X sky130_fd_sc_hd__mux4_2
XFILLER_108_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13645_ _13645_/A vssd1 vssd1 vccd1 vccd1 _14437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10857_ _10857_/A vssd1 vssd1 vccd1 vccd1 _13938_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08815__B _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09199__A _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _12561_/X _14418_/Q _13576_/S vssd1 vssd1 vccd1 vccd1 _13577_/B sky130_fd_sc_hd__mux2_1
X_10788_ _13930_/Q _10788_/B vssd1 vssd1 vccd1 vccd1 _10789_/B sky130_fd_sc_hd__nor2_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12527_ _12913_/A _08896_/A _12537_/S vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__mux2_1
XFILLER_75_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12458_ _12817_/A vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__clkbuf_2
X_11409_ _13946_/Q _13945_/Q vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__nand2_2
X_12389_ _12391_/A vssd1 vssd1 vccd1 vccd1 _12389_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07447__A _14227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ _14152_/CLK _14128_/D vssd1 vssd1 vccd1 vccd1 _14128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06950_ _14428_/Q _06981_/B _14460_/Q vssd1 vssd1 vccd1 vccd1 _06950_/X sky130_fd_sc_hd__and3b_1
XFILLER_113_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14059_ _14164_/CLK _14059_/D vssd1 vssd1 vccd1 vccd1 _14059_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12512__A0 _12218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09084__D _09084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06881_ _14388_/Q vssd1 vssd1 vccd1 vccd1 _06881_/Y sky130_fd_sc_hd__inv_2
X_08620_ _08620_/A _08620_/B _08618_/X vssd1 vssd1 vccd1 vccd1 _08620_/X sky130_fd_sc_hd__or3b_1
XANTENNA__13184__A _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08278__A _09777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08551_ _09092_/C vssd1 vssd1 vccd1 vccd1 _08899_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07502_ hold18/X _14186_/Q _07506_/S vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08482_ _09905_/A vssd1 vssd1 vccd1 vccd1 _08863_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_74_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07433_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07433_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07364_ _14099_/Q _07363_/X vssd1 vssd1 vccd1 vccd1 _07364_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09103_ _09144_/B _09144_/C _09144_/A vssd1 vssd1 vccd1 vccd1 _09103_/Y sky130_fd_sc_hd__a21oi_2
X_07295_ _14244_/Q _07333_/S _07506_/S vssd1 vssd1 vccd1 vccd1 _07296_/A sky130_fd_sc_hd__mux2_1
X_09034_ _08688_/A _08966_/X _09032_/X _09033_/Y vssd1 vssd1 vccd1 vccd1 _09034_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13359__A _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09936_ _10394_/A _09939_/B _09935_/X vssd1 vssd1 vccd1 vccd1 _09937_/A sky130_fd_sc_hd__a21o_1
XFILLER_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09867_ _09887_/A _09887_/B _09866_/X vssd1 vssd1 vccd1 vccd1 _10083_/A sky130_fd_sc_hd__a21oi_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _08818_/A _08856_/A vssd1 vssd1 vccd1 vccd1 _08962_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14392__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10511__A _10597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09798_ _09800_/A _09799_/A vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__or2_1
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _09348_/B _09884_/A _09145_/D _08750_/A vssd1 vssd1 vccd1 vccd1 _08787_/C
+ sky130_fd_sc_hd__a22oi_2
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ input64/X input63/X input35/X input34/X vssd1 vssd1 vccd1 vccd1 _11774_/C
+ sky130_fd_sc_hd__or4_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07820__A _14033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _11244_/A _10727_/B vssd1 vssd1 vccd1 vccd1 _10716_/B sky130_fd_sc_hd__nand2_1
X_11691_ _13768_/Q _13767_/Q _11729_/B vssd1 vssd1 vccd1 vccd1 _11692_/B sky130_fd_sc_hd__or3_1
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12438__A _12485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _08780_/X _08963_/X _09038_/Y vssd1 vssd1 vccd1 vccd1 _10642_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13430_ _13447_/A vssd1 vssd1 vccd1 vccd1 _13443_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__13231__A1 _14439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13361_ _13467_/S vssd1 vssd1 vccd1 vccd1 _13374_/S sky130_fd_sc_hd__clkbuf_2
X_10573_ _10644_/B _09117_/Y _09421_/Y _10632_/A vssd1 vssd1 vccd1 vccd1 _10596_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12312_ _12316_/A vssd1 vssd1 vccd1 vccd1 _12312_/Y sky130_fd_sc_hd__inv_2
X_13292_ _14419_/Q _13284_/X _13290_/X _13291_/X vssd1 vssd1 vccd1 vccd1 _13292_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_108_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input78_A io_wbs_datwr[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08651__A _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12243_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12173__A _12922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07267__A _14165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ _13830_/Q _12095_/A _12173_/X _12161_/X vssd1 vssd1 vccd1 vccd1 _13830_/D
+ sky130_fd_sc_hd__o211a_1
X_11125_ _11125_/A _11125_/B vssd1 vssd1 vccd1 vccd1 _11125_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12901__A _12928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06972__A1 _14281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09482__A _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11056_ _11056_/A _11056_/B vssd1 vssd1 vccd1 vccd1 _11122_/A sky130_fd_sc_hd__xor2_1
XFILLER_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10007_ _10007_/A vssd1 vssd1 vccd1 vccd1 _10007_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11958_ _11959_/A vssd1 vssd1 vccd1 vccd1 _11958_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08826__A _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10909_ _13927_/Q vssd1 vssd1 vccd1 vccd1 _11140_/B sky130_fd_sc_hd__clkbuf_1
X_11889_ _13811_/Q _11882_/X _11887_/X _11888_/Y _11885_/X vssd1 vssd1 vccd1 vccd1
+ _13751_/D sky130_fd_sc_hd__o221a_1
XANTENNA__12348__A _12348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13628_ input87/X _14433_/Q _13628_/S vssd1 vssd1 vccd1 vccd1 _13629_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09426__B1 _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13559_ _12664_/X _14413_/Q _13559_/S vssd1 vssd1 vccd1 vccd1 _13560_/B sky130_fd_sc_hd__mux2_1
X_07080_ _14267_/Q _07046_/X _07079_/X _14363_/Q vssd1 vssd1 vccd1 vccd1 _07080_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14265__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12083__A _12536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07982_ _09286_/B vssd1 vssd1 vccd1 vccd1 _08573_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_114_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06963__A1 _14282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06933_ _14286_/Q _06929_/X _06932_/X _14382_/Q vssd1 vssd1 vccd1 vccd1 _06933_/X
+ sky130_fd_sc_hd__o211a_1
X_09721_ _09614_/Y _09721_/B vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__and2b_1
XFILLER_45_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11839__A2 _11855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08704__A2 _09000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06864_ _13777_/Q vssd1 vssd1 vccd1 vccd1 _06864_/Y sky130_fd_sc_hd__inv_2
X_09652_ _09652_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09663_/A sky130_fd_sc_hd__xnor2_2
XFILLER_41_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08603_ _09132_/B vssd1 vssd1 vccd1 vccd1 _09053_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_94_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09583_ _09538_/A _09538_/B _09582_/X vssd1 vssd1 vccd1 vccd1 _09712_/B sky130_fd_sc_hd__a21boi_1
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08534_ _08534_/A _08537_/A _08534_/C vssd1 vssd1 vccd1 vccd1 _08566_/B sky130_fd_sc_hd__nand3_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08465_ _08468_/B _08815_/B _08703_/B _08925_/A vssd1 vssd1 vccd1 vccd1 _08469_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_24_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12258__A _12259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07416_ _07431_/A _07416_/B vssd1 vssd1 vccd1 vccd1 _07416_/X sky130_fd_sc_hd__or2_1
XFILLER_50_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08396_ _09685_/A _08389_/B _08388_/A vssd1 vssd1 vccd1 vccd1 _08402_/B sky130_fd_sc_hd__a21oi_1
XFILLER_17_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07347_ _07373_/A vssd1 vssd1 vccd1 vccd1 _07347_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_36_io_wbs_clk_A clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_12_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07278_ _07300_/B _14166_/Q _07278_/C vssd1 vssd1 vccd1 vccd1 _07307_/C sky130_fd_sc_hd__nor3_1
XFILLER_12_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09017_ _08135_/A _08925_/C _08547_/D _08208_/B vssd1 vssd1 vccd1 vccd1 _09017_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11527__A1 _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07087__A _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08943__A2 _08937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12721__A _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07815__A _14037_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _09938_/A _09938_/B _09918_/Y vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__a21oi_2
XFILLER_58_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12930_ _12930_/A _12940_/B vssd1 vssd1 vccd1 vccd1 _12930_/X sky130_fd_sc_hd__or2_1
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _14133_/Q _12857_/X _12860_/X _12817_/X vssd1 vssd1 vccd1 vccd1 _14133_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _13787_/Q _11848_/A _11770_/X _14236_/Q vssd1 vssd1 vccd1 vccd1 _11812_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _14138_/Q _12776_/X _12791_/X vssd1 vssd1 vccd1 vccd1 _12792_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__A _14256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _13823_/Q _11718_/X _11740_/B vssd1 vssd1 vccd1 vccd1 _11743_/X sky130_fd_sc_hd__o21ba_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14464_/CLK _14462_/D vssd1 vssd1 vccd1 vccd1 _14462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _13773_/Q _13771_/Q vssd1 vssd1 vccd1 vccd1 _11679_/B sky130_fd_sc_hd__or2b_1
XFILLER_14_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14288__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13698__S _13704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13413_ _12688_/X _14371_/Q _13425_/S vssd1 vssd1 vccd1 vccd1 _13414_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10625_ _10626_/A _10626_/B _10528_/X vssd1 vssd1 vccd1 vccd1 _10625_/X sky130_fd_sc_hd__a21o_1
X_14393_ _14440_/CLK _14393_/D vssd1 vssd1 vccd1 vccd1 _14393_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13344_ _14351_/Q _13332_/X _13342_/X _13343_/X vssd1 vssd1 vccd1 vccd1 _14351_/D
+ sky130_fd_sc_hd__o211a_1
X_10556_ _10556_/A _10556_/B vssd1 vssd1 vccd1 vccd1 _10556_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13275_ _14448_/Q _13315_/A _13204_/X _14400_/Q vssd1 vssd1 vccd1 vccd1 _13275_/X
+ sky130_fd_sc_hd__a22o_1
X_10487_ _10487_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__nor2_1
X_12226_ _13079_/A _12226_/B vssd1 vssd1 vccd1 vccd1 _12229_/S sky130_fd_sc_hd__or2_1
XFILLER_5_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12157_ _12909_/A _12160_/B vssd1 vssd1 vccd1 vccd1 _12157_/X sky130_fd_sc_hd__or2_1
XFILLER_29_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11108_ _11108_/A _11108_/B vssd1 vssd1 vccd1 vccd1 _11108_/Y sky130_fd_sc_hd__nor2_1
X_12088_ _13470_/A vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11039_ _11039_/A _11039_/B vssd1 vssd1 vccd1 vccd1 _11050_/B sky130_fd_sc_hd__xor2_1
XFILLER_83_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10151__A _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07460__A _07460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07122__A1 _14294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08250_ _09762_/A _08621_/A vssd1 vssd1 vccd1 vccd1 _08252_/B sky130_fd_sc_hd__or2_1
X_07201_ _14277_/Q _07200_/X _07201_/S vssd1 vssd1 vccd1 vccd1 _07202_/A sky130_fd_sc_hd__mux2_1
X_08181_ _09696_/A vssd1 vssd1 vccd1 vccd1 _09635_/A sky130_fd_sc_hd__clkbuf_4
X_07132_ _14423_/Q _07131_/Y _06970_/A vssd1 vssd1 vccd1 vccd1 _07132_/X sky130_fd_sc_hd__a21o_1
X_07063_ _14436_/Q _14260_/Q vssd1 vssd1 vccd1 vccd1 _07063_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11509__A1 _10215_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08386__B1 _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08138__A1_N _08621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13637__A _13637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09553__C _09553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _07966_/A _07963_/Y _08002_/A _08684_/A vssd1 vssd1 vccd1 vccd1 _08315_/A
+ sky130_fd_sc_hd__and4bb_1
X_09704_ _09692_/A _09692_/Y _09702_/X _09703_/Y vssd1 vssd1 vccd1 vccd1 _09704_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10061__A _10061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06916_ _14432_/Q _06915_/Y _06877_/X vssd1 vssd1 vccd1 vccd1 _06916_/X sky130_fd_sc_hd__a21o_1
XFILLER_96_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07896_ _07896_/A _07843_/Y vssd1 vssd1 vccd1 vccd1 _07897_/B sky130_fd_sc_hd__or2b_1
XANTENNA__09850__A _10127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09635_ _09635_/A _09635_/B vssd1 vssd1 vccd1 vccd1 _09635_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09566_ _09592_/B _09592_/C _09592_/A vssd1 vssd1 vccd1 vccd1 _09566_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08466__A _14011_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10248__A1 _08980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ _08517_/A _08517_/B _08517_/C vssd1 vssd1 vccd1 vccd1 _08532_/A sky130_fd_sc_hd__nand3_1
XFILLER_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09497_ _09541_/B _09496_/C _09496_/A vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08448_ _09807_/B vssd1 vssd1 vccd1 vccd1 _09011_/B sky130_fd_sc_hd__buf_2
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _09678_/A _09678_/B _09678_/C vssd1 vssd1 vccd1 vccd1 _08379_/Y sky130_fd_sc_hd__nand3_2
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11748__A1 _11745_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10410_ _10459_/B _10411_/A vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__or2b_1
XANTENNA__09297__A _09297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ _13847_/Q _11390_/B vssd1 vssd1 vccd1 vccd1 _11390_/X sky130_fd_sc_hd__or2_1
XFILLER_87_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08632__C _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10341_ _10341_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10345_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ _11990_/B _13059_/A _13059_/B _14240_/Q vssd1 vssd1 vccd1 vccd1 _13060_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_3_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08351__D _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10272_ _09962_/B _10000_/Y _09999_/Y vssd1 vssd1 vccd1 vccd1 _10272_/X sky130_fd_sc_hd__o21a_1
X_12011_ _13786_/Q _12000_/X _12003_/X _13826_/Q vssd1 vssd1 vccd1 vccd1 _12012_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06927__A1 _14319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07545__A _14256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08129__B1 _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13962_ _14020_/CLK _13962_/D _12384_/Y vssd1 vssd1 vccd1 vccd1 _13962_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12913_ _12913_/A _12913_/B vssd1 vssd1 vccd1 vccd1 _12913_/X sky130_fd_sc_hd__or2_1
X_13893_ _13988_/CLK _13893_/D _12300_/Y vssd1 vssd1 vccd1 vccd1 _13893_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _12847_/A _12844_/B vssd1 vssd1 vccd1 vccd1 _12845_/A sky130_fd_sc_hd__and2_1
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _14150_/Q _12772_/X _12774_/X _14126_/Q vssd1 vssd1 vccd1 vccd1 _12775_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07104__A1 _14264_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_io_wbs_clk clkbuf_opt_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13920_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_30_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _13767_/Q _11729_/B _13768_/Q vssd1 vssd1 vccd1 vccd1 _11726_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14445_ _14449_/CLK _14445_/D vssd1 vssd1 vccd1 vccd1 _14445_/Q sky130_fd_sc_hd__dfxtp_1
X_11657_ _13778_/Q _13777_/Q _13776_/Q _13775_/Q vssd1 vssd1 vccd1 vccd1 _11675_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_7_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10608_ _10615_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10608_/X sky130_fd_sc_hd__or2b_1
XFILLER_70_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14376_ _14457_/CLK _14376_/D vssd1 vssd1 vccd1 vccd1 _14376_/Q sky130_fd_sc_hd__dfxtp_1
X_11588_ _11587_/A _11587_/B _11587_/C vssd1 vssd1 vccd1 vccd1 _11588_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _13526_/A vssd1 vssd1 vccd1 vccd1 _13327_/X sky130_fd_sc_hd__clkbuf_2
X_10539_ _09725_/X _09741_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _10540_/B sky130_fd_sc_hd__a21oi_2
XFILLER_50_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13258_ _13299_/A vssd1 vssd1 vccd1 vccd1 _13258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12209_ _12904_/A vssd1 vssd1 vccd1 vccd1 _12209_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10580__S _10585_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09654__B _09663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12361__A _12379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13189_ _13189_/A vssd1 vssd1 vccd1 vccd1 _13189_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07750_ _14065_/Q _07720_/X _07748_/X _07749_/Y vssd1 vssd1 vccd1 vccd1 _14065_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07681_ _14125_/Q _14060_/Q vssd1 vssd1 vccd1 vccd1 _07682_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_65_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14259_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13192__A _13193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09420_ _09420_/A _09420_/B vssd1 vssd1 vccd1 vccd1 _10613_/C sky130_fd_sc_hd__nor2_8
XFILLER_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09351_ _09351_/A _09351_/B _09351_/C vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__or3_1
XFILLER_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08302_ _09336_/A _08334_/B vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__nor2_1
XFILLER_61_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09282_ _09425_/A _08449_/C _09281_/A _09281_/C vssd1 vssd1 vccd1 vccd1 _09284_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08233_ _08403_/A _08233_/B vssd1 vssd1 vccd1 vccd1 _08234_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12536__A _12536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08733__B _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08164_ _09590_/A vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07115_ _07112_/X _14295_/Q _07115_/S vssd1 vssd1 vccd1 vccd1 _07116_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ _09465_/A vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__inv_2
XFILLER_119_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07046_ _07085_/A vssd1 vssd1 vccd1 vccd1 _07046_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12155__A1 _13824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06909__A1 _14262_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08997_ _08997_/A _08997_/B vssd1 vssd1 vccd1 vccd1 _09023_/A sky130_fd_sc_hd__and2_1
XFILLER_60_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07948_ _08976_/A vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__buf_4
XFILLER_21_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09580__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07879_ _07877_/Y _13981_/Q _07912_/S vssd1 vssd1 vccd1 vccd1 _07880_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09618_ _09575_/X _09622_/A _09721_/B _09617_/Y vssd1 vssd1 vccd1 vccd1 _09667_/A
+ sky130_fd_sc_hd__o211a_1
X_10890_ _13973_/Q _10900_/B vssd1 vssd1 vccd1 vccd1 _10890_/X sky130_fd_sc_hd__and2_1
XFILLER_93_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09549_ _09549_/A _09549_/B vssd1 vssd1 vccd1 vccd1 _09592_/A sky130_fd_sc_hd__xor2_1
XFILLER_34_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12560_ _12560_/A vssd1 vssd1 vccd1 vccd1 _14021_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ _11511_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11511_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10641__A1 _13953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12491_ _14036_/Q _12485_/X _12490_/X _12473_/X vssd1 vssd1 vccd1 vccd1 _12491_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14230_ _14244_/CLK _14230_/D _13028_/Y vssd1 vssd1 vccd1 vccd1 _14230_/Q sky130_fd_sc_hd__dfrtp_2
X_11442_ _11442_/A vssd1 vssd1 vccd1 vccd1 _11471_/B sky130_fd_sc_hd__inv_2
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14161_ _14163_/CLK _14161_/D vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_2
X_11373_ _13854_/Q _11377_/B vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__or2_1
X_13112_ _13112_/A vssd1 vssd1 vccd1 vccd1 _14257_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input60_A io_wbs_adr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ _10346_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10326_/A sky130_fd_sc_hd__xnor2_1
X_14092_ _14104_/CLK _14092_/D _12740_/Y vssd1 vssd1 vccd1 vccd1 _14092_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13043_ _14244_/Q _13036_/S _13042_/Y hold34/A _13032_/X vssd1 vssd1 vccd1 vccd1
+ _13043_/X sky130_fd_sc_hd__a221o_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10255_/A _10255_/B vssd1 vssd1 vccd1 vccd1 _10619_/A sky130_fd_sc_hd__or2_1
XFILLER_65_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10186_ _10186_/A _10186_/B vssd1 vssd1 vccd1 vccd1 _10186_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_output147_A _14303_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09314__A2 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13945_ _13946_/CLK _13945_/D _12364_/Y vssd1 vssd1 vccd1 vccd1 _13945_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13876_ _14028_/CLK _13876_/D _12278_/Y vssd1 vssd1 vccd1 vccd1 _13876_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09078__A1 _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ input66/X vssd1 vssd1 vccd1 vccd1 _12827_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_61_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12758_/A vssd1 vssd1 vccd1 vccd1 _12758_/Y sky130_fd_sc_hd__inv_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11709_ _13772_/Q _11706_/Y _11708_/Y vssd1 vssd1 vccd1 vccd1 _13772_/D sky130_fd_sc_hd__a21oi_1
X_12689_ _12688_/X _14055_/Q _12695_/S vssd1 vssd1 vccd1 vccd1 _12690_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12356__A _12360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11260__A _13895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14428_ _14465_/CLK _14428_/D vssd1 vssd1 vccd1 vccd1 _14428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14359_ _14365_/CLK _14359_/D vssd1 vssd1 vccd1 vccd1 _14359_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_115_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08920_ _08934_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08921_/B sky130_fd_sc_hd__and2_1
XFILLER_112_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10604__A _10604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07185__A _07185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ _08811_/Y _08840_/X _08883_/A _08850_/X vssd1 vssd1 vccd1 vccd1 _08858_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_44_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09295__B_N _09223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _11175_/S vssd1 vssd1 vccd1 vccd1 _10670_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08782_ _09943_/B vssd1 vssd1 vccd1 vccd1 _08937_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_38_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07733_ _07732_/Y _14158_/Q _07757_/S vssd1 vssd1 vccd1 vccd1 _07733_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07664_ _14068_/Q _07664_/B vssd1 vssd1 vccd1 vccd1 _07665_/B sky130_fd_sc_hd__or2_1
XFILLER_26_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09403_ _09396_/Y _09397_/X _09329_/A _09329_/Y vssd1 vssd1 vccd1 vccd1 _09404_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_77_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07595_ _07595_/A vssd1 vssd1 vccd1 vccd1 _07604_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_81_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09334_ _09319_/A _09242_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _09335_/B sky130_fd_sc_hd__o21ba_1
XFILLER_51_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10623__A1 _10565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11820__B1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _09187_/X _09190_/Y _09262_/X _09264_/Y vssd1 vssd1 vccd1 vccd1 _09267_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_21_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08216_ _08217_/B _08217_/C _08217_/A vssd1 vssd1 vccd1 vccd1 _08218_/A sky130_fd_sc_hd__a21o_1
X_09196_ _09340_/A _09340_/B vssd1 vssd1 vccd1 vccd1 _09341_/B sky130_fd_sc_hd__xnor2_1
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _08622_/A vssd1 vssd1 vccd1 vccd1 _08317_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__07252__A0 _14078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08078_ _08078_/A _08078_/B _08078_/C vssd1 vssd1 vccd1 vccd1 _08079_/B sky130_fd_sc_hd__or3_1
XFILLER_84_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07029_ _07012_/X _07028_/X _14370_/Q vssd1 vssd1 vccd1 vccd1 _07030_/S sky130_fd_sc_hd__o21a_1
XANTENNA__10514__A _10644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__A2_N _11882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10040_ _09930_/B _10067_/B _10039_/X vssd1 vssd1 vccd1 vccd1 _10042_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__buf_2
XFILLER_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07823__A _14032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11991_ hold6/A _13823_/Q _11991_/S vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13730_ _13730_/A vssd1 vssd1 vccd1 vccd1 _14462_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10942_ _10715_/A _10927_/Y _10941_/X vssd1 vssd1 vccd1 vccd1 _11026_/A sky130_fd_sc_hd__a21bo_1
XFILLER_44_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10862__A1 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13661_ _13661_/A _13661_/B vssd1 vssd1 vccd1 vccd1 _13662_/A sky130_fd_sc_hd__and2_1
XFILLER_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10873_ _10873_/A _10873_/B _10873_/C vssd1 vssd1 vccd1 vccd1 _10874_/B sky130_fd_sc_hd__nor3_1
XFILLER_44_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ _13184_/A _12612_/B vssd1 vssd1 vccd1 vccd1 _12613_/A sky130_fd_sc_hd__or2_1
XANTENNA__12064__B1 _12060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13592_ _13592_/A vssd1 vssd1 vccd1 vccd1 _13607_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12543_ _12543_/A vssd1 vssd1 vccd1 vccd1 _14016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09480__A1 _08623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09480__B2 _08623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12474_ _14032_/Q _12464_/X _12472_/X _12473_/X vssd1 vssd1 vccd1 vccd1 _12474_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_71_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14213_ _14215_/CLK _14213_/D _13007_/Y vssd1 vssd1 vccd1 vccd1 _14213_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09768__C1 _10393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ _11282_/A _11061_/A _11425_/S vssd1 vssd1 vccd1 vccd1 _11426_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12904__A _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07243__A0 _14081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14144_ _14149_/CLK _14144_/D vssd1 vssd1 vccd1 vccd1 _14144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11356_ _11355_/A _10845_/X _11355_/Y _10669_/X vssd1 vssd1 vccd1 vccd1 _13894_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10307_ _10307_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10307_/X sky130_fd_sc_hd__and2_1
XFILLER_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14075_ _14075_/CLK _14075_/D _12719_/Y vssd1 vssd1 vccd1 vccd1 _14075_/Q sky130_fd_sc_hd__dfrtp_1
X_11287_ _11333_/B _11333_/C _11333_/A vssd1 vssd1 vccd1 vccd1 _11334_/A sky130_fd_sc_hd__a21o_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _13028_/A vssd1 vssd1 vccd1 vccd1 _13026_/Y sky130_fd_sc_hd__inv_2
X_10238_ _10151_/X _10169_/Y _10185_/Y _10186_/Y vssd1 vssd1 vccd1 vccd1 _10238_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07546__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10169_ _10186_/A _10186_/B _10168_/X vssd1 vssd1 vccd1 vccd1 _10169_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13928_ _13987_/CLK _13928_/D _12343_/Y vssd1 vssd1 vccd1 vccd1 _13928_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13859_ _13867_/CLK _13859_/D _12256_/Y vssd1 vssd1 vccd1 vccd1 _13859_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13470__A _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07380_ _07376_/X _07377_/X _07378_/X _07379_/X vssd1 vssd1 vccd1 vccd1 _07380_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09050_ _09050_/A _09188_/C vssd1 vssd1 vccd1 vccd1 _09110_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13555__A0 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08001_ _08291_/C vssd1 vssd1 vccd1 vccd1 _08132_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_7_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07908__A _14027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09952_ _10013_/A _10013_/B _09951_/X vssd1 vssd1 vccd1 vccd1 _09954_/B sky130_fd_sc_hd__a21oi_1
XFILLER_103_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08903_ _09044_/A _10215_/B _08906_/A _08902_/X vssd1 vssd1 vccd1 vccd1 _08957_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09883_ _09975_/B vssd1 vssd1 vccd1 vccd1 _09883_/Y sky130_fd_sc_hd__inv_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12530__A1 _08983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08834_ _08834_/A _08834_/B _08834_/C vssd1 vssd1 vccd1 vccd1 _08844_/B sky130_fd_sc_hd__and3_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08765_ _08771_/A vssd1 vssd1 vccd1 vccd1 _08772_/A sky130_fd_sc_hd__inv_2
XFILLER_73_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _07716_/A _07716_/B vssd1 vssd1 vccd1 vccd1 _07716_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08696_ _09348_/B _09865_/A _09884_/A _08750_/A vssd1 vssd1 vccd1 vccd1 _08745_/C
+ sky130_fd_sc_hd__a22o_1
X_07647_ _14072_/Q _14071_/Q _07660_/A vssd1 vssd1 vccd1 vccd1 _07716_/A sky130_fd_sc_hd__and3_2
XFILLER_54_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07578_ _14093_/Q input9/X _07582_/S vssd1 vssd1 vccd1 vccd1 _07579_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12597__A1 _14032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_3_0_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_io_wbs_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_09317_ _08978_/B _08284_/C _08070_/C _08978_/A vssd1 vssd1 vccd1 vccd1 _09317_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_90_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09248_ _09248_/A _09248_/B _09248_/C vssd1 vssd1 vccd1 vccd1 _09248_/X sky130_fd_sc_hd__and3_1
XANTENNA__13546__A0 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ _09177_/X _09176_/Y _09144_/Y _09144_/B vssd1 vssd1 vccd1 vccd1 _09180_/D
+ sky130_fd_sc_hd__o211ai_2
XFILLER_108_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11210_ _13907_/Q vssd1 vssd1 vccd1 vccd1 _11300_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12190_ _12828_/B vssd1 vssd1 vccd1 vccd1 _13194_/C sky130_fd_sc_hd__inv_2
XANTENNA__07818__A _14035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11141_ _10761_/B _11139_/X _11140_/X vssd1 vssd1 vccd1 vccd1 _11141_/X sky130_fd_sc_hd__o21a_1
X_11072_ _11107_/B _11112_/B _11107_/A vssd1 vssd1 vccd1 vccd1 _11108_/B sky130_fd_sc_hd__o21a_1
Xinput100 io_wbs_we vssd1 vssd1 vccd1 vccd1 _12211_/A sky130_fd_sc_hd__buf_4
XFILLER_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10023_ _10055_/A _10021_/X _10216_/A vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__a21boi_2
XFILLER_1_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08649__A _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input23_A dout1[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_43_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_5_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11974_ _11976_/A vssd1 vssd1 vccd1 vccd1 _11974_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13713_ _13713_/A vssd1 vssd1 vccd1 vccd1 _14457_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08087__C _08097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10925_ _10652_/A _10924_/X _10920_/X vssd1 vssd1 vccd1 vccd1 _10990_/A sky130_fd_sc_hd__o21ai_2
XFILLER_60_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13644_ _13644_/A _13644_/B vssd1 vssd1 vccd1 vccd1 _13645_/A sky130_fd_sc_hd__and2_1
X_10856_ _13938_/Q _10855_/X _10871_/S vssd1 vssd1 vccd1 vccd1 _10857_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13592_/A vssd1 vssd1 vccd1 vccd1 _13590_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10599__B1 _10562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ _10899_/A _10899_/B vssd1 vssd1 vccd1 vccd1 _10894_/B sky130_fd_sc_hd__or2_1
XANTENNA__10419__A _10435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12526_ _12526_/A vssd1 vssd1 vccd1 vccd1 _14011_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12457_ _13731_/A vssd1 vssd1 vccd1 vccd1 _12817_/A sky130_fd_sc_hd__buf_2
XANTENNA__07216__A0 _14273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _13876_/Q _11392_/A _11396_/A _11407_/X vssd1 vssd1 vccd1 vccd1 _13876_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09756__A2 _08255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12388_ _12391_/A vssd1 vssd1 vccd1 vccd1 _12388_/Y sky130_fd_sc_hd__inv_2
X_14127_ _14152_/CLK _14127_/D vssd1 vssd1 vccd1 vccd1 _14127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11339_ _11339_/A _11339_/B vssd1 vssd1 vccd1 vccd1 _11339_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_99_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09943__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14058_ _14256_/CLK _14255_/Q _12698_/Y vssd1 vssd1 vccd1 vccd1 _14058_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12512__A1 _08966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13465__A _13485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ _13009_/A vssd1 vssd1 vccd1 vccd1 _13009_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06880_ _14391_/Q vssd1 vssd1 vccd1 vccd1 _06880_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08550_ _08584_/A _08550_/B vssd1 vssd1 vccd1 vccd1 _08568_/A sky130_fd_sc_hd__or2_1
XFILLER_36_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07501_ _07501_/A _07501_/B vssd1 vssd1 vccd1 vccd1 _14187_/D sky130_fd_sc_hd__nand2_1
X_08481_ _09865_/B vssd1 vssd1 vccd1 vccd1 _09905_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07432_ _11746_/S vssd1 vssd1 vccd1 vccd1 _07432_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ _07363_/A vssd1 vssd1 vccd1 vccd1 _07363_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09444__B2 _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09102_ _09144_/A _09144_/B _09144_/C vssd1 vssd1 vccd1 vccd1 _09102_/X sky130_fd_sc_hd__and3_1
X_07294_ _14227_/Q vssd1 vssd1 vccd1 vccd1 _07333_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_108_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09033_ _09030_/Y _09031_/Y _08678_/A _08967_/X vssd1 vssd1 vccd1 vccd1 _09033_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_11_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07207__A0 _14276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13359__B _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09935_ _09978_/A _09933_/B _10394_/B vssd1 vssd1 vccd1 vccd1 _09935_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12503__A1 _14056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09866_ _09866_/A _09905_/A vssd1 vssd1 vccd1 vccd1 _09866_/X sky130_fd_sc_hd__and2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _08814_/X _08815_/X _08818_/A _08816_/Y vssd1 vssd1 vccd1 vccd1 _08856_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_86_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09797_ _08291_/C _09824_/B _09796_/X vssd1 vssd1 vccd1 vccd1 _09799_/A sky130_fd_sc_hd__a21o_1
XFILLER_2_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08748_ _08789_/A _08748_/B vssd1 vssd1 vccd1 vccd1 _08787_/B sky130_fd_sc_hd__nand2_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _08980_/B vssd1 vssd1 vccd1 vccd1 _10486_/S sky130_fd_sc_hd__buf_6
XANTENNA__12719__A _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _13941_/Q vssd1 vssd1 vccd1 vccd1 _10716_/A sky130_fd_sc_hd__inv_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _13766_/Q _11732_/B vssd1 vssd1 vccd1 vccd1 _11729_/B sky130_fd_sc_hd__or2_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10641_ _13953_/Q _10550_/X _10634_/Y _10640_/X vssd1 vssd1 vccd1 vccd1 _13953_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13231__A2 _13336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13360_ _13447_/A vssd1 vssd1 vccd1 vccd1 _13467_/S sky130_fd_sc_hd__buf_6
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10572_ _10572_/A _10572_/B vssd1 vssd1 vccd1 vccd1 _10572_/Y sky130_fd_sc_hd__xnor2_1
X_12311_ _12317_/A vssd1 vssd1 vccd1 vccd1 _12316_/A sky130_fd_sc_hd__buf_2
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13291_ _14371_/Q _13215_/A _13299_/A vssd1 vssd1 vccd1 vccd1 _13291_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08651__B _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12242_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08370__C _13874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12173_ _12922_/A _12173_/B vssd1 vssd1 vccd1 vccd1 _12173_/X sky130_fd_sc_hd__or2_1
XANTENNA__07267__B _14166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11124_ _11124_/A _11124_/B _11124_/C vssd1 vssd1 vccd1 vccd1 _11124_/X sky130_fd_sc_hd__or3_1
XFILLER_111_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11055_ _11124_/B _11124_/C _11124_/A vssd1 vssd1 vccd1 vccd1 _11125_/B sky130_fd_sc_hd__o21a_1
XFILLER_114_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09482__B _09482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10006_ _10382_/B _10006_/B vssd1 vssd1 vccd1 vccd1 _10011_/A sky130_fd_sc_hd__xnor2_1
XFILLER_92_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10421__B _10421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11957_ _11959_/A vssd1 vssd1 vccd1 vccd1 _11957_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08826__B _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11481__A1 _08658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10908_ _13970_/Q _10690_/S _10904_/X _13928_/Q _10907_/X vssd1 vssd1 vccd1 vccd1
+ _13928_/D sky130_fd_sc_hd__o221a_1
XFILLER_33_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11888_ _13751_/Q _11888_/B vssd1 vssd1 vccd1 vccd1 _11888_/Y sky130_fd_sc_hd__nor2_1
X_13627_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13644_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10839_ _10839_/A vssd1 vssd1 vccd1 vccd1 _13941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13558_ _13592_/A vssd1 vssd1 vccd1 vccd1 _13573_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08842__A _08842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12509_ _12209_/X _12210_/X _12567_/B _12508_/X _12216_/X vssd1 vssd1 vccd1 vccd1
+ _14007_/D sky130_fd_sc_hd__o311a_1
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13489_ _13502_/A _13489_/B vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__and2_1
XFILLER_69_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12364__A _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09673__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ _14019_/Q vssd1 vssd1 vccd1 vccd1 _09286_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13195__A _13332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ _09720_/A _09720_/B vssd1 vssd1 vccd1 vccd1 _09723_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06932_ _14430_/Q _06930_/Y _06931_/X vssd1 vssd1 vccd1 vccd1 _06932_/X sky130_fd_sc_hd__a21o_1
XFILLER_68_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09651_ _09651_/A _09647_/C vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__or2b_1
X_06863_ _14402_/Q _06856_/Y _11659_/A _14401_/Q _06862_/X vssd1 vssd1 vccd1 vccd1
+ _06869_/B sky130_fd_sc_hd__a221o_1
XFILLER_28_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08602_ _09055_/A _08684_/A vssd1 vssd1 vccd1 vccd1 _08607_/A sky130_fd_sc_hd__nand2_1
XFILLER_95_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09582_ _09582_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__or2b_1
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07921__A _14024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ _08590_/B _08502_/C _08502_/B vssd1 vssd1 vccd1 vccd1 _08534_/C sky130_fd_sc_hd__a21o_1
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08464_ _09132_/A vssd1 vssd1 vccd1 vccd1 _08925_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07415_ _14206_/Q _14208_/Q _07415_/S vssd1 vssd1 vccd1 vccd1 _07416_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08395_ _09696_/A vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_32_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_1_0_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_io_wbs_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07346_ _14220_/Q _07311_/X _07316_/X _07345_/X vssd1 vssd1 vccd1 vccd1 _14220_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09848__A _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07277_ _14191_/Q _07312_/A _07277_/C _14225_/Q vssd1 vssd1 vccd1 vccd1 _07278_/C
+ sky130_fd_sc_hd__or4b_1
XANTENNA__12274__A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09016_ _09084_/C _09084_/D vssd1 vssd1 vccd1 vccd1 _10092_/A sky130_fd_sc_hd__nand2_4
XFILLER_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07600__A0 _14083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09918_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09918_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10522__A _10644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09849_ _08836_/B _09847_/X _09848_/X vssd1 vssd1 vccd1 vccd1 _09895_/A sky130_fd_sc_hd__o21ai_4
XFILLER_59_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12860_ _12904_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _12860_/X sky130_fd_sc_hd__or2_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _13993_/Q _11845_/B _12254_/B _14112_/Q vssd1 vssd1 vccd1 vccd1 _11811_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07831__A _14024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12809_/A vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09656__A1 _10644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _13764_/Q _11714_/X _11716_/A _11741_/X vssd1 vssd1 vccd1 vccd1 _13764_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11463__A1 _09188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_16_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13987_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14465_/CLK _14461_/D vssd1 vssd1 vccd1 vccd1 _14461_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11673_/A vssd1 vssd1 vccd1 vccd1 _13780_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _13447_/A vssd1 vssd1 vccd1 vccd1 _13425_/S sky130_fd_sc_hd__buf_2
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input90_A io_wbs_datwr[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06890__A1 _14393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ _13955_/Q _10545_/X _10623_/X vssd1 vssd1 vccd1 vccd1 _13955_/D sky130_fd_sc_hd__o21a_1
X_14392_ _14440_/CLK _14392_/D vssd1 vssd1 vccd1 vccd1 _14392_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_70_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13343_ _13343_/A vssd1 vssd1 vccd1 vccd1 _13343_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10555_ _10418_/A _10417_/A _10565_/C _10644_/A vssd1 vssd1 vccd1 vccd1 _10556_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12184__A input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13274_ _13637_/A vssd1 vssd1 vccd1 vccd1 _13315_/A sky130_fd_sc_hd__clkbuf_2
X_10486_ _09998_/A _09188_/B _10486_/S vssd1 vssd1 vccd1 vccd1 _10487_/B sky130_fd_sc_hd__mux2_1
XANTENNA_output177_A _14168_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12225_ _12906_/A _12220_/S _12224_/Y vssd1 vssd1 vccd1 vccd1 _13837_/D sky130_fd_sc_hd__o21a_1
X_12156_ input88/X vssd1 vssd1 vccd1 vccd1 _12909_/A sky130_fd_sc_hd__buf_6
XFILLER_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11107_ _11107_/A _11107_/B _11112_/B vssd1 vssd1 vccd1 vccd1 _11107_/X sky130_fd_sc_hd__or3_1
XFILLER_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12087_ input33/X input44/X _13202_/A _12429_/A vssd1 vssd1 vccd1 vccd1 _13470_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_1_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11038_ _11038_/A vssd1 vssd1 vccd1 vccd1 _11050_/A sky130_fd_sc_hd__inv_2
XFILLER_65_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_55_io_wbs_clk clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14396_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12989_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12989_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12359__A _12360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12651__A0 _12650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07200_ _14093_/Q _07185_/X _07186_/X vssd1 vssd1 vccd1 vccd1 _07200_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08180_ _09336_/A vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08572__A _13859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07131_ _14455_/Q _14279_/Q vssd1 vssd1 vccd1 vccd1 _07131_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12094__A _12146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07062_ _07062_/A vssd1 vssd1 vccd1 vccd1 _14302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07964_ _09233_/D vssd1 vssd1 vccd1 vccd1 _08684_/A sky130_fd_sc_hd__clkbuf_2
X_09703_ _09727_/B _09727_/C _09727_/A vssd1 vssd1 vccd1 vccd1 _09703_/Y sky130_fd_sc_hd__o21ai_1
X_06915_ _14464_/Q _14288_/Q vssd1 vssd1 vccd1 vccd1 _06915_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09886__A1 _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07895_ _07895_/A vssd1 vssd1 vccd1 vccd1 _13977_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09634_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09634_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09850__B _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09565_ _09592_/A _09592_/B _09592_/C vssd1 vssd1 vccd1 vccd1 _09565_/X sky130_fd_sc_hd__and3_1
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08516_ _08867_/A _09152_/B _08503_/A _08503_/C vssd1 vssd1 vccd1 vccd1 _08517_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12642__A0 _12641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09496_ _09496_/A _09541_/B _09496_/C vssd1 vssd1 vccd1 vccd1 _09496_/X sky130_fd_sc_hd__and3_1
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08447_ _09869_/B vssd1 vssd1 vccd1 vccd1 _09807_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _09678_/C sky130_fd_sc_hd__xor2_2
X_07329_ _07491_/A vssd1 vssd1 vccd1 vccd1 _07329_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10517__A _10629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10340_ _10347_/A _10347_/B vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__xor2_1
XFILLER_87_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10271_ _10271_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10274_/A sky130_fd_sc_hd__nor2_1
X_12010_ _12216_/A vssd1 vssd1 vccd1 vccd1 _12026_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__07826__A _14029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10252__A _10421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08129__A1 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13961_ _14020_/CLK _13961_/D _12383_/Y vssd1 vssd1 vccd1 vccd1 _13961_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12912_ _14152_/Q _12901_/X _12911_/X _12907_/X vssd1 vssd1 vccd1 vccd1 _14152_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13892_ _13892_/CLK _13892_/D _12298_/Y vssd1 vssd1 vccd1 vccd1 _13892_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14255__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ _12641_/X _14129_/Q _12846_/S vssd1 vssd1 vccd1 vccd1 _12844_/B sky130_fd_sc_hd__mux2_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12179__A _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11436__A1 _11002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12774_/A vssd1 vssd1 vccd1 vccd1 _12774_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07104__A2 _07085_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _11716_/X _11722_/X _11724_/X vssd1 vssd1 vccd1 vccd1 _13769_/D sky130_fd_sc_hd__a21o_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12907__A _12920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14444_ _14449_/CLK _14444_/D vssd1 vssd1 vccd1 vccd1 _14444_/Q sky130_fd_sc_hd__dfxtp_1
X_11656_ _11585_/S _11651_/B hold41/X _11655_/X vssd1 vssd1 vccd1 vccd1 _13840_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_70_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10607_ _10626_/A _10261_/X _10263_/Y vssd1 vssd1 vccd1 vccd1 _10615_/B sky130_fd_sc_hd__o21bai_1
X_14375_ _14427_/CLK _14375_/D vssd1 vssd1 vccd1 vccd1 _14375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11587_ _11587_/A _11587_/B _11587_/C vssd1 vssd1 vccd1 vccd1 _11587_/X sky130_fd_sc_hd__or3_1
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09000__B _09000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13326_ _14347_/Q _13311_/X _13325_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _14347_/D
+ sky130_fd_sc_hd__o211a_1
X_10538_ _10457_/A _10456_/A _10548_/C _10528_/A vssd1 vssd1 vccd1 vccd1 _10538_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13257_ _14412_/Q _13230_/X _13256_/X vssd1 vssd1 vccd1 vccd1 _13257_/X sky130_fd_sc_hd__a21o_1
X_10469_ _10407_/A _10472_/S _10439_/A vssd1 vssd1 vccd1 vccd1 _10470_/B sky130_fd_sc_hd__a21oi_1
X_12208_ _13834_/Q _12202_/C _12205_/X _12206_/X _12207_/X vssd1 vssd1 vccd1 vccd1
+ _13834_/D sky130_fd_sc_hd__o221a_1
X_13188_ _13189_/A vssd1 vssd1 vccd1 vccd1 _13188_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12139_ input78/X _12143_/B vssd1 vssd1 vccd1 vccd1 _12139_/X sky130_fd_sc_hd__or2_1
XFILLER_111_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07680_ _07687_/A _07687_/B vssd1 vssd1 vccd1 vccd1 _07680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07471__A _07471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09350_ _08791_/B _09543_/C _09543_/D _08791_/A vssd1 vssd1 vccd1 vccd1 _09351_/C
+ sky130_fd_sc_hd__a22oi_2
X_08301_ _09694_/A _08301_/B vssd1 vssd1 vccd1 vccd1 _08334_/B sky130_fd_sc_hd__xnor2_1
X_09281_ _09281_/A _09281_/B _09281_/C vssd1 vssd1 vccd1 vccd1 _09284_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12817__A _12817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08232_ _09634_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08233_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12927__A1 _14158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13772__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08163_ _08201_/A _08163_/B vssd1 vssd1 vccd1 vccd1 _08167_/C sky130_fd_sc_hd__or2_1
XFILLER_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07114_ _07090_/X _07113_/X _14359_/Q vssd1 vssd1 vccd1 vccd1 _07115_/S sky130_fd_sc_hd__o21a_1
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08094_ _09537_/A vssd1 vssd1 vccd1 vccd1 _09465_/A sky130_fd_sc_hd__clkbuf_4
X_07045_ _07045_/A vssd1 vssd1 vccd1 vccd1 _14304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06909__A2 _06873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08996_ _09045_/A _08994_/Y _08665_/A _08667_/B vssd1 vssd1 vccd1 vccd1 _09025_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_60_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09861__A _10305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07947_ _13871_/Q vssd1 vssd1 vccd1 vccd1 _08976_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07878_ _07878_/A vssd1 vssd1 vccd1 vccd1 _07912_/S sky130_fd_sc_hd__buf_2
XANTENNA__08477__A _13859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09617_ _09614_/Y _09615_/X _09580_/X _09581_/X vssd1 vssd1 vccd1 vccd1 _09617_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_83_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_48_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11418__A1 _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ _09548_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09479_ _09479_/A _09479_/B _09803_/A _09479_/D vssd1 vssd1 vccd1 vccd1 _09481_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_106_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11510_ _11510_/A vssd1 vssd1 vccd1 vccd1 _11510_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12490_ _08150_/A _12486_/X _12476_/X _14052_/Q vssd1 vssd1 vccd1 vccd1 _12490_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12918__A1 _14154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ _11300_/A _11079_/A _11446_/S vssd1 vssd1 vccd1 vccd1 _11442_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08598__A1 _08823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__B2 _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14160_ _14163_/CLK _14160_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_2
X_11372_ _13891_/Q _11363_/X _11370_/X _11371_/X vssd1 vssd1 vccd1 vccd1 _13891_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13111_ _14257_/Q _13111_/B _13111_/C vssd1 vssd1 vccd1 vccd1 _13112_/A sky130_fd_sc_hd__and3b_1
XANTENNA__13558__A _13592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10323_ _10323_/A _10323_/B vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__or2_1
XFILLER_3_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14091_ _14104_/CLK _14091_/D _12739_/Y vssd1 vssd1 vccd1 vccd1 _14091_/Q sky130_fd_sc_hd__dfrtp_1
X_13042_ _13042_/A _13042_/B vssd1 vssd1 vccd1 vccd1 _13042_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_input53_A io_wbs_adr[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10254_ _10254_/A _10254_/B _10254_/C vssd1 vssd1 vccd1 vccd1 _10255_/B sky130_fd_sc_hd__and3_1
XFILLER_106_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11354__B1 _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07022__A1 _14307_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10185_ _10279_/B _10225_/B _10184_/X vssd1 vssd1 vccd1 vccd1 _10185_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_6_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14215_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13944_ _13947_/CLK _13944_/D _12363_/Y vssd1 vssd1 vccd1 vccd1 _13944_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13875_ _13986_/CLK _13875_/D _12277_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12826_ _12209_/X _12210_/X _12900_/B _12825_/Y _12008_/A vssd1 vssd1 vccd1 vccd1
+ _14124_/D sky130_fd_sc_hd__o311a_1
XFILLER_50_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09078__A2 _09076_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13795__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07089__A1 _14266_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _12758_/A vssd1 vssd1 vccd1 vccd1 _12757_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10856__S _10871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11541__A _14052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11708_ _13772_/Q _11706_/Y hold38/X vssd1 vssd1 vccd1 vccd1 _11708_/Y sky130_fd_sc_hd__o21ai_1
X_12688_ input72/X vssd1 vssd1 vccd1 vccd1 _12688_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09011__A _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14427_ _14427_/CLK _14427_/D vssd1 vssd1 vccd1 vccd1 _14427_/Q sky130_fd_sc_hd__dfxtp_1
X_11639_ _11639_/A _11639_/B vssd1 vssd1 vccd1 vccd1 _11639_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_50_io_wbs_clk_A clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14358_ _14365_/CLK _14358_/D vssd1 vssd1 vccd1 vccd1 _14358_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13309_ _14423_/Q _13306_/X _13308_/X _13299_/X vssd1 vssd1 vccd1 vccd1 _13309_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13468__A _13485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14289_ _14365_/CLK _14289_/D _13152_/Y vssd1 vssd1 vccd1 vccd1 _14289_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12372__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09002__A2 _08794_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ _08850_/A _08879_/A _08850_/C vssd1 vssd1 vccd1 vccd1 _08850_/X sky130_fd_sc_hd__and3_1
XANTENNA__08210__B1 _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07801_ _10946_/B vssd1 vssd1 vccd1 vccd1 _11175_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08781_ _08781_/A _08781_/B vssd1 vssd1 vccd1 vccd1 _08962_/A sky130_fd_sc_hd__xor2_1
XFILLER_84_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07732_ _07732_/A vssd1 vssd1 vccd1 vccd1 _07732_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_66_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07663_ _07663_/A _07663_/B vssd1 vssd1 vccd1 vccd1 _07732_/A sky130_fd_sc_hd__or2_2
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09402_ _09402_/A _09644_/B vssd1 vssd1 vccd1 vccd1 _09404_/B sky130_fd_sc_hd__xor2_1
XFILLER_80_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07594_ _07594_/A vssd1 vssd1 vccd1 vccd1 _14086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09333_ _09248_/X _09333_/B vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__and2b_1
XFILLER_90_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ _09263_/X _09261_/Y _09191_/Y _09192_/Y vssd1 vssd1 vccd1 vccd1 _09264_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_21_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08215_ _08215_/A _08247_/B vssd1 vssd1 vccd1 vccd1 _08217_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10067__A _10067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09195_ _09133_/A _09135_/B _09133_/B vssd1 vssd1 vccd1 vccd1 _09340_/B sky130_fd_sc_hd__o21ba_1
XFILLER_88_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09278__D _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _08146_/A vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09856__A _10305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12781__C1 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13378__A _13467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08077_ _08078_/B _08078_/C _08295_/A vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__o21ai_2
XFILLER_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07028_ _14418_/Q _07059_/B _14450_/Q vssd1 vssd1 vccd1 vccd1 _07028_/X sky130_fd_sc_hd__and3b_1
XANTENNA__07376__A _07376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07095__B _14265_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__clkbuf_4
XFILLER_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08979_ _08979_/A _08979_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__nor2_1
XFILLER_5_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11990_ _11994_/A _11990_/B vssd1 vssd1 vccd1 vccd1 _11991_/S sky130_fd_sc_hd__nor2_1
XFILLER_99_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10941_ _10936_/A _10938_/X _10940_/X _10971_/A vssd1 vssd1 vccd1 vccd1 _10941_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08000__A _13872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13660_ input94/X _14442_/Q _13670_/S vssd1 vssd1 vccd1 vccd1 _13661_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10872_ _10872_/A vssd1 vssd1 vccd1 vccd1 _13935_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _12610_/X _14036_/Q _12611_/S vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__mux2_1
X_13591_ _13591_/A vssd1 vssd1 vccd1 vccd1 _14422_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12457__A _13731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12542_ _12551_/A _12542_/B vssd1 vssd1 vccd1 vccd1 _12543_/A sky130_fd_sc_hd__and2_1
XANTENNA__11811__B2 _14112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09480__A2 _09818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12473_ _12473_/A vssd1 vssd1 vccd1 vccd1 _12473_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14212_ _14217_/CLK _14212_/D _13006_/Y vssd1 vssd1 vccd1 vccd1 _14212_/Q sky130_fd_sc_hd__dfrtp_1
X_11424_ _11506_/A _11506_/B vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14443__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14149_/CLK _14143_/D vssd1 vssd1 vccd1 vccd1 _14143_/Q sky130_fd_sc_hd__dfxtp_1
X_11355_ _11355_/A _11355_/B vssd1 vssd1 vccd1 vccd1 _11355_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _10306_/A _10306_/B vssd1 vssd1 vccd1 vccd1 _10338_/A sky130_fd_sc_hd__xnor2_1
X_14074_ _14075_/CLK hold4/X _12718_/Y vssd1 vssd1 vccd1 vccd1 _14074_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11286_ _11330_/B _11286_/B vssd1 vssd1 vccd1 vccd1 _11333_/A sky130_fd_sc_hd__nand2_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ _13028_/A vssd1 vssd1 vccd1 vccd1 _13025_/Y sky130_fd_sc_hd__inv_2
X_10237_ _10204_/Y _10224_/X _10234_/X _10235_/X _10236_/Y vssd1 vssd1 vccd1 vccd1
+ _10237_/X sky130_fd_sc_hd__a32o_2
XFILLER_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12920__A _12920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10168_ _10167_/B _10168_/B vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__and2b_1
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10099_ _10099_/A _10099_/B vssd1 vssd1 vccd1 vccd1 _10100_/B sky130_fd_sc_hd__xnor2_2
XFILLER_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13927_ _13927_/CLK _13927_/D _12341_/Y vssd1 vssd1 vccd1 vccd1 _13927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _14258_/CLK _13858_/D vssd1 vssd1 vccd1 vccd1 _13858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13470__B _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12809_ _12809_/A vssd1 vssd1 vccd1 vccd1 _12809_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12367__A _12379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13789_ _13809_/CLK _13789_/D vssd1 vssd1 vccd1 vccd1 _13789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08000_ _13872_/Q vssd1 vssd1 vccd1 vccd1 _08291_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__08580__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13198__A _13526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13810__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _09950_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09951_/X sky130_fd_sc_hd__and2b_1
XFILLER_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11318__B1 _10851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08902_ _08921_/A _08902_/B vssd1 vssd1 vccd1 vccd1 _08902_/X sky130_fd_sc_hd__and2_1
XFILLER_98_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09882_ _09882_/A _09882_/B vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__xnor2_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12830__A _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08833_ _08820_/A _08820_/B _08820_/C vssd1 vssd1 vccd1 vccd1 _08834_/C sky130_fd_sc_hd__a21o_1
XFILLER_98_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07924__A _09788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13960__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08764_ _08764_/A _08805_/C _08764_/C vssd1 vssd1 vccd1 vccd1 _08771_/A sky130_fd_sc_hd__or3_1
XFILLER_26_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ _07715_/A vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__clkbuf_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13491__A0 _12650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08695_ _13861_/Q vssd1 vssd1 vccd1 vccd1 _09884_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07646_ _14070_/Q _07663_/A vssd1 vssd1 vccd1 vccd1 _07660_/A sky130_fd_sc_hd__and2_1
XFILLER_54_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07577_ _07577_/A vssd1 vssd1 vccd1 vccd1 _14094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12277__A _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09316_ _09316_/A _09316_/B _09316_/C vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__nand3_1
XFILLER_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09247_ _09245_/A _09245_/C _09245_/B vssd1 vssd1 vccd1 vccd1 _09248_/C sky130_fd_sc_hd__a21o_1
XFILLER_108_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09178_ _09144_/B _09144_/Y _09176_/Y _09177_/X vssd1 vssd1 vccd1 vccd1 _09180_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_119_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08129_ _08150_/A _08128_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _08130_/B sky130_fd_sc_hd__o21ai_1
X_11140_ _11152_/S _11140_/B vssd1 vssd1 vccd1 vccd1 _11140_/X sky130_fd_sc_hd__or2_1
XANTENNA__12506__C1 _12498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _11104_/B _11071_/B vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08725__A1 _08966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__nand2_1
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10532__A1 _10528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input16_A dout1[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _11976_/A vssd1 vssd1 vccd1 vccd1 _11973_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13482__B1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10924_ _10765_/B _10923_/X _10916_/X vssd1 vssd1 vccd1 vccd1 _10924_/X sky130_fd_sc_hd__o21a_2
X_13712_ _13712_/A _13712_/B vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__and2_1
XFILLER_44_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13643_ _13084_/X _14437_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13644_/B sky130_fd_sc_hd__mux2_1
X_10855_ _11119_/A _10846_/C _10853_/X _10854_/X vssd1 vssd1 vccd1 vccd1 _10855_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13574_ _13574_/A vssd1 vssd1 vccd1 vccd1 _14417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10599__A1 _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09199__C _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _13929_/Q _10786_/B vssd1 vssd1 vccd1 vccd1 _10899_/B sky130_fd_sc_hd__xnor2_1
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10419__B _10435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12525_ _12534_/A _12525_/B vssd1 vssd1 vccd1 vccd1 _12526_/A sky130_fd_sc_hd__and2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12915__A _12928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12456_ _14028_/Q _12438_/X _12455_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _12456_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07216__A1 _07215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ _13840_/Q _11407_/B vssd1 vssd1 vccd1 vccd1 _11407_/X sky130_fd_sc_hd__or2_1
X_12387_ _12391_/A vssd1 vssd1 vccd1 vccd1 _12387_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10435__A _10435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14126_ _14152_/CLK _14126_/D vssd1 vssd1 vccd1 vccd1 _14126_/Q sky130_fd_sc_hd__dfxtp_1
X_11338_ _11338_/A _11342_/A vssd1 vssd1 vccd1 vccd1 _11339_/B sky130_fd_sc_hd__or2_1
XFILLER_67_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14057_ _14363_/CLK _14057_/D vssd1 vssd1 vccd1 vccd1 _14057_/Q sky130_fd_sc_hd__dfxtp_2
X_11269_ _11269_/A _11269_/B vssd1 vssd1 vccd1 vccd1 _11351_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09943__B _09943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12650__A input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13008_ _13009_/A vssd1 vssd1 vccd1 vccd1 _13008_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13473__B1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07500_ _07274_/A _07399_/A _14187_/Q vssd1 vssd1 vccd1 vccd1 _07501_/B sky130_fd_sc_hd__a21bo_1
XFILLER_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08480_ _13861_/Q vssd1 vssd1 vccd1 vccd1 _09865_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_39_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07431_ _07431_/A _07431_/B vssd1 vssd1 vccd1 vccd1 _07431_/X sky130_fd_sc_hd__or2_1
XFILLER_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07362_ _14217_/Q _07347_/X _07348_/X _07361_/X vssd1 vssd1 vccd1 vccd1 _14217_/D
+ sky130_fd_sc_hd__a22o_1
X_09101_ _09100_/A _09100_/C _09100_/B vssd1 vssd1 vccd1 vccd1 _09144_/C sky130_fd_sc_hd__a21o_1
XANTENNA__07455__A1 _14083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07293_ _07293_/A vssd1 vssd1 vccd1 vccd1 _14228_/D sky130_fd_sc_hd__clkbuf_1
X_09032_ _08678_/A _08967_/X _09030_/Y _09031_/Y vssd1 vssd1 vccd1 vccd1 _09032_/X
+ sky130_fd_sc_hd__a211o_4
XFILLER_50_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07207__A1 _07205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12200__A1 _07323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13656__A _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09934_ _10394_/B _09934_/B vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07654__A _14146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _09865_/A _09865_/B vssd1 vssd1 vccd1 vccd1 _09887_/B sky130_fd_sc_hd__xor2_4
XANTENNA_input8_A dout1[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _08772_/B _08812_/Y _08811_/Y _08811_/A vssd1 vssd1 vccd1 vccd1 _08816_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09796_ _09796_/A _09817_/A vssd1 vssd1 vccd1 vccd1 _09796_/X sky130_fd_sc_hd__and2_1
XFILLER_22_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08747_ _09234_/A _09887_/A _08745_/A _08745_/C vssd1 vssd1 vccd1 vccd1 _08758_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13464__A0 input89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08678_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _08967_/A sky130_fd_sc_hd__nand2_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08485__A _09865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _14126_/Q _14061_/Q vssd1 vssd1 vccd1 vccd1 _07684_/B sky130_fd_sc_hd__nor2_1
XFILLER_41_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_1_io_wbs_clk clkbuf_1_1_1_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_io_wbs_clk/A
+ sky130_fd_sc_hd__clkbuf_2
X_10640_ _10634_/A _10639_/Y _09788_/X vssd1 vssd1 vccd1 vccd1 _10640_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10571_ _10583_/A _10583_/B _10377_/B vssd1 vssd1 vccd1 vccd1 _10572_/B sky130_fd_sc_hd__o21ba_1
X_12310_ _12310_/A vssd1 vssd1 vccd1 vccd1 _12310_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07829__A _14027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ _14451_/Q _13315_/A _13218_/X _14403_/Q vssd1 vssd1 vccd1 vccd1 _13290_/X
+ sky130_fd_sc_hd__a22o_1
X_12241_ _12245_/A vssd1 vssd1 vccd1 vccd1 _12241_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12172_ input95/X vssd1 vssd1 vccd1 vccd1 _12922_/A sky130_fd_sc_hd__buf_6
XANTENNA__07267__C _11663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10753__A1 _11240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ _11119_/X _11120_/C _11122_/X _11100_/X _11056_/A vssd1 vssd1 vccd1 vccd1
+ _13916_/D sky130_fd_sc_hd__a32o_1
XFILLER_110_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054_ _11054_/A _11054_/B vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__xor2_1
XFILLER_77_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10005_ _10205_/A _10017_/B _09872_/A vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__o21ba_2
Xclkbuf_leaf_45_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14464_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output122_A _11849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11956_ _11959_/A vssd1 vssd1 vccd1 vccd1 _11956_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08395__A _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ _10899_/A _10905_/X _11125_/A vssd1 vssd1 vccd1 vccd1 _10907_/X sky130_fd_sc_hd__a21o_1
X_11887_ _13751_/Q _11888_/B vssd1 vssd1 vccd1 vccd1 _11887_/X sky130_fd_sc_hd__and2_1
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13626_ _13626_/A vssd1 vssd1 vccd1 vccd1 _14432_/D sky130_fd_sc_hd__clkbuf_1
X_10838_ _13941_/Q _10836_/X _10871_/S vssd1 vssd1 vccd1 vccd1 _10839_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10149__B _10149_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10769_ _10769_/A _11164_/S vssd1 vssd1 vccd1 vccd1 _10770_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13557_ _13557_/A vssd1 vssd1 vccd1 vccd1 _14412_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12645__A input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08842__B _10171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12508_ _11990_/B _13059_/A _13111_/C _14007_/Q vssd1 vssd1 vccd1 vccd1 _12508_/X
+ sky130_fd_sc_hd__a31o_1
X_13488_ _12645_/X _14393_/Q _13494_/S vssd1 vssd1 vccd1 vccd1 _13489_/B sky130_fd_sc_hd__mux2_1
X_12439_ _12486_/A vssd1 vssd1 vccd1 vccd1 _12439_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13476__A _13485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ _14149_/CLK _14109_/D vssd1 vssd1 vccd1 vccd1 _14109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07980_ _09286_/A vssd1 vssd1 vccd1 vccd1 _08012_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06931_ _06970_/A vssd1 vssd1 vccd1 vccd1 _06931_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13694__A0 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12497__A1 _14038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ _09650_/A _09649_/Y vssd1 vssd1 vccd1 vccd1 _10592_/A sky130_fd_sc_hd__or2b_1
X_06862_ _14401_/Q _11659_/A _06858_/Y _14400_/Q vssd1 vssd1 vccd1 vccd1 _06862_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08601_ _08670_/A _08670_/B vssd1 vssd1 vccd1 vccd1 _08608_/A sky130_fd_sc_hd__xnor2_1
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09581_ _09690_/A _09581_/B vssd1 vssd1 vccd1 vccd1 _09581_/X sky130_fd_sc_hd__or2_1
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08532_ _08532_/A _08719_/A vssd1 vssd1 vccd1 vccd1 _08534_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07125__B1 _06970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _08796_/A vssd1 vssd1 vccd1 vccd1 _09132_/A sky130_fd_sc_hd__buf_2
XFILLER_51_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07414_ _07399_/X _07412_/X _07413_/X _07408_/X _14208_/Q vssd1 vssd1 vccd1 vccd1
+ _14208_/D sky130_fd_sc_hd__a32o_1
X_08394_ _08391_/X _08392_/Y _09698_/A _08390_/Y vssd1 vssd1 vccd1 vccd1 _09729_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_10_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07345_ _07321_/X _07343_/X _07344_/X _07329_/X vssd1 vssd1 vccd1 vccd1 _07345_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09848__B _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07276_ _14190_/Q _07276_/B vssd1 vssd1 vccd1 vccd1 _07277_/C sky130_fd_sc_hd__or2_1
X_09015_ _09015_/A _09015_/B vssd1 vssd1 vccd1 vccd1 _09098_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__14192__D _14192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09864__A _09892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09917_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09938_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12488__A1 _14035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09848_ _09848_/A _09848_/B vssd1 vssd1 vccd1 vccd1 _09848_/X sky130_fd_sc_hd__or2_2
XFILLER_86_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13437__A0 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09779_ _09779_/A _09779_/B vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__xnor2_2
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _12768_/A vssd1 vssd1 vccd1 vccd1 _12254_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _14154_/Q _12783_/X _12774_/X _14130_/Q vssd1 vssd1 vccd1 vccd1 _12790_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _13824_/Q _11718_/X _11739_/X _11740_/Y vssd1 vssd1 vccd1 vccd1 _11741_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11672_ _11669_/X _11672_/B _11680_/D vssd1 vssd1 vccd1 vccd1 _11673_/A sky130_fd_sc_hd__and3b_1
X_14460_ _14465_/CLK _14460_/D vssd1 vssd1 vccd1 vccd1 _14460_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13411_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13426_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__07419__A1 _07399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10623_ _10565_/B _10619_/Y _10622_/Y _09788_/X vssd1 vssd1 vccd1 vccd1 _10623_/X
+ sky130_fd_sc_hd__a211o_1
X_14391_ _14450_/CLK _14391_/D vssd1 vssd1 vccd1 vccd1 _14391_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12465__A _12486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13342_ _14431_/Q _13327_/X _13340_/X _13341_/X vssd1 vssd1 vccd1 vccd1 _13342_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_input83_A io_wbs_datwr[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10554_ _10417_/A _10565_/C _10418_/A vssd1 vssd1 vccd1 vccd1 _10556_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12184__B _13609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13273_ _14335_/Q _13265_/X _13272_/X _13254_/X vssd1 vssd1 vccd1 vccd1 _14335_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07278__B _14166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14184__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10485_ _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__or2_1
XFILLER_108_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_55_io_wbs_clk_A clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12224_ _07263_/A _12220_/S _13193_/A vssd1 vssd1 vccd1 vccd1 _12224_/Y sky130_fd_sc_hd__a21oi_1
X_12155_ _13824_/Q _12146_/X _12154_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _13824_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09493__B _09493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11106_ _11002_/B _10701_/X _11104_/X _11105_/Y vssd1 vssd1 vccd1 vccd1 _13922_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07294__A _14227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12086_ _12086_/A vssd1 vssd1 vccd1 vccd1 _13806_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11037_ _13913_/Q vssd1 vssd1 vccd1 vccd1 _11038_/A sky130_fd_sc_hd__buf_2
XFILLER_65_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07107__B1 _14360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12988_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12988_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07658__A1 _14145_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11939_ _11940_/A vssd1 vssd1 vccd1 vccd1 _11939_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13600__A0 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ _13609_/A vssd1 vssd1 vccd1 vccd1 _13680_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07130_ _07130_/A vssd1 vssd1 vccd1 vccd1 _14293_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08291__C _08291_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07061_ _07058_/X _14302_/Q _07061_/S vssd1 vssd1 vccd1 vccd1 _07062_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13667__A0 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07963_ _08208_/B _09434_/B _08983_/C _08132_/A vssd1 vssd1 vccd1 vccd1 _07963_/Y
+ sky130_fd_sc_hd__a22oi_1
X_06914_ _06914_/A vssd1 vssd1 vccd1 vccd1 _14321_/D sky130_fd_sc_hd__clkbuf_1
X_09702_ _09727_/A _09727_/B _09727_/C vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__or3_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07894_ _07893_/Y _13977_/Q _07912_/S vssd1 vssd1 vccd1 vccd1 _07895_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07932__A _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13419__A0 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09633_ _09631_/A _09631_/Y _09527_/X _09632_/Y vssd1 vssd1 vccd1 vccd1 _09638_/A
+ sky130_fd_sc_hd__a211o_1
X_09564_ _09563_/A _09563_/B _09563_/C vssd1 vssd1 vccd1 vccd1 _09592_/C sky130_fd_sc_hd__a21o_1
XFILLER_110_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08515_ _09234_/A vssd1 vssd1 vccd1 vccd1 _08867_/A sky130_fd_sc_hd__buf_4
XFILLER_70_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09495_ _09541_/A _09494_/B _09491_/Y vssd1 vssd1 vccd1 vccd1 _09496_/C sky130_fd_sc_hd__a21bo_1
XFILLER_93_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08446_ _09508_/B _09882_/A _09092_/C _08445_/X vssd1 vssd1 vccd1 vccd1 _08503_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09859__A _10091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1_0_io_wbs_clk_A clkbuf_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08377_ _08384_/A _08384_/B vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__xor2_2
XFILLER_104_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07328_ _14222_/Q _14224_/Q _07333_/S vssd1 vssd1 vccd1 vccd1 _07328_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07098__B _07098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07259_ _14260_/Q _07258_/X _07259_/S vssd1 vssd1 vccd1 vccd1 _07260_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09594__A _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ _09970_/A _09970_/B _09967_/A vssd1 vssd1 vccd1 vccd1 _10293_/A sky130_fd_sc_hd__o21ai_1
XFILLER_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08129__A2 _08128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13960_ _14020_/CLK _13960_/D _12382_/Y vssd1 vssd1 vccd1 vccd1 _13960_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11133__A1 _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11133__B2 _10826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12911_ _12911_/A _12913_/B vssd1 vssd1 vccd1 vccd1 _12911_/X sky130_fd_sc_hd__or2_1
XFILLER_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13891_ _14107_/CLK _13891_/D _12297_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12842_ _12842_/A vssd1 vssd1 vccd1 vccd1 _14128_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12773_ _12773_/A _13200_/B vssd1 vssd1 vccd1 vccd1 _12774_/A sky130_fd_sc_hd__and2_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11692_/B _11872_/A hold38/A _13769_/Q vssd1 vssd1 vccd1 vccd1 _11724_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14443_ _14449_/CLK _14443_/D vssd1 vssd1 vccd1 vccd1 _14443_/Q sky130_fd_sc_hd__dfxtp_1
X_11655_ _13840_/Q _11655_/B vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__and2_1
XANTENNA__12195__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10606_ _09421_/C _10604_/Y _10605_/Y vssd1 vssd1 vccd1 vccd1 _10606_/X sky130_fd_sc_hd__o21a_1
XFILLER_11_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14374_ _14453_/CLK _14374_/D vssd1 vssd1 vccd1 vccd1 _14374_/Q sky130_fd_sc_hd__dfxtp_1
X_11586_ _11586_/A vssd1 vssd1 vccd1 vccd1 _13857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13325_ _14427_/Q _13306_/X _13324_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13325_/X
+ sky130_fd_sc_hd__a211o_1
X_10537_ _10456_/A _10548_/C _10457_/A vssd1 vssd1 vccd1 vccd1 _10537_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_115_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13256_ _14444_/Q _13250_/X _13245_/X _14396_/Q vssd1 vssd1 vccd1 vccd1 _13256_/X
+ sky130_fd_sc_hd__a22o_1
X_10468_ _10491_/A _10468_/B vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12207_ _12216_/A vssd1 vssd1 vccd1 vccd1 _12207_/X sky130_fd_sc_hd__buf_2
XANTENNA__11539__A _14054_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ _13189_/A vssd1 vssd1 vccd1 vccd1 _13187_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07576__A0 _14094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ _10426_/B _10399_/B vssd1 vssd1 vccd1 vccd1 _10430_/S sky130_fd_sc_hd__xnor2_2
X_12138_ _13818_/Q _12133_/X _12137_/X _12131_/X vssd1 vssd1 vccd1 vccd1 _13818_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09317__A1 _08978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09317__B2 _08978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12069_ _12081_/A _12069_/B vssd1 vssd1 vccd1 vccd1 _12070_/A sky130_fd_sc_hd__and2_1
XFILLER_78_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08300_ _09777_/B _08301_/B vssd1 vssd1 vccd1 vccd1 _08343_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09280_ _09145_/B _09869_/B _08748_/B _09145_/A vssd1 vssd1 vccd1 vccd1 _09281_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08231_ _08245_/A _08169_/B _08168_/A vssd1 vssd1 vccd1 vccd1 _08278_/B sky130_fd_sc_hd__a21oi_1
XFILLER_60_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08162_ _09685_/A vssd1 vssd1 vccd1 vccd1 _08245_/A sky130_fd_sc_hd__buf_2
XFILLER_14_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07113_ _14407_/Q _07134_/B _14439_/Q vssd1 vssd1 vccd1 vccd1 _07113_/X sky130_fd_sc_hd__and3b_1
XFILLER_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08093_ _08093_/A _09319_/A vssd1 vssd1 vccd1 vccd1 _09537_/A sky130_fd_sc_hd__xnor2_2
XFILLER_109_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12833__A _12853_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07044_ _07041_/X _14304_/Q _07044_/S vssd1 vssd1 vccd1 vccd1 _07045_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13352__A2 _13216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07567__A0 _14098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08995_ _08665_/A _08667_/B _09045_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _09048_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_69_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07946_ _09425_/A vssd1 vssd1 vccd1 vccd1 _08135_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ _07877_/A _07877_/B vssd1 vssd1 vccd1 vccd1 _07877_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_29_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09616_ _09580_/X _09581_/X _09614_/Y _09615_/X vssd1 vssd1 vccd1 vccd1 _09721_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09547_ _09593_/B _09547_/B vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__nor2_1
XFILLER_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09478_ _09478_/A _09478_/B _09478_/C vssd1 vssd1 vccd1 vccd1 _09485_/A sky130_fd_sc_hd__nand3_1
XFILLER_93_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08429_ _13864_/Q vssd1 vssd1 vccd1 vccd1 _09869_/A sky130_fd_sc_hd__buf_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10528__A _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11440_ _11478_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11471_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08598__A2 _09811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _13855_/Q _11377_/B vssd1 vssd1 vccd1 vccd1 _11371_/X sky130_fd_sc_hd__or2_1
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13110_ _13115_/A vssd1 vssd1 vccd1 vccd1 _13110_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10322_ _10374_/A _10374_/B _10374_/C vssd1 vssd1 vccd1 vccd1 _10323_/B sky130_fd_sc_hd__a21oi_1
X_14090_ _14104_/CLK _14090_/D _12738_/Y vssd1 vssd1 vccd1 vccd1 _14090_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041_ _13041_/A vssd1 vssd1 vccd1 vccd1 _13041_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11359__A _14057_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10253_ _10254_/A _10254_/B _10254_/C vssd1 vssd1 vccd1 vccd1 _10255_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07558__A0 _14102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__A1 _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10184_ _10183_/A _10184_/B vssd1 vssd1 vccd1 vccd1 _10184_/X sky130_fd_sc_hd__and2b_1
XANTENNA_input46_A io_wbs_adr[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11106__A1 _11002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13943_ _13943_/CLK _13943_/D _12362_/Y vssd1 vssd1 vccd1 vccd1 _13943_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07325__A3 _07521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14372__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13874_ _13946_/CLK _13874_/D _12276_/Y vssd1 vssd1 vccd1 vccd1 _13874_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12825_ _12210_/X _12900_/B _11745_/Y vssd1 vssd1 vccd1 vccd1 _12825_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07089__A2 _07085_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08286__A1 _08716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12758_/A vssd1 vssd1 vccd1 vccd1 _12756_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08286__B2 _08632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10093__A1 _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ hold6/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__buf_2
XFILLER_37_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _12687_/A vssd1 vssd1 vccd1 vccd1 _14054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14426_ _14427_/CLK _14426_/D vssd1 vssd1 vccd1 vccd1 _14426_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08038__A1 _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11638_ _11638_/A _11548_/X vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__or2b_1
XFILLER_7_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14357_ _14410_/CLK _14357_/D vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_4
X_11569_ _14049_/Q _13961_/Q _11568_/X vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__o21ai_4
X_13308_ _14375_/Q _13307_/X _13294_/X _14455_/Q vssd1 vssd1 vccd1 vccd1 _13308_/X
+ sky130_fd_sc_hd__a22o_1
X_14288_ _14365_/CLK _14288_/D _13151_/Y vssd1 vssd1 vccd1 vccd1 _14288_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13239_ _14328_/Q _13196_/X _13238_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _14328_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09962__A _10000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__A1 _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08210__B2 _08249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07800_ _10931_/A vssd1 vssd1 vccd1 vccd1 _10946_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08780_ _09038_/A _09038_/B _08778_/X _08779_/Y vssd1 vssd1 vccd1 vccd1 _08780_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08578__A _09491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07731_ _07731_/A vssd1 vssd1 vccd1 vccd1 _14070_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07662_ _07662_/A _07665_/A vssd1 vssd1 vccd1 vccd1 _07663_/B sky130_fd_sc_hd__and2_1
XFILLER_37_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09401_ _09401_/A _09401_/B vssd1 vssd1 vccd1 vccd1 _09644_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07593_ _14086_/Q input2/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07594_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09332_ _09329_/Y _09330_/X _09275_/X _09276_/X vssd1 vssd1 vccd1 vccd1 _09345_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_80_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09263_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09263_/X sky130_fd_sc_hd__buf_2
XFILLER_21_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08214_ _08214_/A _08246_/A vssd1 vssd1 vccd1 vccd1 _08247_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09194_ _09140_/X _09194_/B vssd1 vssd1 vccd1 vccd1 _09340_/A sky130_fd_sc_hd__and2b_1
XFILLER_119_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08145_ _08221_/B _08145_/B vssd1 vssd1 vccd1 vccd1 _08195_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12563__A _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10387__A2 _10421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ _08076_/A _08076_/B _08076_/C vssd1 vssd1 vccd1 vccd1 _08081_/B sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_3_4_0_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_84_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07027_ _07027_/A vssd1 vssd1 vccd1 vccd1 _07059_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10083__A _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12533__A0 _12919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13394__A _13411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14395__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08488__A _09865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08978_ _08978_/A _08978_/B _09857_/A _09233_/D vssd1 vssd1 vccd1 vccd1 _08979_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_29_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07929_ _10578_/A vssd1 vssd1 vccd1 vccd1 _10547_/A sky130_fd_sc_hd__buf_2
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10940_ _13899_/Q _13900_/Q _13901_/Q _13902_/Q _10960_/S _10662_/A vssd1 vssd1 vccd1
+ vccd1 _10940_/X sky130_fd_sc_hd__mux4_2
XFILLER_95_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10871_ _13935_/Q _10870_/X _10871_/S vssd1 vssd1 vccd1 vccd1 _10872_/A sky130_fd_sc_hd__mux2_1
X_12610_ input69/X vssd1 vssd1 vccd1 vccd1 _12610_/X sky130_fd_sc_hd__buf_4
XANTENNA_input100_A io_wbs_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12064__A2 _12059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13590_ _13590_/A _13590_/B vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__and2_1
XFILLER_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13261__B2 _14397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12541_ _12924_/A _08716_/A _12555_/S vssd1 vssd1 vccd1 vccd1 _12542_/B sky130_fd_sc_hd__mux2_1
XFILLER_101_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12472_ _08716_/A _12465_/X _12454_/X _14048_/Q vssd1 vssd1 vccd1 vccd1 _12472_/X
+ sky130_fd_sc_hd__a22o_1
X_14211_ _14211_/CLK _14211_/D _13005_/Y vssd1 vssd1 vccd1 vccd1 _14211_/Q sky130_fd_sc_hd__dfrtp_1
X_11423_ _11279_/A _11058_/A _11436_/S vssd1 vssd1 vccd1 vccd1 _11506_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11354_ _11108_/A _11350_/B _11353_/Y _11319_/A _11264_/A vssd1 vssd1 vccd1 vccd1
+ _13895_/D sky130_fd_sc_hd__o32ai_4
X_14142_ _14149_/CLK _14142_/D vssd1 vssd1 vccd1 vccd1 _14142_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10705__B _10705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ _10463_/S _10305_/B vssd1 vssd1 vccd1 vccd1 _10306_/B sky130_fd_sc_hd__xnor2_1
XFILLER_4_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11285_ _11285_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11286_/B sky130_fd_sc_hd__or2_1
X_14073_ _14075_/CLK hold8/X _12717_/Y vssd1 vssd1 vccd1 vccd1 _14073_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12524__A0 _12911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10236_ _10236_/A _10236_/B vssd1 vssd1 vccd1 vccd1 _10236_/Y sky130_fd_sc_hd__nand2_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13024_ _13028_/A vssd1 vssd1 vccd1 vccd1 _13024_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output152_A _14308_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11878__A2 _11872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10167_ _10168_/B _10167_/B vssd1 vssd1 vccd1 vccd1 _10186_/B sky130_fd_sc_hd__xnor2_1
XFILLER_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08398__A _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10098_ _10098_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10099_/A sky130_fd_sc_hd__xnor2_1
XFILLER_94_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13926_ _13927_/CLK _13926_/D _12340_/Y vssd1 vssd1 vccd1 vccd1 _13926_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07703__B1 hold37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13857_ _13988_/CLK _13857_/D _12253_/Y vssd1 vssd1 vccd1 vccd1 _13857_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12808_ _14117_/Q _12800_/X _12807_/X _12805_/X vssd1 vssd1 vccd1 vccd1 _14117_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13788_ _14163_/CLK _13788_/D vssd1 vssd1 vccd1 vccd1 _13788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _12740_/A vssd1 vssd1 vccd1 vccd1 _12739_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11802__A2 _11870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14268__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409_ _14410_/CLK _14409_/D vssd1 vssd1 vccd1 vccd1 _14409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08580__B _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09950_ _09950_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11318__A1 _11119_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08901_ _08921_/A _08902_/B vssd1 vssd1 vccd1 vccd1 _08906_/A sky130_fd_sc_hd__xor2_1
X_09881_ _09881_/A _09881_/B vssd1 vssd1 vccd1 vccd1 _09882_/B sky130_fd_sc_hd__xor2_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08832_ _08861_/B _08861_/C _08861_/A vssd1 vssd1 vccd1 vccd1 _08834_/B sky130_fd_sc_hd__a21bo_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10631__A _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08763_ _08729_/B _08729_/C _08729_/A vssd1 vssd1 vccd1 vccd1 _08764_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__12818__A1 _14121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08101__A _14013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07714_ _14073_/Q _07713_/X _07730_/S vssd1 vssd1 vccd1 vccd1 _07715_/A sky130_fd_sc_hd__mux2_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _09349_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _08745_/B sky130_fd_sc_hd__and2_1
XFILLER_54_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07940__A _14022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07645_ _07662_/A _07665_/A vssd1 vssd1 vccd1 vccd1 _07663_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08755__B _08796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07576_ _14094_/Q input10/X _07582_/S vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09315_ _09236_/B _09236_/C _09236_/A vssd1 vssd1 vccd1 vccd1 _09316_/C sky130_fd_sc_hd__a21bo_1
XFILLER_22_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _09173_/A _09173_/C _09173_/B vssd1 vssd1 vccd1 vccd1 _09248_/B sky130_fd_sc_hd__a21bo_1
X_09177_ _09177_/A _09198_/B _09198_/C vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__and3_1
XFILLER_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12293__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08128_ _08128_/A _08128_/B _10000_/A vssd1 vssd1 vccd1 vccd1 _08130_/A sky130_fd_sc_hd__and3_1
XFILLER_108_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08059_ _13871_/Q vssd1 vssd1 vccd1 vccd1 _09796_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11070_ _11007_/B _11070_/B vssd1 vssd1 vccd1 vccd1 _11071_/B sky130_fd_sc_hd__and2b_1
XFILLER_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10021_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10021_/X sky130_fd_sc_hd__or2_1
XFILLER_27_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08725__A2 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_io_wbs_clk clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14020_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10532__A2 _10524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08011__A _09792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11972_ _11976_/A vssd1 vssd1 vccd1 vccd1 _11972_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08946__A _08946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13711_ input79/X _14457_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13712_/B sky130_fd_sc_hd__mux2_1
X_10923_ _13910_/Q _10922_/X _10923_/S vssd1 vssd1 vccd1 vccd1 _10923_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07161__A1 _14104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13642_ _13642_/A vssd1 vssd1 vccd1 vccd1 _14436_/D sky130_fd_sc_hd__clkbuf_1
X_10854_ _13980_/Q _10895_/B vssd1 vssd1 vccd1 vccd1 _10854_/X sky130_fd_sc_hd__and2_1
XFILLER_73_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _13573_/A _13573_/B vssd1 vssd1 vccd1 vccd1 _13574_/A sky130_fd_sc_hd__and2_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10785_ _13928_/Q _10905_/B vssd1 vssd1 vccd1 vccd1 _10899_/A sky130_fd_sc_hd__nand2_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09777__A _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12524_ _12911_/A _08891_/A _12537_/S vssd1 vssd1 vccd1 vccd1 _12525_/B sky130_fd_sc_hd__mux2_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08661__B2 _08925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12455_ _08896_/A _12439_/X _12454_/X _14044_/Q vssd1 vssd1 vccd1 vccd1 _12455_/X
+ sky130_fd_sc_hd__a22o_1
X_11406_ _13877_/Q _11392_/A _11396_/X _11405_/X vssd1 vssd1 vccd1 vccd1 _13877_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_74_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14152_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12386_ _12410_/A vssd1 vssd1 vccd1 vccd1 _12391_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_114_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10435__B _10435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14125_ _14239_/CLK _14125_/D vssd1 vssd1 vccd1 vccd1 _14125_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11337_ _10826_/A _11333_/C _11336_/Y _10851_/B _11282_/A vssd1 vssd1 vccd1 vccd1
+ _13901_/D sky130_fd_sc_hd__a32o_1
XFILLER_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14056_ _14411_/CLK _14056_/D vssd1 vssd1 vccd1 vccd1 _14056_/Q sky130_fd_sc_hd__dfxtp_2
X_11268_ _11268_/A _11268_/B _11268_/C vssd1 vssd1 vccd1 vccd1 _11350_/B sky130_fd_sc_hd__and3_1
XFILLER_97_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _13009_/A vssd1 vssd1 vccd1 vccd1 _13007_/Y sky130_fd_sc_hd__inv_2
X_10219_ _10220_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10219_/Y sky130_fd_sc_hd__nand2_1
X_11199_ _10652_/A _11147_/X _11143_/X vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__o21a_1
XFILLER_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13909_ _13949_/CLK _13909_/D _12319_/Y vssd1 vssd1 vccd1 vccd1 _13909_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_62_io_wbs_clk_A clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_78_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07430_ _14203_/Q _14205_/Q _07442_/S vssd1 vssd1 vccd1 vccd1 _07431_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12097__B _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07361_ _07349_/X _07359_/X _07360_/X _07352_/X vssd1 vssd1 vccd1 vccd1 _07361_/X
+ sky130_fd_sc_hd__a22o_1
X_09100_ _09100_/A _09100_/B _09100_/C vssd1 vssd1 vccd1 vccd1 _09144_/B sky130_fd_sc_hd__nand3_4
XANTENNA__13701__S _13704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07292_ _14241_/Q _14228_/Q _07506_/S vssd1 vssd1 vccd1 vccd1 _07293_/A sky130_fd_sc_hd__mux2_1
X_09031_ _09029_/B _09029_/C _09029_/A vssd1 vssd1 vccd1 vccd1 _09031_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_102_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06966__A1 _14314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09933_ _09978_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09934_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07935__A _13870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__A1 _08547_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09864_ _09892_/A vssd1 vssd1 vccd1 vccd1 _10126_/B sky130_fd_sc_hd__clkbuf_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08815_ _09188_/A _08815_/B _08815_/C vssd1 vssd1 vccd1 vccd1 _08815_/X sky130_fd_sc_hd__and3_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09795_ _13871_/Q _09817_/A vssd1 vssd1 vccd1 vccd1 _09824_/B sky130_fd_sc_hd__xor2_4
XFILLER_39_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08746_ _09200_/B vssd1 vssd1 vccd1 vccd1 _09887_/A sky130_fd_sc_hd__buf_4
XFILLER_96_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _08675_/Y _08674_/X _08620_/X _08618_/X vssd1 vssd1 vccd1 vccd1 _08678_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _14127_/Q _14062_/Q vssd1 vssd1 vccd1 vccd1 _07628_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ _07559_/A vssd1 vssd1 vccd1 vccd1 _14102_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11920__A _11920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10570_ _10587_/A _10327_/X _10375_/X vssd1 vssd1 vccd1 vccd1 _10583_/B sky130_fd_sc_hd__o21ba_1
XFILLER_22_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09229_ _09277_/A _09277_/B _09277_/C vssd1 vssd1 vccd1 vccd1 _09229_/X sky130_fd_sc_hd__and3_1
X_12240_ _12252_/A vssd1 vssd1 vccd1 vccd1 _12245_/A sky130_fd_sc_hd__buf_2
XANTENNA__08006__A _14019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ _13829_/Q _12095_/A _12170_/X _12161_/X vssd1 vssd1 vccd1 vccd1 _13829_/D
+ sky130_fd_sc_hd__o211a_1
X_11122_ _11122_/A _11122_/B _11125_/B vssd1 vssd1 vccd1 vccd1 _11122_/X sky130_fd_sc_hd__or3_1
XANTENNA__07845__A _14031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11053_ _11127_/B _11127_/C _11127_/A vssd1 vssd1 vccd1 vccd1 _11124_/C sky130_fd_sc_hd__a21oi_1
XFILLER_77_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10004_ _10004_/A _10004_/B vssd1 vssd1 vccd1 vccd1 _10382_/B sky130_fd_sc_hd__xnor2_2
XFILLER_88_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_io_wbs_clk clkbuf_2_3_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_io_wbs_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_92_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11955_ _11959_/A vssd1 vssd1 vccd1 vccd1 _11955_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output115_A _11832_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10906_ _10906_/A vssd1 vssd1 vccd1 vccd1 _11125_/A sky130_fd_sc_hd__buf_4
XFILLER_83_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11886_ _13810_/Q _11882_/X _11883_/X _11884_/Y _11885_/X vssd1 vssd1 vccd1 vccd1
+ _13750_/D sky130_fd_sc_hd__o221a_1
XFILLER_44_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13625_ _13625_/A _13625_/B vssd1 vssd1 vccd1 vccd1 _13626_/A sky130_fd_sc_hd__and2_1
XFILLER_16_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10837_ _10902_/S vssd1 vssd1 vccd1 vccd1 _10871_/S sky130_fd_sc_hd__buf_2
XANTENNA__12926__A _12926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13556_ _13556_/A _13556_/B vssd1 vssd1 vccd1 vccd1 _13557_/A sky130_fd_sc_hd__and2_1
XFILLER_73_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10768_ _10768_/A _10768_/B _13932_/Q vssd1 vssd1 vccd1 vccd1 _10879_/B sky130_fd_sc_hd__or3b_1
XFILLER_40_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12507_ _13358_/A _13111_/C vssd1 vssd1 vccd1 vccd1 _12567_/B sky130_fd_sc_hd__nand2_1
XFILLER_73_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13487_ _13504_/A vssd1 vssd1 vccd1 vccd1 _13502_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10699_ _11220_/A vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__clkbuf_2
X_12438_ _12485_/A vssd1 vssd1 vccd1 vccd1 _12438_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13391__A0 _12664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12369_ _12372_/A vssd1 vssd1 vccd1 vccd1 _12369_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06948__A1 _14284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14306__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14108_ _14239_/CLK _14108_/D vssd1 vssd1 vccd1 vccd1 _14108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06930_ _14462_/Q _14286_/Q vssd1 vssd1 vccd1 vccd1 _06930_/Y sky130_fd_sc_hd__nand2_1
X_14039_ _14054_/CLK _14039_/D vssd1 vssd1 vccd1 vccd1 _14039_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06861_ _13780_/Q vssd1 vssd1 vccd1 vccd1 _11659_/A sky130_fd_sc_hd__clkinv_2
XFILLER_41_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08600_ _08600_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08670_/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09580_ _09673_/A _09580_/B vssd1 vssd1 vccd1 vccd1 _09580_/X sky130_fd_sc_hd__or2_1
XFILLER_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08531_ _08532_/A _08531_/B _08531_/C vssd1 vssd1 vccd1 vccd1 _08719_/A sky130_fd_sc_hd__nand3_1
XANTENNA__07921__C _07921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08462_ _09811_/A vssd1 vssd1 vccd1 vccd1 _08703_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_91_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07413_ _14091_/Q _07404_/X _07406_/X _13891_/Q _07521_/B vssd1 vssd1 vccd1 vccd1
+ _07413_/X sky130_fd_sc_hd__a221o_1
X_08393_ _09698_/A _08390_/Y _08391_/X _08392_/Y vssd1 vssd1 vccd1 vccd1 _09729_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07344_ _14219_/Q _14221_/Q _07360_/S vssd1 vssd1 vccd1 vccd1 _07344_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07275_ _14189_/Q _14188_/Q _14187_/Q vssd1 vssd1 vccd1 vccd1 _07276_/B sky130_fd_sc_hd__or3_1
X_09014_ _09014_/A _09014_/B vssd1 vssd1 vccd1 vccd1 _09015_/B sky130_fd_sc_hd__nor2_1
XFILLER_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13382__A0 _12650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09916_ _10197_/A _09940_/B _09915_/X vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__10091__A _10091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _09848_/A _09848_/B vssd1 vssd1 vccd1 vccd1 _09847_/X sky130_fd_sc_hd__and2_2
XFILLER_101_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09778_ _09778_/A _09778_/B vssd1 vssd1 vccd1 vccd1 _09779_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _08729_/A _08729_/B _08729_/C vssd1 vssd1 vccd1 vccd1 _08764_/A sky130_fd_sc_hd__and3_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _13764_/Q _11740_/B vssd1 vssd1 vccd1 vccd1 _11740_/Y sky130_fd_sc_hd__nor2_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _13779_/Q _11675_/A _11682_/C _13780_/Q vssd1 vssd1 vccd1 vccd1 _11672_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13410_ _13410_/A vssd1 vssd1 vccd1 vccd1 _14370_/D sky130_fd_sc_hd__clkbuf_1
X_10622_ _10622_/A _10622_/B vssd1 vssd1 vccd1 vccd1 _10622_/Y sky130_fd_sc_hd__nor2_1
X_14390_ _14450_/CLK _14390_/D vssd1 vssd1 vccd1 vccd1 _14390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08662__C _09482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ _13341_/A vssd1 vssd1 vccd1 vccd1 _13341_/X sky130_fd_sc_hd__clkbuf_2
X_10553_ _10564_/A _10564_/B _10564_/C vssd1 vssd1 vccd1 vccd1 _10565_/C sky130_fd_sc_hd__a21o_1
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input76_A io_wbs_datwr[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ _14367_/Q _13208_/X _13271_/X _13258_/X vssd1 vssd1 vccd1 vccd1 _13272_/X
+ sky130_fd_sc_hd__a211o_1
X_10484_ _10470_/B _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10495_/A sky130_fd_sc_hd__mux2_1
X_12223_ _12223_/A vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__buf_6
XFILLER_29_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12154_ _12906_/A _12160_/B vssd1 vssd1 vccd1 vccd1 _12154_/X sky130_fd_sc_hd__or2_1
XFILLER_68_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11105_ _11108_/A _11105_/B vssd1 vssd1 vccd1 vccd1 _11105_/Y sky130_fd_sc_hd__nor2_1
X_12085_ _12517_/A _12085_/B vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__and2_1
XFILLER_1_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11036_ _11052_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11124_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07107__A1 _07090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12987_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12987_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11938_ _11940_/A vssd1 vssd1 vccd1 vccd1 _11938_/Y sky130_fd_sc_hd__inv_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10875__S _10875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ _11869_/A vssd1 vssd1 vccd1 vccd1 _11869_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13608_ _13608_/A vssd1 vssd1 vccd1 vccd1 _14427_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13061__C1 _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13539_ _13539_/A _13539_/B vssd1 vssd1 vccd1 vccd1 _13540_/A sky130_fd_sc_hd__and2_1
XFILLER_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09280__A1 _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09280__B2 _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07060_ _07051_/X _07059_/X _14366_/Q vssd1 vssd1 vccd1 vccd1 _07061_/S sky130_fd_sc_hd__o21a_1
XANTENNA__08291__D _09233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13487__A _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10904__A _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07962_ _09803_/B vssd1 vssd1 vccd1 vccd1 _08983_/C sky130_fd_sc_hd__buf_2
X_09701_ _09698_/X _09699_/Y _09687_/A _09687_/Y vssd1 vssd1 vccd1 vccd1 _09727_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_96_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06913_ _06909_/X _14321_/Q _06913_/S vssd1 vssd1 vccd1 vccd1 _06914_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11678__B1 _13778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ _07893_/A _07893_/B vssd1 vssd1 vccd1 vccd1 _07893_/Y sky130_fd_sc_hd__xnor2_1
X_09632_ _09527_/A _09527_/C _09527_/B vssd1 vssd1 vccd1 vccd1 _09632_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09563_ _09563_/A _09563_/B _09563_/C vssd1 vssd1 vccd1 vccd1 _09592_/B sky130_fd_sc_hd__nand3_2
XFILLER_71_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08514_ _08693_/B _08693_/C _08693_/A vssd1 vssd1 vccd1 vccd1 _08517_/B sky130_fd_sc_hd__o21bai_1
XFILLER_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09494_ _09491_/Y _09494_/B _09541_/A vssd1 vssd1 vccd1 vccd1 _09541_/B sky130_fd_sc_hd__nand3b_1
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08445_ _08750_/A vssd1 vssd1 vccd1 vccd1 _08445_/X sky130_fd_sc_hd__buf_4
XFILLER_93_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09859__B _10090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08376_ _08376_/A _08376_/B vssd1 vssd1 vccd1 vccd1 _08384_/B sky130_fd_sc_hd__and2_1
XFILLER_17_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07327_ _14106_/Q _07323_/X vssd1 vssd1 vccd1 vccd1 _07327_/X sky130_fd_sc_hd__or2b_1
XFILLER_20_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09875__A _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07258_ _14076_/Q _13876_/Q _07258_/S vssd1 vssd1 vccd1 vccd1 _07258_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12158__A1 _13825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07189_ _14281_/Q _07187_/X _07201_/S vssd1 vssd1 vccd1 vccd1 _07190_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07395__A _14093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11133__A2 _11110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12910_ _14151_/Q _12901_/X _12909_/X _12907_/X vssd1 vssd1 vccd1 vccd1 _14151_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13890_ _14107_/CLK _13890_/D _12296_/Y vssd1 vssd1 vccd1 vccd1 _13890_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12841_ _12847_/A _12841_/B vssd1 vssd1 vccd1 vccd1 _12842_/A sky130_fd_sc_hd__and2_1
XFILLER_46_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12772_ _12801_/A vssd1 vssd1 vccd1 vccd1 _12772_/X sky130_fd_sc_hd__buf_2
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11882_/A vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__buf_2
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09769__B _09769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14442_ _14442_/CLK _14442_/D vssd1 vssd1 vccd1 vccd1 _14442_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _14040_/Q _13952_/Q vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__or2_1
XFILLER_70_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10605_ _09421_/C _10604_/Y _10597_/A vssd1 vssd1 vccd1 vccd1 _10605_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_11_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14373_ _14453_/CLK _14373_/D vssd1 vssd1 vccd1 vccd1 _14373_/Q sky130_fd_sc_hd__dfxtp_1
X_11585_ _13857_/Q _11584_/Y _11585_/S vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13324_ _14379_/Q _13307_/X _13315_/X _14459_/Q vssd1 vssd1 vccd1 vccd1 _13324_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07273__B1 _14166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10536_ _10546_/B _10546_/C _10546_/A vssd1 vssd1 vccd1 vccd1 _10548_/C sky130_fd_sc_hd__a21o_1
XFILLER_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12149__A1 _13822_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13255_ _14331_/Q _13240_/X _13253_/X _13254_/X vssd1 vssd1 vccd1 vccd1 _14331_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _10467_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _10468_/B sky130_fd_sc_hd__or2_1
X_12206_ _13837_/Q _12201_/A _12202_/C vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__a21bo_1
X_13186_ _13189_/A vssd1 vssd1 vccd1 vccd1 _13186_/Y sky130_fd_sc_hd__inv_2
X_10398_ _10383_/A _10396_/Y _10397_/X vssd1 vssd1 vccd1 vccd1 _10399_/B sky130_fd_sc_hd__a21oi_4
XFILLER_96_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ input76/X _12143_/B vssd1 vssd1 vccd1 vccd1 _12137_/X sky130_fd_sc_hd__or2_1
XFILLER_36_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12068_ _13801_/Q _12059_/X _12060_/X _13817_/Q vssd1 vssd1 vccd1 vccd1 _12069_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11019_ _13917_/Q vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11832__B1 _11823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12386__A _12410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08230_ _09673_/A vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08161_ _08389_/A vssd1 vssd1 vccd1 vccd1 _09685_/A sky130_fd_sc_hd__buf_2
XFILLER_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07112_ _14263_/Q _07085_/X _07111_/X _14359_/Q vssd1 vssd1 vccd1 vccd1 _07112_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09695__A _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08092_ _14009_/Q _09821_/A vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__nand2_4
X_07043_ _07012_/X _07042_/X _14368_/Q vssd1 vssd1 vccd1 vccd1 _07044_/S sky130_fd_sc_hd__o21a_1
XANTENNA__10634__A _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13010__A _13010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08104__A _08789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07567__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08994_ _08993_/B _08993_/C _08993_/A vssd1 vssd1 vccd1 vccd1 _08994_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07943__A _09818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _14021_/Q vssd1 vssd1 vccd1 vccd1 _09425_/A sky130_fd_sc_hd__buf_2
XFILLER_68_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07876_ _07876_/A _07876_/B vssd1 vssd1 vccd1 vccd1 _07877_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09615_ _09611_/X _09613_/Y _09573_/B _09573_/Y vssd1 vssd1 vccd1 vccd1 _09615_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13680__A _13680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09546_ _09545_/C _08070_/C _09593_/A _09544_/Y vssd1 vssd1 vccd1 vccd1 _09547_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09477_ _09427_/B _09427_/C _09427_/A vssd1 vssd1 vccd1 vccd1 _09478_/C sky130_fd_sc_hd__o21bai_1
XFILLER_34_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09492__B2 _09443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08428_ _09881_/B vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13576__A0 _12561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08047__A2 _09800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ _09479_/A _09479_/B _09796_/A _09123_/C vssd1 vssd1 vccd1 vccd1 _08360_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07255__A0 _14077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ _11396_/A vssd1 vssd1 vccd1 vccd1 _11370_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10321_ _10374_/A _10374_/B _10374_/C vssd1 vssd1 vccd1 vccd1 _10323_/A sky130_fd_sc_hd__and3_1
XFILLER_106_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13040_ _13032_/X _13036_/X _13038_/X _13039_/X vssd1 vssd1 vccd1 vccd1 _14232_/D
+ sky130_fd_sc_hd__o211a_1
X_10252_ _10421_/B _10252_/B vssd1 vssd1 vccd1 vccd1 _10254_/C sky130_fd_sc_hd__xnor2_1
XFILLER_79_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07558__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10183_ _10183_/A _10184_/B vssd1 vssd1 vccd1 vccd1 _10225_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07853__A _14035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input39_A io_wbs_adr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13942_ _13943_/CLK _13942_/D _12360_/Y vssd1 vssd1 vccd1 vccd1 _13942_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10865__A1 _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13873_ _13946_/CLK _13873_/D _12275_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12824_ _12902_/B vssd1 vssd1 vccd1 vccd1 _12900_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11814__B1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _12758_/A vssd1 vssd1 vccd1 vccd1 _12755_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_67_io_wbs_clk_A clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08286__A2 _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11706_ _11730_/B _11882_/A vssd1 vssd1 vccd1 vccd1 _11706_/Y sky130_fd_sc_hd__nor2_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12686_ _12696_/A _12686_/B vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__and2_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _14427_/CLK _14425_/D vssd1 vssd1 vccd1 vccd1 _14425_/Q sky130_fd_sc_hd__dfxtp_1
X_11637_ _11585_/S _11634_/X _11635_/Y _11636_/X vssd1 vssd1 vccd1 vccd1 _13845_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09235__A1 _09233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__A _13254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09235__B2 _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__A0 _14080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14356_ _14365_/CLK _14356_/D vssd1 vssd1 vccd1 vccd1 _14356_/Q sky130_fd_sc_hd__dfxtp_2
X_11568_ _14049_/Q _13961_/Q _11619_/A vssd1 vssd1 vccd1 vccd1 _11568_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12790__A1 _14154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13307_ _13328_/A vssd1 vssd1 vccd1 vccd1 _13307_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10519_ _07924_/X _10511_/X _10516_/Y _10518_/X vssd1 vssd1 vccd1 vccd1 _13968_/D
+ sky130_fd_sc_hd__o31a_1
X_14287_ _14365_/CLK _14287_/D _13150_/Y vssd1 vssd1 vccd1 vccd1 _14287_/Q sky130_fd_sc_hd__dfrtp_4
X_11499_ _11499_/A vssd1 vssd1 vccd1 vccd1 _11499_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13238_ _14408_/Q _13199_/X _13235_/X _13237_/X vssd1 vssd1 vccd1 vccd1 _13238_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10173__B _10173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13169_ _13171_/A vssd1 vssd1 vccd1 vccd1 _13169_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08210__A2 _09800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__B _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07730_ _14070_/Q _07729_/X _07730_/S vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07661_ _14143_/Q _07727_/A vssd1 vssd1 vccd1 vccd1 _07661_/X sky130_fd_sc_hd__or2_1
XFILLER_26_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13704__S _13704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09400_ _09999_/B _08091_/A _09319_/A _09317_/Y vssd1 vssd1 vccd1 vccd1 _09401_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07592_ _07592_/A vssd1 vssd1 vccd1 vccd1 _14087_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ _09275_/X _09276_/X _09329_/Y _09330_/X vssd1 vssd1 vccd1 vccd1 _09345_/A
+ sky130_fd_sc_hd__a211o_2
XANTENNA__11805__B1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09262_ _09191_/Y _09192_/Y _09263_/A _09261_/Y vssd1 vssd1 vccd1 vccd1 _09262_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08213_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08246_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09193_ _09402_/A vssd1 vssd1 vccd1 vccd1 _09629_/A sky130_fd_sc_hd__buf_4
X_08144_ _08144_/A _08144_/B _08144_/C vssd1 vssd1 vccd1 vccd1 _08145_/B sky130_fd_sc_hd__or3_1
XFILLER_119_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08985__B1 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08075_ _08076_/B _08076_/C _08076_/A vssd1 vssd1 vccd1 vccd1 _08081_/A sky130_fd_sc_hd__a21o_1
XFILLER_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07026_ _14274_/Q _07007_/X _07025_/X _14370_/Q vssd1 vssd1 vccd1 vccd1 _07026_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12533__A1 _08983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13927_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_103_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_103_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_08977_ _08468_/B _09857_/A _09482_/B _08925_/A vssd1 vssd1 vccd1 vccd1 _08979_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07928_ _08249_/A vssd1 vssd1 vccd1 vccd1 _10578_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07859_ _07868_/B _07857_/Y _07858_/Y vssd1 vssd1 vccd1 vccd1 _07859_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10870_ _13977_/Q _10869_/Y _10875_/S vssd1 vssd1 vccd1 vccd1 _10870_/X sky130_fd_sc_hd__mux2_1
XFILLER_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11642__B _13955_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09529_ _09516_/A _09516_/B _09528_/X vssd1 vssd1 vccd1 vccd1 _09580_/B sky130_fd_sc_hd__a21oi_2
XFILLER_25_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ _12562_/S vssd1 vssd1 vccd1 vccd1 _12555_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_52_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13549__A0 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12471_ _13996_/Q _12460_/X _12470_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _13996_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14210_ _14217_/CLK _14210_/D _13003_/Y vssd1 vssd1 vccd1 vccd1 _14210_/Q sky130_fd_sc_hd__dfrtp_1
X_11422_ _11425_/S vssd1 vssd1 vccd1 vccd1 _11436_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_64_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14365_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_14141_ _14149_/CLK _14141_/D vssd1 vssd1 vccd1 vccd1 _14141_/Q sky130_fd_sc_hd__dfxtp_2
X_11353_ _11268_/A _11268_/B _11268_/C vssd1 vssd1 vccd1 vccd1 _11353_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06987__C1 hold33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ _10333_/A _10333_/B vssd1 vssd1 vccd1 vccd1 _10306_/A sky130_fd_sc_hd__xor2_1
X_14072_ _14075_/CLK _14072_/D _12715_/Y vssd1 vssd1 vccd1 vccd1 _14072_/Q sky130_fd_sc_hd__dfrtp_1
X_11284_ _11336_/B _11336_/C _11336_/A vssd1 vssd1 vccd1 vccd1 _11333_/C sky130_fd_sc_hd__a21o_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13721__A0 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12524__A1 _08891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13023_ _13116_/A vssd1 vssd1 vccd1 vccd1 _13028_/A sky130_fd_sc_hd__buf_2
XFILLER_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10235_ _10236_/A _10236_/B _10231_/Y _10233_/Y vssd1 vssd1 vccd1 vccd1 _10235_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08679__A _08980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ _10166_/A _10166_/B vssd1 vssd1 vccd1 vccd1 _10167_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output145_A _14301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10097_ _10086_/X _10139_/B _10096_/X vssd1 vssd1 vccd1 vccd1 _10100_/A sky130_fd_sc_hd__a21o_1
XFILLER_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13925_ _13927_/CLK _13925_/D _12339_/Y vssd1 vssd1 vccd1 vccd1 _13925_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__07703__A1 _14148_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13856_ _13988_/CLK _13856_/D _12251_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12807_ _14158_/Q _12801_/X _12803_/X _14142_/Q _12791_/X vssd1 vssd1 vccd1 vccd1
+ _12807_/X sky130_fd_sc_hd__a221o_2
XANTENNA__11552__B _13953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13787_ _13809_/CLK _13787_/D vssd1 vssd1 vccd1 vccd1 _13787_/Q sky130_fd_sc_hd__dfxtp_1
X_10999_ _11220_/A _10999_/B vssd1 vssd1 vccd1 vccd1 _11000_/B sky130_fd_sc_hd__nor2_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12740_/A vssd1 vssd1 vccd1 vccd1 _12738_/Y sky130_fd_sc_hd__inv_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09208__A1 _08623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12669_ _12669_/A vssd1 vssd1 vccd1 vccd1 _12685_/S sky130_fd_sc_hd__buf_2
XANTENNA__09208__B2 _08623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07219__A0 _14272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14408_ _14411_/CLK _14408_/D vssd1 vssd1 vccd1 vccd1 _14408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14339_ _14400_/CLK _14339_/D vssd1 vssd1 vccd1 vccd1 _14339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09973__A _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08900_ _08937_/B _10061_/A _08866_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08902_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09880_ _09880_/A _09880_/B vssd1 vssd1 vccd1 vccd1 _09986_/A sky130_fd_sc_hd__xnor2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10526__B1 _10562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__A _10912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08831_/A _08869_/A _08831_/C vssd1 vssd1 vccd1 vccd1 _08861_/A sky130_fd_sc_hd__nand3_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08762_/A _08774_/B _08762_/C vssd1 vssd1 vccd1 vccd1 _08805_/C sky130_fd_sc_hd__or3_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07713_ _07700_/B hold7/X _07723_/A vssd1 vssd1 vccd1 vccd1 _07713_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08693_ _08693_/A _08693_/B _08693_/C vssd1 vssd1 vccd1 vccd1 _08701_/A sky130_fd_sc_hd__or3_1
XFILLER_39_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07644_ _14068_/Q _07664_/B vssd1 vssd1 vccd1 vccd1 _07665_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07575_ _07575_/A vssd1 vssd1 vccd1 vccd1 _14095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09314_ _08867_/A _09822_/A _09313_/A _09313_/C vssd1 vssd1 vccd1 vccd1 _09316_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08474__D _13859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09245_ _09245_/A _09245_/B _09245_/C vssd1 vssd1 vccd1 vccd1 _09248_/A sky130_fd_sc_hd__nand3_2
XFILLER_90_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09176_ _09198_/A _09198_/C _09198_/B vssd1 vssd1 vccd1 vccd1 _09176_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11557__A2 _13955_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08127_ _09508_/C vssd1 vssd1 vccd1 vccd1 _10000_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08058_ _09472_/A _09472_/B _09543_/D _09493_/D vssd1 vssd1 vccd1 vccd1 _08140_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07009_ _07087_/A vssd1 vssd1 vccd1 vccd1 _07009_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10020_ _10092_/B _10191_/B vssd1 vssd1 vccd1 vccd1 _10054_/B sky130_fd_sc_hd__xnor2_2
XFILLER_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10532__A3 _10530_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11971_ _11971_/A vssd1 vssd1 vccd1 vccd1 _11976_/A sky130_fd_sc_hd__buf_2
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08946__B _10206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ _13710_/A vssd1 vssd1 vccd1 vccd1 _14456_/D sky130_fd_sc_hd__clkbuf_1
X_10922_ _13908_/Q _13909_/Q _10931_/A vssd1 vssd1 vccd1 vccd1 _10922_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13641_ _13644_/A _13641_/B vssd1 vssd1 vccd1 vccd1 _13642_/A sky130_fd_sc_hd__and2_1
XFILLER_60_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10853_ _10853_/A _10853_/B _10853_/C vssd1 vssd1 vccd1 vccd1 _10853_/X sky130_fd_sc_hd__or3_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _12681_/X _14417_/Q _13576_/S vssd1 vssd1 vccd1 vccd1 _13573_/B sky130_fd_sc_hd__mux2_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _13929_/Q _10786_/B vssd1 vssd1 vccd1 vccd1 _10894_/A sky130_fd_sc_hd__nand2_1
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12562_/S vssd1 vssd1 vccd1 vccd1 _12537_/S sky130_fd_sc_hd__clkbuf_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09777__B _09777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08661__A2 _09482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12454_ _12476_/A vssd1 vssd1 vccd1 vccd1 _12454_/X sky130_fd_sc_hd__clkbuf_2
X_11405_ _13841_/Q _11407_/B vssd1 vssd1 vccd1 vccd1 _11405_/X sky130_fd_sc_hd__or2_1
X_12385_ _12385_/A vssd1 vssd1 vccd1 vccd1 _12410_/A sky130_fd_sc_hd__clkbuf_2
X_14124_ _14239_/CLK _14124_/D vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__09793__A _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11336_ _11336_/A _11336_/B _11336_/C vssd1 vssd1 vccd1 vccd1 _11336_/Y sky130_fd_sc_hd__nand3_1
XFILLER_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14055_ _14363_/CLK _14055_/D vssd1 vssd1 vccd1 vccd1 _14055_/Q sky130_fd_sc_hd__dfxtp_2
X_11267_ _11355_/B _11355_/A vssd1 vssd1 vccd1 vccd1 _11268_/C sky130_fd_sc_hd__and2b_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13006_ _13009_/A vssd1 vssd1 vccd1 vccd1 _13006_/Y sky130_fd_sc_hd__inv_2
X_10218_ _10067_/A _10216_/X _10217_/X vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__a21oi_1
XFILLER_97_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11198_ _11220_/B _11221_/A vssd1 vssd1 vccd1 vccd1 _11216_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10149_ _10149_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10150_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09126__B1 _09218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12659__A _13072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11484__A1 _11002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13908_ _13949_/CLK _13908_/D _12318_/Y vssd1 vssd1 vccd1 vccd1 _13908_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11282__B _11282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ _14259_/CLK _13839_/D vssd1 vssd1 vccd1 vccd1 _13839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13225__A2 _13336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07360_ _14216_/Q _14218_/Q _07360_/S vssd1 vssd1 vccd1 vccd1 _07360_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07291_ _07521_/D vssd1 vssd1 vccd1 vccd1 _07506_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09030_ _09030_/A vssd1 vssd1 vccd1 vccd1 _09030_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07000__B _14277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09932_ _10195_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__and2b_1
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09863_ _09863_/A _09875_/B vssd1 vssd1 vccd1 vccd1 _09892_/A sky130_fd_sc_hd__xnor2_4
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _08809_/B _08814_/B vssd1 vssd1 vccd1 vccd1 _08814_/X sky130_fd_sc_hd__and2b_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _10279_/A vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__buf_4
XFILLER_61_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07951__A _09362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08745_ _08745_/A _08745_/B _08745_/C vssd1 vssd1 vccd1 vccd1 _08758_/A sky130_fd_sc_hd__nand3_1
XFILLER_100_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08676_ _08618_/X _08620_/X _08674_/X _08675_/Y vssd1 vssd1 vccd1 vccd1 _08678_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07162__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _14128_/Q _14063_/Q vssd1 vssd1 vccd1 vccd1 _07675_/A sky130_fd_sc_hd__or2_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07558_ _14102_/Q input19/X _07560_/S vssd1 vssd1 vccd1 vccd1 _07559_/A sky130_fd_sc_hd__mux2_1
XANTENNA__08782__A _09943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07489_ _07277_/C _07329_/X _07399_/A vssd1 vssd1 vccd1 vccd1 _07489_/X sky130_fd_sc_hd__a21bo_1
XFILLER_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09228_ _09215_/A _09215_/B _09215_/C vssd1 vssd1 vccd1 vccd1 _09277_/C sky130_fd_sc_hd__a21o_1
XFILLER_10_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09159_ _09158_/A _09158_/C _09158_/B vssd1 vssd1 vccd1 vccd1 _09161_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ _12919_/A _12173_/B vssd1 vssd1 vccd1 vccd1 _12170_/X sky130_fd_sc_hd__or2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11121_ _11119_/X _11117_/C _11120_/Y _11100_/X _11058_/A vssd1 vssd1 vccd1 vccd1
+ _13917_/D sky130_fd_sc_hd__a32o_1
XFILLER_107_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11052_ _11052_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11127_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10271__B _10271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _10003_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _10030_/A sky130_fd_sc_hd__xnor2_2
XFILLER_40_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input21_A dout1[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07861__A _14039_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12479__A _12817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11954_ _11971_/A vssd1 vssd1 vccd1 vccd1 _11959_/A sky130_fd_sc_hd__buf_2
XFILLER_44_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10905_ _13928_/Q _10905_/B vssd1 vssd1 vccd1 vccd1 _10905_/X sky130_fd_sc_hd__or2_1
XFILLER_45_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11885_ _11920_/A vssd1 vssd1 vccd1 vccd1 _11885_/X sky130_fd_sc_hd__clkbuf_2
X_13624_ input86/X _14432_/Q _13628_/S vssd1 vssd1 vccd1 vccd1 _13625_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09788__A _09788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10836_ _13983_/Q _10835_/Y _10836_/S vssd1 vssd1 vccd1 vccd1 _10836_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13555_ _12660_/X _14412_/Q _13559_/S vssd1 vssd1 vccd1 vccd1 _13556_/B sky130_fd_sc_hd__mux2_1
X_10767_ _11020_/A _10767_/B vssd1 vssd1 vccd1 vccd1 _10768_/A sky130_fd_sc_hd__xnor2_1
XFILLER_9_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09831__A1 _10435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12506_ _14006_/Q _12460_/A _12505_/X _12498_/X vssd1 vssd1 vccd1 vccd1 _14006_/D
+ sky130_fd_sc_hd__o211a_1
X_13486_ _13486_/A vssd1 vssd1 vccd1 vccd1 _14392_/D sky130_fd_sc_hd__clkbuf_1
X_10698_ _11228_/A vssd1 vssd1 vccd1 vccd1 _11220_/A sky130_fd_sc_hd__clkbuf_2
X_12437_ _13989_/Q _12422_/X _12436_/X _12203_/X vssd1 vssd1 vccd1 vccd1 _13989_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12942__A _12942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13391__A1 _14365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12368_ _12372_/A vssd1 vssd1 vccd1 vccd1 _12368_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14107_ _14107_/CLK _14107_/D _12758_/Y vssd1 vssd1 vccd1 vccd1 _14107_/Q sky130_fd_sc_hd__dfrtp_4
X_11319_ _11319_/A vssd1 vssd1 vccd1 vccd1 _11319_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12299_ _12317_/A vssd1 vssd1 vccd1 vccd1 _12304_/A sky130_fd_sc_hd__buf_4
XFILLER_113_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14038_ _14054_/CLK _14038_/D vssd1 vssd1 vccd1 vccd1 _14038_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11154__A0 _11032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06860_ _14396_/Q _13775_/Q vssd1 vssd1 vccd1 vccd1 _06869_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08867__A _08867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08530_ _08530_/A _08530_/B vssd1 vssd1 vccd1 vccd1 _08531_/C sky130_fd_sc_hd__xnor2_1
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08461_ _09165_/C vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__buf_2
XFILLER_36_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07412_ _07431_/A _07412_/B vssd1 vssd1 vccd1 vccd1 _07412_/X sky130_fd_sc_hd__or2_1
X_08392_ _08391_/A _08391_/B _08391_/C vssd1 vssd1 vccd1 vccd1 _08392_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07343_ _14103_/Q _07336_/X vssd1 vssd1 vccd1 vccd1 _07343_/X sky130_fd_sc_hd__or2b_1
XFILLER_52_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07274_ _07274_/A vssd1 vssd1 vccd1 vccd1 _07300_/B sky130_fd_sc_hd__inv_2
XANTENNA__08107__A _14013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09013_ _08573_/B _08494_/D _09942_/A _08012_/A vssd1 vssd1 vccd1 vccd1 _09014_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_89_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07946__A _09425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07061__A1 _14302_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09915_ _09912_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _09915_/X sky130_fd_sc_hd__and2b_1
XFILLER_63_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09846_ _10126_/A vssd1 vssd1 vccd1 vccd1 _10205_/A sky130_fd_sc_hd__clkbuf_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07681__A _14125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09778_/B sky130_fd_sc_hd__xor2_1
XFILLER_74_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06989_ _14405_/Q _07020_/B _14437_/Q vssd1 vssd1 vccd1 vccd1 _06989_/X sky130_fd_sc_hd__and3b_1
XANTENNA__12299__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08728_ _08723_/B _08723_/C _08723_/A vssd1 vssd1 vccd1 vccd1 _08729_/C sky130_fd_sc_hd__a21o_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08659_ _13870_/Q vssd1 vssd1 vccd1 vccd1 _09818_/A sky130_fd_sc_hd__buf_2
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11931__A _12216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _13781_/Q _11669_/X _11664_/Y vssd1 vssd1 vccd1 vccd1 _13781_/D sky130_fd_sc_hd__o21a_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _10621_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _10622_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10547__A _10547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13340_ _14383_/Q _13328_/X _13336_/X _14463_/Q vssd1 vssd1 vccd1 vccd1 _13340_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11620__A1 _11619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10552_ _13964_/Q _10545_/X _10548_/X _10551_/Y vssd1 vssd1 vccd1 vccd1 _13964_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08017__A _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ _14415_/Q _13306_/A _13270_/X vssd1 vssd1 vccd1 vccd1 _13271_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10483_ _10458_/X _10461_/X _10462_/X _10482_/Y vssd1 vssd1 vccd1 vccd1 _10520_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12222_ _12222_/A vssd1 vssd1 vccd1 vccd1 _13836_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input69_A io_wbs_datwr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14472__184 vssd1 vssd1 vccd1 vccd1 _14472__184/HI io_oeb[4] sky130_fd_sc_hd__conb_1
XFILLER_68_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12153_ input77/X vssd1 vssd1 vccd1 vccd1 _12906_/A sky130_fd_sc_hd__buf_6
XFILLER_29_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11104_ _11104_/A _11104_/B _11108_/B vssd1 vssd1 vccd1 vccd1 _11104_/X sky130_fd_sc_hd__or3_1
XFILLER_2_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12084_ _13806_/Q _12000_/A _12021_/A _13822_/Q vssd1 vssd1 vccd1 vccd1 _12085_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11035_ _11035_/A _11035_/B vssd1 vssd1 vccd1 vccd1 _11052_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11439__A1 _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12002__A _12060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12986_ _13004_/A vssd1 vssd1 vccd1 vccd1 _12991_/A sky130_fd_sc_hd__buf_2
XFILLER_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13798__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11937_ _11940_/A vssd1 vssd1 vccd1 vccd1 _11937_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13532__S _13542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11868_ _14354_/Q _11870_/B vssd1 vssd1 vccd1 vccd1 _11869_/A sky130_fd_sc_hd__and2_1
XANTENNA__09311__A _09349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13607_ _13607_/A _13607_/B vssd1 vssd1 vccd1 vccd1 _13608_/A sky130_fd_sc_hd__and2_1
X_10819_ _10840_/A _10840_/B _10841_/A vssd1 vssd1 vccd1 vccd1 _10819_/X sky130_fd_sc_hd__o21ba_1
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11799_ _12773_/A vssd1 vssd1 vccd1 vccd1 _12768_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11611__A1 _11610_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13538_ input91/X _14407_/Q _13542_/S vssd1 vssd1 vccd1 vccd1 _13539_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13469_ _13469_/A vssd1 vssd1 vccd1 vccd1 _14387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_74_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_4_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07961_ _09818_/B vssd1 vssd1 vccd1 vccd1 _09434_/B sky130_fd_sc_hd__buf_2
XFILLER_4_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _09687_/A _09687_/Y _09698_/X _09699_/Y vssd1 vssd1 vccd1 vccd1 _09727_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06912_ _06894_/X _06911_/X _14358_/Q vssd1 vssd1 vccd1 vccd1 _06913_/S sky130_fd_sc_hd__o21a_1
XFILLER_68_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12611__S _12611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ _07824_/Y _07892_/B vssd1 vssd1 vccd1 vccd1 _07893_/B sky130_fd_sc_hd__and2b_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09631_ _09631_/A _09631_/B _09631_/C vssd1 vssd1 vccd1 vccd1 _09631_/Y sky130_fd_sc_hd__nand3_2
XFILLER_110_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12627__A0 _12218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _09485_/B _09485_/C _09485_/A vssd1 vssd1 vccd1 vccd1 _09563_/C sky130_fd_sc_hd__a21bo_1
XFILLER_36_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08513_ _09457_/A _09348_/B _09200_/B _08748_/B vssd1 vssd1 vccd1 vccd1 _08693_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_64_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10102__A1 _10333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09493_ _09493_/A _09493_/B _09792_/B _09493_/D vssd1 vssd1 vccd1 vccd1 _09541_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08444_ _09869_/B vssd1 vssd1 vccd1 vccd1 _09092_/C sky130_fd_sc_hd__buf_2
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08375_ _08287_/B _08287_/C _09596_/A vssd1 vssd1 vccd1 vccd1 _08376_/B sky130_fd_sc_hd__o21ai_1
X_07326_ _14224_/Q _07311_/X _07316_/X _07325_/X vssd1 vssd1 vccd1 vccd1 _14224_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07257_ _07257_/A vssd1 vssd1 vccd1 vccd1 _14261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10169__A1 _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07188_ _07259_/S vssd1 vssd1 vccd1 vccd1 _07201_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__07034__A1 _14273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09891__A _10092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11118__B1 _11100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09829_ _10435_/B _09829_/B vssd1 vssd1 vccd1 vccd1 _09901_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08300__A _09777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12840_ _12579_/X _14128_/Q _12846_/S vssd1 vssd1 vccd1 vccd1 _12841_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12618__A0 _12940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12800_/A vssd1 vssd1 vccd1 vccd1 _12771_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _13829_/Q _13770_/Q _11719_/B vssd1 vssd1 vccd1 vccd1 _11722_/X sky130_fd_sc_hd__o21ba_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14441_ _14441_/CLK _14441_/D vssd1 vssd1 vccd1 vccd1 _14441_/Q sky130_fd_sc_hd__dfxtp_1
X_11653_ _11653_/A vssd1 vssd1 vccd1 vccd1 _13841_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10604_ _10604_/A _10614_/B vssd1 vssd1 vccd1 vccd1 _10604_/Y sky130_fd_sc_hd__nand2_1
X_14372_ _14417_/CLK _14372_/D vssd1 vssd1 vccd1 vccd1 _14372_/Q sky130_fd_sc_hd__dfxtp_1
X_11584_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _11584_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_70_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14446__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13323_ _14346_/Q _13311_/X _13321_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _14346_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10535_ _10564_/A _10564_/B _10418_/X vssd1 vssd1 vccd1 vccd1 _10546_/B sky130_fd_sc_hd__a21o_1
X_13254_ _13254_/A vssd1 vssd1 vccd1 vccd1 _13254_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ _10467_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _10491_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output175_A _14300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ _12205_/A _12205_/B vssd1 vssd1 vccd1 vccd1 _12205_/X sky130_fd_sc_hd__and2_1
X_13185_ _13189_/A vssd1 vssd1 vccd1 vccd1 _13185_/Y sky130_fd_sc_hd__inv_2
X_10397_ _10382_/B _10397_/B vssd1 vssd1 vccd1 vccd1 _10397_/X sky130_fd_sc_hd__and2b_1
XFILLER_97_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12136_ _13817_/Q _12133_/X _12135_/X _12131_/X vssd1 vssd1 vccd1 vccd1 _13817_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12067_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12081_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11018_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11114_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12969_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12969_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08160_ _08160_/A _08160_/B _08160_/C vssd1 vssd1 vccd1 vccd1 _08170_/B sky130_fd_sc_hd__nor3_1
XANTENNA__09789__B1 _09788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12793__C1 _12216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07111_ _14407_/Q _07110_/Y _07087_/X vssd1 vssd1 vccd1 vccd1 _07111_/X sky130_fd_sc_hd__a21o_1
XFILLER_119_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08091_ _08091_/A _08091_/B vssd1 vssd1 vccd1 vccd1 _08093_/A sky130_fd_sc_hd__nor2_2
XFILLER_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13813__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07042_ _14416_/Q _07059_/B _14448_/Q vssd1 vssd1 vccd1 vccd1 _07042_/X sky130_fd_sc_hd__and3b_1
XFILLER_103_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13986_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08993_ _08993_/A _08993_/B _08993_/C vssd1 vssd1 vccd1 vccd1 _09045_/A sky130_fd_sc_hd__and3_1
XFILLER_102_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07944_ _08251_/A _09233_/D _08982_/B _08132_/A vssd1 vssd1 vccd1 vccd1 _07944_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_60_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08516__A1 _08867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09216__A _09216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _07875_/A vssd1 vssd1 vccd1 vccd1 _13982_/D sky130_fd_sc_hd__clkbuf_1
X_09614_ _09573_/B _09573_/Y _09611_/X _09613_/Y vssd1 vssd1 vccd1 vccd1 _09614_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_44_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ _09593_/A _09544_/Y _09545_/C _09545_/D vssd1 vssd1 vccd1 vccd1 _09593_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_34_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09476_ _08312_/A _10007_/A _09475_/A _09475_/C vssd1 vssd1 vccd1 vccd1 _09478_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08427_ _08983_/A _08449_/B _09152_/B _09091_/B vssd1 vssd1 vccd1 vccd1 _08592_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11912__A2_N _11872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ _14019_/Q vssd1 vssd1 vccd1 vccd1 _09479_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_54_io_wbs_clk clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13809_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07309_ _14165_/D _07543_/B _07301_/Y vssd1 vssd1 vccd1 vccd1 _07462_/A sky130_fd_sc_hd__a21o_2
X_08289_ _08289_/A vssd1 vssd1 vccd1 vccd1 _09962_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_4_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13201__A _13637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ _10369_/C _10320_/B vssd1 vssd1 vccd1 vccd1 _10374_/C sky130_fd_sc_hd__nand2_1
X_10251_ _10395_/A _10256_/B vssd1 vssd1 vccd1 vccd1 _10254_/B sky130_fd_sc_hd__or2b_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10182_ _10182_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10184_/B sky130_fd_sc_hd__xnor2_1
XFILLER_106_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13941_ _13947_/CLK _13941_/D _12359_/Y vssd1 vssd1 vccd1 vccd1 _13941_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13872_ _13946_/CLK _13872_/D _12273_/Y vssd1 vssd1 vccd1 vccd1 _13872_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12823_ _12828_/A _12952_/B _12823_/C vssd1 vssd1 vccd1 vccd1 _12902_/B sky130_fd_sc_hd__or3_1
XFILLER_28_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12758_/A vssd1 vssd1 vccd1 vccd1 _12754_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11710_/B vssd1 vssd1 vccd1 vccd1 _11882_/A sky130_fd_sc_hd__buf_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12940_/A _14054_/Q _12685_/S vssd1 vssd1 vccd1 vccd1 _12686_/B sky130_fd_sc_hd__mux2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14424_ _14427_/CLK _14424_/D vssd1 vssd1 vccd1 vccd1 _14424_/Q sky130_fd_sc_hd__dfxtp_1
X_11636_ _13845_/Q _11655_/B vssd1 vssd1 vccd1 vccd1 _11636_/X sky130_fd_sc_hd__and2_1
X_14478__190 vssd1 vssd1 vccd1 vccd1 _14478__190/HI io_oeb[10] sky130_fd_sc_hd__conb_1
X_14355_ _14464_/CLK _14355_/D vssd1 vssd1 vccd1 vccd1 _14355_/Q sky130_fd_sc_hd__dfxtp_1
X_11567_ _11544_/Y _11623_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _11619_/A sky130_fd_sc_hd__o21ai_4
XFILLER_10_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13306_ _13306_/A vssd1 vssd1 vccd1 vccd1 _13306_/X sky130_fd_sc_hd__clkbuf_2
X_10518_ _13968_/Q _10562_/B vssd1 vssd1 vccd1 vccd1 _10518_/X sky130_fd_sc_hd__or2_1
X_14286_ _14365_/CLK _14286_/D _13149_/Y vssd1 vssd1 vccd1 vccd1 _14286_/Q sky130_fd_sc_hd__dfrtp_4
X_11498_ _11493_/A _11497_/X _10686_/X vssd1 vssd1 vccd1 vccd1 _11498_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13237_ _14360_/Q _13236_/X _13210_/X vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__a21o_1
X_10449_ _10449_/A _10449_/B _10453_/A vssd1 vssd1 vccd1 vccd1 _10450_/B sky130_fd_sc_hd__and3_1
XFILLER_41_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13168_ _13171_/A vssd1 vssd1 vccd1 vccd1 _13168_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12119_ _12147_/A vssd1 vssd1 vccd1 vccd1 _12130_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13099_ _12645_/X hold25/A _13105_/S vssd1 vssd1 vccd1 vccd1 _13100_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07255__S _07258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__B _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07660_ _07660_/A _07660_/B vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__or2_2
XFILLER_26_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07591_ _14087_/Q input3/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07592_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _09399_/B _09329_/C _09329_/D _09329_/A vssd1 vssd1 vccd1 vccd1 _09330_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11805__B2 _14111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09261_ _09257_/X _09259_/Y _09184_/B _09184_/Y vssd1 vssd1 vccd1 vccd1 _09261_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08212_ _08212_/A _08212_/B vssd1 vssd1 vccd1 vccd1 _08214_/A sky130_fd_sc_hd__xnor2_4
X_09192_ _09635_/A _09192_/B vssd1 vssd1 vccd1 vccd1 _09192_/Y sky130_fd_sc_hd__nor2_2
XFILLER_105_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08143_ _08144_/B _08144_/C _08144_/A vssd1 vssd1 vccd1 vccd1 _08221_/B sky130_fd_sc_hd__o21ai_1
XFILLER_53_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13021__A _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ _08125_/A _08125_/B vssd1 vssd1 vccd1 vccd1 _08076_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07025_ _14418_/Q _07024_/Y _07009_/X vssd1 vssd1 vccd1 vccd1 _07025_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12860__A _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__buf_2
X_08976_ _08976_/A vssd1 vssd1 vccd1 vccd1 _09857_/A sky130_fd_sc_hd__buf_4
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__07165__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13494__A0 _12654_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07927_ _08132_/A vssd1 vssd1 vccd1 vccd1 _08249_/A sky130_fd_sc_hd__buf_2
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07858_ _14038_/Q _13984_/Q vssd1 vssd1 vccd1 vccd1 _07858_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07789_ _10655_/A _07806_/B _07786_/A vssd1 vssd1 vccd1 vccd1 _10875_/S sky130_fd_sc_hd__nor3b_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _09515_/A _09528_/B vssd1 vssd1 vccd1 vccd1 _09528_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12100__A _12924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07476__A1 _14079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ _09459_/A _09459_/B _09459_/C vssd1 vssd1 vccd1 vccd1 _09462_/A sky130_fd_sc_hd__or3_1
XFILLER_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12470_ _14031_/Q _12464_/X _12469_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _12470_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11421_ _11511_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11506_/A sky130_fd_sc_hd__or2_1
X_14140_ _14149_/CLK _14140_/D vssd1 vssd1 vccd1 vccd1 _14140_/Q sky130_fd_sc_hd__dfxtp_2
X_11352_ _11269_/A _10904_/X _11351_/Y _07784_/X vssd1 vssd1 vccd1 vccd1 _13896_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12509__C1 _12216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ _10420_/B _10328_/B vssd1 vssd1 vccd1 vccd1 _10310_/A sky130_fd_sc_hd__xor2_1
X_14071_ _14075_/CLK _14071_/D _12714_/Y vssd1 vssd1 vccd1 vccd1 _14071_/Q sky130_fd_sc_hd__dfrtp_2
X_11283_ _11333_/B _11283_/B vssd1 vssd1 vccd1 vccd1 _11336_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13022_ _13022_/A vssd1 vssd1 vccd1 vccd1 _13022_/Y sky130_fd_sc_hd__inv_2
X_10234_ _10236_/A _10236_/B _10231_/Y _10233_/Y vssd1 vssd1 vccd1 vccd1 _10234_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_input51_A io_wbs_adr[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10165_ _10155_/Y _10182_/B _10164_/Y vssd1 vssd1 vccd1 vccd1 _10168_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10096_ _10138_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _10096_/X sky130_fd_sc_hd__and2_1
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output138_A _11807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13924_ _13927_/CLK _13924_/D _12338_/Y vssd1 vssd1 vccd1 vccd1 _13924_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_75_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08695__A _13861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08900__A1 _08937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07703__A2 _07548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13855_ _13892_/CLK _13855_/D _12250_/Y vssd1 vssd1 vccd1 vccd1 _13855_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12806_ _14116_/Q _12800_/X _12804_/X _12805_/X vssd1 vssd1 vccd1 vccd1 _14116_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12010__A _12216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10998_ _11076_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__nand2_1
X_13786_ _13809_/CLK _13786_/D vssd1 vssd1 vccd1 vccd1 _13786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07467__A1 _14081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12740_/A vssd1 vssd1 vccd1 vccd1 _12737_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12668_ input67/X vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__buf_4
X_14407_ _14442_/CLK _14407_/D vssd1 vssd1 vccd1 vccd1 _14407_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07219__A1 _07218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ _11619_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _11619_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_117_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12599_ _12599_/A vssd1 vssd1 vccd1 vccd1 _14032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08580__D _09870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14338_ _14400_/CLK _14338_/D vssd1 vssd1 vccd1 vccd1 _14338_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_13_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14269_ _14365_/CLK _14269_/D _13128_/Y vssd1 vssd1 vccd1 vccd1 _14269_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12680__A _13072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10526__A1 _10597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _08830_/A _08830_/B vssd1 vssd1 vccd1 vccd1 _08861_/C sky130_fd_sc_hd__xnor2_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08760_/A _08760_/B _08760_/C vssd1 vssd1 vccd1 vccd1 _08762_/C sky130_fd_sc_hd__a21oi_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07712_ _07712_/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__clkbuf_1
XFILLER_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08692_ _08692_/A _08965_/A vssd1 vssd1 vccd1 vccd1 _09038_/A sky130_fd_sc_hd__xnor2_2
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07643_ _07666_/A _07667_/A _07642_/Y vssd1 vssd1 vccd1 vccd1 _07664_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07574_ _14095_/Q input11/X _07582_/S vssd1 vssd1 vccd1 vccd1 _07575_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ _09313_/A _09313_/B _09313_/C vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__nand3_2
XFILLER_81_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09244_ _09239_/A _09239_/B _09239_/C vssd1 vssd1 vccd1 vccd1 _09245_/C sky130_fd_sc_hd__a21o_1
XANTENNA__10273__B1_N _10272_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09175_ _09175_/A _09175_/B vssd1 vssd1 vccd1 vccd1 _09198_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_5_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14211_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08126_ _08126_/A vssd1 vssd1 vccd1 vccd1 _08128_/B sky130_fd_sc_hd__buf_4
XFILLER_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08057_ _13871_/Q vssd1 vssd1 vccd1 vccd1 _09493_/D sky130_fd_sc_hd__clkbuf_2
X_07008_ _14452_/Q _14276_/Q vssd1 vssd1 vccd1 vccd1 _07008_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09383__A1 _09553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09383__B2 _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13467__A0 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _08856_/A _08856_/C _08856_/B vssd1 vssd1 vccd1 vccd1 _08959_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11934__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _11970_/A vssd1 vssd1 vccd1 vccd1 _13774_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09404__A _09641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ _10652_/X _10917_/X _10920_/X vssd1 vssd1 vccd1 vccd1 _10987_/A sky130_fd_sc_hd__o21ai_2
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13640_ _12827_/X _14436_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13641_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10852_ _10845_/X _10849_/X _10851_/Y vssd1 vssd1 vccd1 vccd1 _13939_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__09123__B _09457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_25_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _13571_/A vssd1 vssd1 vccd1 vccd1 _14416_/D sky130_fd_sc_hd__clkbuf_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10783_ _10783_/A _10783_/B vssd1 vssd1 vccd1 vccd1 _10786_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12522_ _12522_/A vssd1 vssd1 vccd1 vccd1 _14010_/D sky130_fd_sc_hd__clkbuf_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input99_A io_wbs_stb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12453_ _13992_/Q _12422_/X _12452_/X _12203_/X vssd1 vssd1 vccd1 vccd1 _13992_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14187__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ _13878_/Q _11392_/X _11396_/X _11403_/X vssd1 vssd1 vccd1 vccd1 _13878_/D
+ sky130_fd_sc_hd__a22o_1
X_12384_ _12384_/A vssd1 vssd1 vccd1 vccd1 _12384_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_4_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11335_ _11285_/A _11319_/X _11334_/X _11322_/X vssd1 vssd1 vccd1 vccd1 _13902_/D
+ sky130_fd_sc_hd__o22a_1
X_14123_ _14164_/CLK _14123_/D vssd1 vssd1 vccd1 vccd1 _14123_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11266_ _13894_/Q vssd1 vssd1 vccd1 vccd1 _11355_/A sky130_fd_sc_hd__clkbuf_2
X_14054_ _14054_/CLK _14054_/D vssd1 vssd1 vccd1 vccd1 _14054_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10217_ _10067_/A _10216_/X _10061_/X _10054_/B vssd1 vssd1 vccd1 vccd1 _10217_/X
+ sky130_fd_sc_hd__o211a_1
X_13005_ _13009_/A vssd1 vssd1 vccd1 vccd1 _13005_/Y sky130_fd_sc_hd__inv_2
X_11197_ _10651_/A _11152_/X _11143_/X vssd1 vssd1 vccd1 vccd1 _11221_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12005__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10148_ _10149_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10636_/A sky130_fd_sc_hd__or2_1
XANTENNA__09126__A1 _09508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13535__S _13542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__B2 _08445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10079_ _10079_/A _10079_/B vssd1 vssd1 vccd1 vccd1 _10106_/A sky130_fd_sc_hd__xnor2_2
XFILLER_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13907_ _13949_/CLK _13907_/D _12316_/Y vssd1 vssd1 vccd1 vccd1 _13907_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13838_ _14259_/CLK _13838_/D vssd1 vssd1 vccd1 vccd1 _13838_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13769_ _13820_/CLK _13769_/D _11962_/Y vssd1 vssd1 vccd1 vccd1 _13769_/Q sky130_fd_sc_hd__dfrtp_1
X_07290_ _07290_/A vssd1 vssd1 vccd1 vccd1 _14229_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07860__A1 _14038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07073__C1 _14364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09931_ _10090_/B vssd1 vssd1 vccd1 vccd1 _10195_/A sky130_fd_sc_hd__buf_2
XANTENNA__09365__A1 _09425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _09966_/C _09862_/B vssd1 vssd1 vccd1 vccd1 _09880_/A sky130_fd_sc_hd__nand2_1
XFILLER_113_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08813_ _08811_/A _08811_/Y _08812_/Y _08772_/B vssd1 vssd1 vccd1 vccd1 _08818_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07009__A _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09793_ _09793_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__xnor2_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08744_ _08709_/A _08708_/B _08708_/C vssd1 vssd1 vccd1 vccd1 _08760_/B sky130_fd_sc_hd__a21o_1
XFILLER_39_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08675_ _08971_/B _08675_/B _08675_/C _08675_/D vssd1 vssd1 vccd1 vccd1 _08675_/Y
+ sky130_fd_sc_hd__nor4_4
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10683__A0 _10826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07626_ _07626_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__nand2_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13621__A0 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07557_ _07557_/A vssd1 vssd1 vccd1 vccd1 _14103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07488_ _07348_/A _07486_/X _07487_/X _07373_/A _14193_/Q vssd1 vssd1 vccd1 vccd1
+ _14193_/D sky130_fd_sc_hd__a32o_1
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09227_ _09227_/A _09227_/B vssd1 vssd1 vccd1 vccd1 _09277_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09158_ _09158_/A _09158_/B _09158_/C vssd1 vssd1 vccd1 vccd1 _09161_/A sky130_fd_sc_hd__nand3_1
X_08109_ _08595_/A _08791_/B _09821_/A vssd1 vssd1 vccd1 vccd1 _09535_/A sky130_fd_sc_hd__and3_1
XFILLER_108_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09089_ _09087_/A _09087_/C _09087_/B vssd1 vssd1 vccd1 vccd1 _09090_/C sky130_fd_sc_hd__a21o_1
XFILLER_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11120_ _11059_/X _11120_/B _11120_/C vssd1 vssd1 vccd1 vccd1 _11120_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _11129_/A _11129_/B vssd1 vssd1 vccd1 vccd1 _11127_/C sky130_fd_sc_hd__or2_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10002_ _10420_/B vssd1 vssd1 vccd1 vccd1 _10421_/B sky130_fd_sc_hd__buf_2
XFILLER_107_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09134__A _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input14_A dout1[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _11953_/A vssd1 vssd1 vccd1 vccd1 _11953_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10904_ _11319_/A vssd1 vssd1 vccd1 vccd1 _10904_/X sky130_fd_sc_hd__buf_2
X_11884_ _11888_/B vssd1 vssd1 vccd1 vccd1 _11884_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13623_ _13623_/A vssd1 vssd1 vccd1 vccd1 _14431_/D sky130_fd_sc_hd__clkbuf_1
X_10835_ _10835_/A _10835_/B vssd1 vssd1 vccd1 vccd1 _10835_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11603__S _11611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _13554_/A vssd1 vssd1 vccd1 vccd1 _14411_/D sky130_fd_sc_hd__clkbuf_1
X_10766_ _10715_/A _10670_/Y _10748_/B _10765_/X vssd1 vssd1 vccd1 vccd1 _10767_/B
+ sky130_fd_sc_hd__o211a_1
X_12505_ _14057_/Q _12442_/X _12435_/X vssd1 vssd1 vccd1 vccd1 _12505_/X sky130_fd_sc_hd__a21o_1
X_13485_ _13485_/A _13485_/B vssd1 vssd1 vccd1 vccd1 _13486_/A sky130_fd_sc_hd__and2_1
X_10697_ _11236_/A vssd1 vssd1 vccd1 vccd1 _11228_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12436_ _12425_/X _12432_/X _12435_/X vssd1 vssd1 vccd1 vccd1 _12436_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12367_ _12379_/A vssd1 vssd1 vccd1 vccd1 _12372_/A sky130_fd_sc_hd__buf_4
XFILLER_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14106_ _14107_/CLK _14106_/D _12757_/Y vssd1 vssd1 vccd1 vccd1 _14106_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_114_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11318_ _11119_/X _11315_/C _11317_/X _10851_/B _11300_/A vssd1 vssd1 vccd1 vccd1
+ _13907_/D sky130_fd_sc_hd__a32o_1
X_12298_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12298_/Y sky130_fd_sc_hd__inv_2
X_11249_ _11249_/A _11249_/B vssd1 vssd1 vccd1 vccd1 _11273_/B sky130_fd_sc_hd__xnor2_1
X_14037_ _14367_/CLK _14037_/D vssd1 vssd1 vccd1 vccd1 _14037_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_80_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11574__A _14052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__B _07921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09044__A _09044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08460_ _09875_/A vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__08246__B_N _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07530__B1 _07521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07411_ _14207_/Q _14209_/Q _07415_/S vssd1 vssd1 vccd1 vccd1 _07412_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13603__A0 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08391_ _08391_/A _08391_/B _08391_/C vssd1 vssd1 vccd1 vccd1 _08391_/X sky130_fd_sc_hd__or3_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07342_ _14221_/Q _07311_/X _07316_/X _07341_/X vssd1 vssd1 vccd1 vccd1 _14221_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10968__A1 _10722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__B2 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07273_ _07274_/A _07308_/A _14166_/Q vssd1 vssd1 vccd1 vccd1 _07307_/B sky130_fd_sc_hd__o21a_1
X_09012_ _09153_/A _09153_/B _09092_/D _09085_/B vssd1 vssd1 vccd1 vccd1 _09014_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10653__A _10875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12590__A0 _12919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09914_ _09914_/A _09914_/B vssd1 vssd1 vccd1 vccd1 _09940_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07962__A _09803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _09091_/B _09843_/X _09844_/X vssd1 vssd1 vccd1 vccd1 _10126_/A sky130_fd_sc_hd__a21oi_4
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A dout1[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12893__A1 _14145_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09776_ _08266_/A _08266_/B _09775_/X vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__o21ba_1
XFILLER_86_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06988_ _07027_/A vssd1 vssd1 vccd1 vccd1 _07020_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08727_ _08727_/A _08727_/B vssd1 vssd1 vccd1 vccd1 _08729_/A sky130_fd_sc_hd__and2_1
XFILLER_6_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08980_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _08664_/A sky130_fd_sc_hd__nand2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07609_ _14079_/Q input26/X _07615_/S vssd1 vssd1 vccd1 vccd1 _07610_/A sky130_fd_sc_hd__mux2_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08619_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _08611_/A sky130_fd_sc_hd__xor2_1
XFILLER_109_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13204__A _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _10627_/A _10627_/B _09273_/A vssd1 vssd1 vccd1 vccd1 _10621_/B sky130_fd_sc_hd__a21boi_1
XFILLER_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ _10540_/B _10549_/X _10550_/X vssd1 vssd1 vccd1 vccd1 _10551_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13270_ _14447_/Q _13250_/X _13245_/X _14399_/Q vssd1 vssd1 vccd1 vccd1 _13270_/X
+ sky130_fd_sc_hd__a22o_1
X_10482_ _10520_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10482_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12221_ _12517_/A _12221_/B vssd1 vssd1 vccd1 vccd1 _12222_/A sky130_fd_sc_hd__and2_1
XFILLER_108_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ _13823_/Q _12146_/X _12151_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _13823_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08033__A _14017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ _10831_/X _11099_/C _11102_/X _11100_/X _11076_/A vssd1 vssd1 vccd1 vccd1
+ _13923_/D sky130_fd_sc_hd__a32o_1
X_12083_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12517_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08968__A _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11136__B2 _10826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _11252_/A _11039_/A _11039_/B vssd1 vssd1 vccd1 vccd1 _11035_/B sky130_fd_sc_hd__o21ai_1
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12985_ _12985_/A vssd1 vssd1 vccd1 vccd1 _12985_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11936_ _11940_/A vssd1 vssd1 vccd1 vccd1 _11936_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _11867_/A vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__06935__B _06942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13606_ input81/X _14427_/Q _13611_/S vssd1 vssd1 vccd1 vccd1 _13607_/B sky130_fd_sc_hd__mux2_1
XFILLER_14_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13061__A1 _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10818_ _13940_/Q _10818_/B vssd1 vssd1 vccd1 vccd1 _10841_/A sky130_fd_sc_hd__xnor2_1
X_11798_ _13035_/A vssd1 vssd1 vccd1 vccd1 _13037_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08208__A _08249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13537_ _13537_/A vssd1 vssd1 vccd1 vccd1 _14406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10749_ _10730_/A _10735_/X _10748_/X vssd1 vssd1 vccd1 vccd1 _10750_/S sky130_fd_sc_hd__o21a_1
XFILLER_71_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09017__B1 _08547_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13468_ _13485_/A _13468_/B vssd1 vssd1 vccd1 vccd1 _13469_/A sky130_fd_sc_hd__and2_1
X_12419_ _12703_/A vssd1 vssd1 vccd1 vccd1 _12419_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_12_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13399_ _12673_/X _14367_/Q _13408_/S vssd1 vssd1 vccd1 vccd1 _13400_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12572__A0 _12515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07258__S _07258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11288__B _11288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09400__A2_N _08091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07960_ _09084_/B vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_io_wbs_clk clkbuf_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_io_wbs_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_96_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06911_ _14406_/Q _06942_/B _14438_/Q vssd1 vssd1 vccd1 vccd1 _06911_/X sky130_fd_sc_hd__and3b_1
XFILLER_110_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07891_ _13978_/Q _07890_/A _07890_/Y _07848_/B vssd1 vssd1 vccd1 vccd1 _13978_/D
+ sky130_fd_sc_hd__a22o_1
X_09630_ _09470_/X _09624_/X _09396_/C _09396_/Y vssd1 vssd1 vccd1 vccd1 _09631_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_95_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09561_ _09560_/B _09560_/C _09560_/A vssd1 vssd1 vccd1 vccd1 _09563_/B sky130_fd_sc_hd__a21o_1
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09669__A_N _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08512_ _13863_/Q vssd1 vssd1 vccd1 vccd1 _09200_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_24_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09492_ _09543_/B _09543_/D _09493_/D _09443_/A vssd1 vssd1 vccd1 vccd1 _09494_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08443_ _13863_/Q vssd1 vssd1 vccd1 vccd1 _09869_/B sky130_fd_sc_hd__buf_2
XFILLER_24_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08374_ _08571_/A _08980_/B _08362_/A _08360_/B vssd1 vssd1 vccd1 vccd1 _08384_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_56_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07325_ _11925_/S _14223_/Q _07521_/B _07321_/X _07324_/X vssd1 vssd1 vccd1 vccd1
+ _07325_/X sky130_fd_sc_hd__a32o_1
XFILLER_108_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14465_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_108_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07256_ _14261_/Q _07255_/X _07259_/S vssd1 vssd1 vccd1 vccd1 _07257_/A sky130_fd_sc_hd__mux2_1
XANTENNA__07957__A _13868_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07282__A2 _14166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13355__A2 _13216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07187_ _14097_/Q _07185_/X _07186_/X vssd1 vssd1 vccd1 vccd1 _07187_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14398__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11118__B2 _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09828_ _09926_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _10435_/A sky130_fd_sc_hd__nor2_4
XFILLER_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12103__A _12926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12618__A1 _14038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ _09759_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10629__A0 _13954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11942__A _11971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12760_/X _12767_/X _12769_/X _12498_/X vssd1 vssd1 vccd1 vccd1 _14108_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _13770_/Q _11714_/X _11716_/X _11720_/Y vssd1 vssd1 vccd1 vccd1 _13770_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14440_/CLK _14440_/D vssd1 vssd1 vccd1 vccd1 _14440_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _13841_/Q _11651_/Y _11652_/S vssd1 vssd1 vccd1 vccd1 _11653_/A sky130_fd_sc_hd__mux2_1
XANTENNA__08028__A _14017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10603_ _10613_/A _10613_/B _10613_/C vssd1 vssd1 vccd1 vccd1 _10614_/B sky130_fd_sc_hd__o21ai_1
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14371_ _14417_/CLK _14371_/D vssd1 vssd1 vccd1 vccd1 _14371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11583_ _11587_/B _11587_/C _11587_/A vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__o21bai_1
XFILLER_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13322_ _13343_/A vssd1 vssd1 vccd1 vccd1 _13322_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input81_A io_wbs_datwr[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10534_ _10534_/A vssd1 vssd1 vccd1 vccd1 _13966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13253_ _14363_/Q _13215_/X _13252_/X _13222_/X vssd1 vssd1 vccd1 vccd1 _13253_/X
+ sky130_fd_sc_hd__a211o_1
X_10465_ _10465_/A _10465_/B vssd1 vssd1 vccd1 vccd1 _10467_/B sky130_fd_sc_hd__xor2_1
X_12204_ _13833_/Q _12202_/C _12202_/Y _12203_/X vssd1 vssd1 vccd1 vccd1 _13833_/D
+ sky130_fd_sc_hd__o211a_1
X_13184_ _13184_/A vssd1 vssd1 vccd1 vccd1 _13189_/A sky130_fd_sc_hd__buf_2
X_10396_ _10396_/A vssd1 vssd1 vccd1 vccd1 _10396_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output168_A _14322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12135_ input75/X _12143_/B vssd1 vssd1 vccd1 vccd1 _12135_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_18_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08698__A _08791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__A1 _11007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ _12066_/A vssd1 vssd1 vccd1 vccd1 _13800_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13765__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11017_ _11017_/A _11017_/B vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__xnor2_1
XFILLER_93_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13109__A _13115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08930__C1 _10061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12968_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12968_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11919_ hold5/X _11919_/B vssd1 vssd1 vccd1 vccd1 _13761_/D sky130_fd_sc_hd__nor2_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11832__A2 _11808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12899_ _14148_/Q _12885_/A _12898_/X _12892_/X vssd1 vssd1 vccd1 vccd1 _14148_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13034__B2 _14240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09789__A1 _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07110_ _14439_/Q _14263_/Q vssd1 vssd1 vccd1 vccd1 _07110_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08090_ _08796_/A _08828_/B _09821_/A vssd1 vssd1 vccd1 vccd1 _08091_/B sky130_fd_sc_hd__o21ai_1
XFILLER_118_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07041_ _14272_/Q _07007_/X _07040_/X _14368_/Q vssd1 vssd1 vccd1 vccd1 _07041_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08992_ _08991_/B _08991_/C _08991_/A vssd1 vssd1 vccd1 vccd1 _08993_/C sky130_fd_sc_hd__a21o_1
X_07943_ _09818_/B vssd1 vssd1 vccd1 vccd1 _08982_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13019__A _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__A1 _08403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07874_ _07873_/X _13982_/Q _07874_/S vssd1 vssd1 vccd1 vccd1 _07875_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11520__A1 _10061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09613_ _09708_/B _09708_/C _09708_/A vssd1 vssd1 vccd1 vccd1 _09613_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _08580_/B _09543_/C _09792_/B _08580_/A vssd1 vssd1 vccd1 vccd1 _09544_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09475_ _09475_/A _09475_/B _09475_/C vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__nand3_1
X_08426_ _09806_/A vssd1 vssd1 vccd1 vccd1 _09091_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08357_ _14020_/Q vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07308_ _07308_/A _07319_/A vssd1 vssd1 vccd1 vccd1 _07543_/B sky130_fd_sc_hd__nor2_2
X_08288_ _08287_/B _08376_/A vssd1 vssd1 vccd1 vccd1 _08323_/A sky130_fd_sc_hd__and2b_1
XFILLER_30_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07239_ _14082_/Q _13882_/Q _07252_/S vssd1 vssd1 vccd1 vccd1 _07239_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10250_ _10250_/A _10250_/B vssd1 vssd1 vccd1 vccd1 _10256_/B sky130_fd_sc_hd__xor2_1
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_9_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13628__S _13628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _10188_/A _10188_/B _10180_/B _10227_/A _10227_/B vssd1 vssd1 vccd1 vccd1
+ _10183_/A sky130_fd_sc_hd__o32a_1
XFILLER_105_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13940_ _13947_/CLK _13940_/D _12358_/Y vssd1 vssd1 vccd1 vccd1 _13940_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13871_ _13946_/CLK _13871_/D _12272_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__07191__A1 _14096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12822_ _14123_/Q _12771_/X _12821_/X _12817_/X vssd1 vssd1 vccd1 vccd1 _14123_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14413__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _12753_/A vssd1 vssd1 vccd1 vccd1 _12758_/A sky130_fd_sc_hd__buf_2
XFILLER_37_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _13762_/Q _11920_/C vssd1 vssd1 vccd1 vccd1 _11710_/B sky130_fd_sc_hd__or2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12684_/A vssd1 vssd1 vccd1 vccd1 _14053_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14423_ _14427_/CLK _14423_/D vssd1 vssd1 vccd1 vccd1 _14423_/Q sky130_fd_sc_hd__dfxtp_1
X_11635_ _11634_/A _11634_/B _11634_/C vssd1 vssd1 vccd1 vccd1 _11635_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_11_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11611__S _11611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ _14354_/CLK _14354_/D vssd1 vssd1 vccd1 vccd1 _14354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11566_ _14048_/Q _13960_/Q vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ _14342_/Q _13289_/X _13304_/X _13301_/X vssd1 vssd1 vccd1 vccd1 _14342_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10517_ _10629_/S vssd1 vssd1 vccd1 vccd1 _10562_/B sky130_fd_sc_hd__buf_4
X_14285_ _14365_/CLK _14285_/D _13148_/Y vssd1 vssd1 vccd1 vccd1 _14285_/Q sky130_fd_sc_hd__dfrtp_4
X_11497_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11497_/X sky130_fd_sc_hd__and2_1
XANTENNA__12008__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12527__A0 _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13236_ _13236_/A vssd1 vssd1 vccd1 vccd1 _13236_/X sky130_fd_sc_hd__buf_2
XFILLER_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10448_ _10449_/B _10453_/A _10449_/A vssd1 vssd1 vccd1 vccd1 _10450_/A sky130_fd_sc_hd__a21oi_1
XFILLER_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13538__S _13542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11847__A _11870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _13171_/A vssd1 vssd1 vccd1 vccd1 _13167_/Y sky130_fd_sc_hd__inv_2
X_10379_ _10407_/A vssd1 vssd1 vccd1 vccd1 _10478_/A sky130_fd_sc_hd__clkbuf_2
X_12118_ input70/X vssd1 vssd1 vccd1 vccd1 _12938_/A sky130_fd_sc_hd__buf_6
X_13098_ _13098_/A vssd1 vssd1 vccd1 vccd1 _14250_/D sky130_fd_sc_hd__clkbuf_1
X_12049_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12065_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07182__A1 _14098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11582__A _14056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07590_ _07590_/A vssd1 vssd1 vccd1 vccd1 _14088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14093__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09260_ _09184_/B _09184_/Y _09257_/X _09259_/Y vssd1 vssd1 vccd1 vccd1 _09263_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08891__A _08891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ _08208_/X _08211_/B vssd1 vssd1 vccd1 vccd1 _08212_/B sky130_fd_sc_hd__and2b_1
X_09191_ _09191_/A _09191_/B vssd1 vssd1 vccd1 vccd1 _09191_/Y sky130_fd_sc_hd__nor2_2
XFILLER_14_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08142_ _08215_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__xor2_1
XFILLER_105_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10645__B _10645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08985__A2 _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ _08131_/A _08073_/B vssd1 vssd1 vccd1 vccd1 _08125_/B sky130_fd_sc_hd__xor2_1
X_07024_ _14450_/Q _14274_/Q vssd1 vssd1 vccd1 vccd1 _07024_/Y sky130_fd_sc_hd__nand2_1
XFILLER_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11741__A1 _13824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08975_ _08639_/B _08639_/C _08639_/A vssd1 vssd1 vccd1 vccd1 _08993_/A sky130_fd_sc_hd__a21bo_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07926_ _09472_/A vssd1 vssd1 vccd1 vccd1 _08132_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13494__A1 _14395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07970__A _14019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14436__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07857_ _07868_/A _07869_/A vssd1 vssd1 vccd1 vccd1 _07857_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07173__A1 _14101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06920__A1 _14320_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07788_ _11452_/A _11452_/B _10664_/B vssd1 vssd1 vccd1 vccd1 _11510_/A sky130_fd_sc_hd__or3b_4
XFILLER_25_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09527_ _09527_/A _09527_/B _09527_/C vssd1 vssd1 vccd1 vccd1 _09527_/X sky130_fd_sc_hd__and3_1
XFILLER_40_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09458_ _08823_/A _09821_/B _09792_/A _08445_/X vssd1 vssd1 vccd1 vccd1 _09459_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_51_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08409_ _09749_/C _08409_/B vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09389_ _09376_/A _09376_/B _09376_/C vssd1 vssd1 vccd1 vccd1 _09423_/C sky130_fd_sc_hd__a21o_1
XFILLER_32_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ _11276_/A _11056_/A _11425_/S vssd1 vssd1 vccd1 vccd1 _11511_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08306__A _13867_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ _11351_/A _11351_/B vssd1 vssd1 vccd1 vccd1 _11351_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__06987__A1 _14261_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10302_ _10302_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10328_/B sky130_fd_sc_hd__xnor2_1
X_14070_ _14075_/CLK _14070_/D _12713_/Y vssd1 vssd1 vccd1 vccd1 _14070_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11282_ _11282_/A _11282_/B vssd1 vssd1 vccd1 vccd1 _11283_/B sky130_fd_sc_hd__or2_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13021_ _13022_/A vssd1 vssd1 vccd1 vccd1 _13021_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10233_ _10271_/B _10233_/B vssd1 vssd1 vccd1 vccd1 _10233_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10164_ _10164_/A _10164_/B vssd1 vssd1 vccd1 vccd1 _10164_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_input44_A io_wbs_adr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10095_ _10333_/A _10095_/B vssd1 vssd1 vccd1 vccd1 _10139_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13923_ _13927_/CLK _13923_/D _12337_/Y vssd1 vssd1 vccd1 vccd1 _13923_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12498__A _12817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07164__A1 _14103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08900__A2 _10061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13237__A1 _14360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _14107_/CLK _13854_/D _12249_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11248__B1 _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ _12817_/A vssd1 vssd1 vccd1 vccd1 _12805_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13785_ _13809_/CLK _13785_/D vssd1 vssd1 vccd1 vccd1 _13785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10997_ _10997_/A _10997_/B vssd1 vssd1 vccd1 vccd1 _11076_/B sky130_fd_sc_hd__xnor2_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _12740_/A vssd1 vssd1 vccd1 vccd1 _12736_/Y sky130_fd_sc_hd__inv_2
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13953__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12667_ _12667_/A vssd1 vssd1 vccd1 vccd1 _14049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14406_ _14450_/CLK _14406_/D vssd1 vssd1 vccd1 vccd1 _14406_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13122__A _13153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11618_ _14049_/Q _13961_/Q vssd1 vssd1 vccd1 vccd1 _11619_/B sky130_fd_sc_hd__xnor2_2
X_12598_ _12615_/A _12598_/B vssd1 vssd1 vccd1 vccd1 _12599_/A sky130_fd_sc_hd__and2_1
XFILLER_117_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14337_ _14400_/CLK _14337_/D vssd1 vssd1 vccd1 vccd1 _14337_/Q sky130_fd_sc_hd__dfxtp_1
X_11549_ _14042_/Q _13954_/Q vssd1 vssd1 vccd1 vccd1 _11646_/A sky130_fd_sc_hd__nor2_1
XANTENNA__14309__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14268_ _14365_/CLK _14268_/D _13127_/Y vssd1 vssd1 vccd1 vccd1 _14268_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_83_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13219_ _14437_/Q _13336_/A _13218_/X _14389_/Q vssd1 vssd1 vccd1 vccd1 _13219_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _14224_/CLK _14199_/D _12990_/Y vssd1 vssd1 vccd1 vccd1 _14199_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08760_ _08760_/A _08760_/B _08760_/C vssd1 vssd1 vccd1 vccd1 _08774_/B sky130_fd_sc_hd__and3_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07790__A _10875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07711_ _14074_/Q _07709_/X _07730_/S vssd1 vssd1 vccd1 vccd1 _07712_/A sky130_fd_sc_hd__mux2_1
X_08691_ _08964_/A _08964_/B vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07155__A1 _14106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07642_ _14132_/Q _14067_/Q vssd1 vssd1 vccd1 vccd1 _07642_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07573_ _07595_/A vssd1 vssd1 vccd1 vccd1 _07582_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09312_ _08823_/A _09543_/D _09493_/D _08445_/X vssd1 vssd1 vccd1 vccd1 _09313_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09243_ _09319_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09245_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09174_ _09173_/B _09173_/C _09173_/A vssd1 vssd1 vccd1 vccd1 _09175_/B sky130_fd_sc_hd__a21oi_1
XFILLER_108_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11411__A0 _13895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _08125_/A _08125_/B vssd1 vssd1 vccd1 vccd1 _08144_/C sky130_fd_sc_hd__and2_1
XFILLER_107_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08056_ _13872_/Q vssd1 vssd1 vccd1 vccd1 _09543_/D sky130_fd_sc_hd__clkbuf_2
X_07007_ _07085_/A vssd1 vssd1 vccd1 vccd1 _07007_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09383__A2 _09074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08958_ _08887_/Y _08913_/Y _08924_/Y _08956_/Y _08957_/Y vssd1 vssd1 vccd1 vccd1
+ _08958_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07909_ _07909_/A _07909_/B _07909_/C vssd1 vssd1 vccd1 vccd1 _07911_/A sky130_fd_sc_hd__and3_1
XFILLER_57_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08889_ _09241_/A vssd1 vssd1 vccd1 vccd1 _08891_/A sky130_fd_sc_hd__buf_4
XFILLER_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10920_ _10920_/A vssd1 vssd1 vccd1 vccd1 _10920_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13207__A _13328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10851_ _13939_/Q _10851_/B vssd1 vssd1 vccd1 vccd1 _10851_/Y sky130_fd_sc_hd__nand2_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _13573_/A _13570_/B vssd1 vssd1 vccd1 vccd1 _13571_/A sky130_fd_sc_hd__and2_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10782_/A _10905_/B vssd1 vssd1 vccd1 vccd1 _10783_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12534_/A _12521_/B vssd1 vssd1 vccd1 vccd1 _12522_/A sky130_fd_sc_hd__and2_1
XFILLER_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12452_ _14027_/Q _12438_/X _12449_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _12452_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11403_ hold22/X _11403_/B vssd1 vssd1 vccd1 vccd1 _11403_/X sky130_fd_sc_hd__or2_1
X_12383_ _12384_/A vssd1 vssd1 vccd1 vccd1 _12383_/Y sky130_fd_sc_hd__inv_2
X_14122_ _14164_/CLK _14122_/D vssd1 vssd1 vccd1 vccd1 _14122_/Q sky130_fd_sc_hd__dfxtp_1
X_11334_ _11334_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11334_/X sky130_fd_sc_hd__and2_1
XANTENNA__07082__B1 _14363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14053_ _14054_/CLK _14053_/D vssd1 vssd1 vccd1 vccd1 _14053_/Q sky130_fd_sc_hd__dfxtp_2
X_11265_ _11264_/B _11264_/C _11264_/A vssd1 vssd1 vccd1 vccd1 _11268_/B sky130_fd_sc_hd__o21ai_1
XFILLER_106_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ _13004_/A vssd1 vssd1 vccd1 vccd1 _13009_/A sky130_fd_sc_hd__buf_2
X_10216_ _10216_/A _10216_/B vssd1 vssd1 vccd1 vccd1 _10216_/X sky130_fd_sc_hd__xor2_1
XFILLER_80_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output150_A _14306_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196_ _11228_/B _11229_/A _11225_/A vssd1 vssd1 vccd1 vccd1 _11220_/B sky130_fd_sc_hd__and3_1
XFILLER_80_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _10151_/A _10145_/Y _10146_/X vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__o21a_2
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10078_ _10076_/Y _10078_/B vssd1 vssd1 vccd1 vccd1 _10079_/B sky130_fd_sc_hd__and2b_1
XFILLER_43_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13906_ _13949_/CLK _13906_/D _12315_/Y vssd1 vssd1 vccd1 vccd1 _13906_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__12021__A _12021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13837_ _14365_/CLK _13837_/D vssd1 vssd1 vccd1 vccd1 _13837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13768_ _13820_/CLK _13768_/D _11961_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12719_ _12721_/A vssd1 vssd1 vccd1 vccd1 _12719_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13699_ _13712_/A _13699_/B vssd1 vssd1 vccd1 vccd1 _13700_/A sky130_fd_sc_hd__and2_1
XFILLER_102_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09930_ _10090_/A _09930_/B vssd1 vssd1 vccd1 vccd1 _09978_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09365__A2 _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _10305_/B _09861_/B vssd1 vssd1 vccd1 vccd1 _09862_/B sky130_fd_sc_hd__or2_1
XFILLER_113_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _08771_/A _08771_/B _08771_/C vssd1 vssd1 vccd1 vccd1 _08812_/Y sky130_fd_sc_hd__a21oi_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _09792_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__xnor2_4
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08743_/A _08743_/B vssd1 vssd1 vccd1 vccd1 _08762_/A sky130_fd_sc_hd__or2_1
XFILLER_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07128__A1 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _08675_/B _08675_/C _08675_/D _08971_/B vssd1 vssd1 vccd1 vccd1 _08674_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07625_ _14129_/Q _14064_/Q vssd1 vssd1 vccd1 vccd1 _07626_/B sky130_fd_sc_hd__or2_1
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12866__A _12920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07556_ _14103_/Q input20/X _07560_/S vssd1 vssd1 vccd1 vccd1 _07557_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07487_ _07333_/S _14194_/Q _07528_/A vssd1 vssd1 vccd1 vccd1 _07487_/X sky130_fd_sc_hd__a21o_1
XFILLER_10_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09226_ _09225_/B _09225_/C _09225_/A vssd1 vssd1 vccd1 vccd1 _09227_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__13385__A0 _12654_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13697__A _13731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14008__D _14008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09157_ _09151_/A _09151_/B _09151_/C vssd1 vssd1 vccd1 vccd1 _09158_/C sky130_fd_sc_hd__a21o_1
X_08108_ _08750_/B vssd1 vssd1 vccd1 vccd1 _08791_/B sky130_fd_sc_hd__buf_2
XANTENNA__07064__B1 _07048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09088_ _09088_/A _10092_/A vssd1 vssd1 vccd1 vccd1 _09090_/B sky130_fd_sc_hd__nor2_1
X_08039_ _08039_/A _08039_/B vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__nor2_2
XANTENNA__12106__A _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11050_ _11050_/A _11050_/B vssd1 vssd1 vccd1 vccd1 _11129_/B sky130_fd_sc_hd__xnor2_1
XFILLER_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11163__A2 _10912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10001_ _09998_/Y _09999_/Y _10000_/Y vssd1 vssd1 vccd1 vccd1 _10420_/B sky130_fd_sc_hd__a21oi_4
XFILLER_103_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11945__A _11947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11952_ _11953_/A vssd1 vssd1 vccd1 vccd1 _11952_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09134__B _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06878__B1 _06877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _10903_/A vssd1 vssd1 vccd1 vccd1 _13929_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11883_ _13750_/Q _11883_/B vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__and2_1
XFILLER_72_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13622_ _13625_/A _13622_/B vssd1 vssd1 vccd1 vccd1 _13623_/A sky130_fd_sc_hd__and2_1
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10834_ _10834_/A _10834_/B vssd1 vssd1 vccd1 vccd1 _10835_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ _13556_/A _13553_/B vssd1 vssd1 vccd1 vccd1 _13554_/A sky130_fd_sc_hd__and2_1
X_10765_ _10765_/A _10765_/B _11186_/S _10757_/B vssd1 vssd1 vccd1 vccd1 _10765_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12504_ _14005_/Q _12460_/A _12503_/X _12498_/X vssd1 vssd1 vccd1 vccd1 _14005_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13484_ input92/X _14392_/Q _13494_/S vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__mux2_1
X_10696_ _11240_/A vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ _12450_/A vssd1 vssd1 vccd1 vccd1 _12435_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12366_ _12366_/A vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14105_ _14107_/CLK _14105_/D _12756_/Y vssd1 vssd1 vccd1 vccd1 _14105_/Q sky130_fd_sc_hd__dfrtp_4
X_11317_ _11317_/A _11317_/B _11317_/C vssd1 vssd1 vccd1 vccd1 _11317_/X sky130_fd_sc_hd__or3_1
XFILLER_10_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12297_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12297_/Y sky130_fd_sc_hd__inv_2
X_14036_ _14054_/CLK _14036_/D vssd1 vssd1 vccd1 vccd1 _14036_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_45_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11248_ _11252_/B _11253_/A _11020_/A vssd1 vssd1 vccd1 vccd1 _11249_/B sky130_fd_sc_hd__a21o_1
XFILLER_45_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13546__S _13559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11855__A _11855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11179_ _11249_/A _11253_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__nand3b_1
XFILLER_67_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09044__B _09188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07410_ _07464_/A vssd1 vssd1 vccd1 vccd1 _07431_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08390_ _09698_/A _09698_/B _09698_/C vssd1 vssd1 vccd1 vccd1 _08390_/Y sky130_fd_sc_hd__nor3_1
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_25_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07341_ _07321_/X _07337_/X _07340_/X _07329_/X vssd1 vssd1 vccd1 vccd1 _07341_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07272_ _07312_/A vssd1 vssd1 vccd1 vccd1 _07308_/A sky130_fd_sc_hd__inv_2
X_09011_ _09152_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _09015_/A sky130_fd_sc_hd__nand2_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12590__A1 _14030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09913_ _10271_/B _09913_/B vssd1 vssd1 vccd1 vccd1 _09914_/B sky130_fd_sc_hd__and2_1
XFILLER_113_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11765__A input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09844_ _09844_/A _09844_/B vssd1 vssd1 vccd1 vccd1 _09844_/X sky130_fd_sc_hd__and2_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09775_ _08273_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _09775_/X sky130_fd_sc_hd__and2b_1
XFILLER_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06987_ _14261_/Q _06968_/X _06986_/X hold33/X vssd1 vssd1 vccd1 vccd1 _06987_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08726_ _08726_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _08727_/B sky130_fd_sc_hd__nand2_1
XFILLER_96_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_73_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14250_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08657_ _08656_/B _08656_/C _08656_/A vssd1 vssd1 vccd1 vccd1 _08665_/B sky130_fd_sc_hd__a21o_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07608_ _07608_/A vssd1 vssd1 vccd1 vccd1 _14080_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08588_ _08643_/A _08643_/B vssd1 vssd1 vccd1 vccd1 _08619_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07539_ _14181_/Q _07526_/X _07538_/Y _14192_/D vssd1 vssd1 vccd1 vccd1 _14173_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10550_ _10629_/S vssd1 vssd1 vccd1 vccd1 _10550_/X sky130_fd_sc_hd__buf_2
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _09209_/A _09209_/B vssd1 vssd1 vccd1 vccd1 _09210_/B sky130_fd_sc_hd__nor2_2
XFILLER_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10481_ _10498_/C _10480_/B _10480_/C vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__a21o_1
X_12220_ _12218_/X _07323_/X _12220_/S vssd1 vssd1 vccd1 vccd1 _12221_/B sky130_fd_sc_hd__mux2_1
XFILLER_68_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12151_ _12904_/A _12160_/B vssd1 vssd1 vccd1 vccd1 _12151_/X sky130_fd_sc_hd__or2_1
XFILLER_29_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11102_ _11102_/A _11102_/B _11105_/B vssd1 vssd1 vccd1 vccd1 _11102_/X sky130_fd_sc_hd__or3_1
X_12082_ _12082_/A vssd1 vssd1 vccd1 vccd1 _13805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11136__A2 _11110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11033_ _11134_/B _10963_/B _10963_/C _11262_/A vssd1 vssd1 vccd1 vccd1 _11039_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09145__A _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12984_ _12985_/A vssd1 vssd1 vccd1 vccd1 _12984_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10647__A1 _13952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ _11935_/A vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__buf_2
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _14353_/Q _11870_/B vssd1 vssd1 vccd1 vccd1 _11867_/A sky130_fd_sc_hd__and2_1
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13597__A0 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13605_ _13605_/A vssd1 vssd1 vccd1 vccd1 _14426_/D sky130_fd_sc_hd__clkbuf_1
X_10817_ _10846_/B _10846_/C _10846_/A vssd1 vssd1 vccd1 vccd1 _10840_/B sky130_fd_sc_hd__a21oi_1
X_11797_ _11797_/A vssd1 vssd1 vccd1 vccd1 _11797_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13536_ _13539_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13537_/A sky130_fd_sc_hd__and2_1
X_10748_ _10748_/A _10748_/B vssd1 vssd1 vccd1 vccd1 _10748_/X sky130_fd_sc_hd__and2_1
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13467_ input90/X _14387_/Q _13467_/S vssd1 vssd1 vccd1 vccd1 _13468_/B sky130_fd_sc_hd__mux2_1
X_10679_ _10679_/A vssd1 vssd1 vccd1 vccd1 _10967_/S sky130_fd_sc_hd__buf_2
XFILLER_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12418_ _12722_/A vssd1 vssd1 vccd1 vccd1 _12703_/A sky130_fd_sc_hd__clkbuf_4
X_13398_ _13398_/A vssd1 vssd1 vccd1 vccd1 _14366_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12572__A1 _14025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12349_ _12353_/A vssd1 vssd1 vccd1 vccd1 _12349_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06910_ _07027_/A vssd1 vssd1 vccd1 vccd1 _06942_/B sky130_fd_sc_hd__clkbuf_4
X_14019_ _14020_/CLK _14019_/D vssd1 vssd1 vccd1 vccd1 _14019_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07890_ _07890_/A _07890_/B vssd1 vssd1 vccd1 vccd1 _07890_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09055__A _09055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09560_ _09560_/A _09560_/B _09560_/C vssd1 vssd1 vccd1 vccd1 _09563_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08894__A _09055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08511_ _14014_/Q vssd1 vssd1 vccd1 vccd1 _09457_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09491_ _09491_/A _09792_/A vssd1 vssd1 vccd1 vccd1 _09491_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08442_ _09869_/A vssd1 vssd1 vccd1 vccd1 _09882_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07303__A _07471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08373_ _09824_/A vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__buf_4
X_07324_ _14107_/Q _07323_/X vssd1 vssd1 vccd1 vccd1 _07324_/X sky130_fd_sc_hd__or2b_1
XFILLER_104_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07255_ _14077_/Q _13877_/Q _07258_/S vssd1 vssd1 vccd1 vccd1 _07255_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07186_ _07186_/A vssd1 vssd1 vccd1 vccd1 _07186_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09827_ _10271_/A _09926_/B vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__nor2_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09758_ _09771_/A _08264_/B _08263_/A vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__o21a_1
XFILLER_104_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08709_ _08709_/A _08760_/A vssd1 vssd1 vccd1 vccd1 _08723_/A sky130_fd_sc_hd__nand2_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09689_ _09607_/B _09675_/Y _09687_/Y _09688_/X vssd1 vssd1 vccd1 vccd1 _09692_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11717_/Y _11718_/X _11719_/Y vssd1 vssd1 vccd1 vccd1 _11720_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08309__A _13868_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11651_/A _11651_/B vssd1 vssd1 vccd1 vccd1 _11651_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_70_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07258__A0 _14076_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ _10627_/A _10621_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10613_/A sky130_fd_sc_hd__and3_1
XFILLER_74_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14370_ _14417_/CLK _14370_/D vssd1 vssd1 vccd1 vccd1 _14370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11582_ _14056_/Q _13968_/Q vssd1 vssd1 vccd1 vccd1 _11587_/A sky130_fd_sc_hd__and2_1
XFILLER_70_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12773__B _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13321_ _14426_/Q _13306_/X _13319_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13321_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10533_ _13966_/Q _10532_/X _10585_/S vssd1 vssd1 vccd1 vccd1 _10534_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ _14411_/Q _13230_/X _13251_/X vssd1 vssd1 vccd1 vccd1 _13252_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input74_A io_wbs_datwr[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ _10302_/A _09969_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _10465_/A sky130_fd_sc_hd__a21bo_1
X_12203_ _12203_/A vssd1 vssd1 vccd1 vccd1 _12203_/X sky130_fd_sc_hd__clkbuf_2
X_13183_ _13183_/A vssd1 vssd1 vccd1 vccd1 _13183_/Y sky130_fd_sc_hd__inv_2
X_10395_ _10395_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _10426_/B sky130_fd_sc_hd__xnor2_2
XFILLER_97_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _12147_/A vssd1 vssd1 vccd1 vccd1 _12143_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08698__B _09457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12065_ _12065_/A _12065_/B vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__and2_1
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11016_ _11244_/A _11016_/B vssd1 vssd1 vccd1 vccd1 _11017_/B sky130_fd_sc_hd__and2_1
XFILLER_49_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07733__A1 _14158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11817__B1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12967_ _12973_/A vssd1 vssd1 vccd1 vccd1 _12972_/A sky130_fd_sc_hd__buf_2
XFILLER_18_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06946__B _14284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11918_ _13761_/Q _11703_/B _11917_/X vssd1 vssd1 vccd1 vccd1 _11919_/B sky130_fd_sc_hd__a21oi_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12898_ _12942_/A _12898_/B vssd1 vssd1 vccd1 vccd1 _12898_/X sky130_fd_sc_hd__or2_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11849_ _14342_/Q _11847_/X _11848_/X _13801_/Q vssd1 vssd1 vccd1 vccd1 _11849_/X
+ sky130_fd_sc_hd__a22o_2
XANTENNA__09238__A1 _09127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__A0 _14079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13519_ _13519_/A vssd1 vssd1 vccd1 vccd1 _14402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07040_ _14416_/Q _07039_/Y _07009_/X vssd1 vssd1 vccd1 vccd1 _07040_/X sky130_fd_sc_hd__a21o_1
XFILLER_115_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08889__A _09241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08991_ _08991_/A _08991_/B _08991_/C vssd1 vssd1 vccd1 vccd1 _08993_/B sky130_fd_sc_hd__nand3_2
XFILLER_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07942_ _13869_/Q vssd1 vssd1 vccd1 vccd1 _09818_/B sky130_fd_sc_hd__buf_2
XFILLER_87_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07873_ _07873_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07873_/X sky130_fd_sc_hd__xor2_1
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09612_ _09612_/A vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07017__B _14275_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09543_ _09543_/A _09543_/B _09543_/C _09543_/D vssd1 vssd1 vccd1 vccd1 _09593_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10659__A _11322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09474_ _09424_/B _09843_/A _09863_/A _09424_/A vssd1 vssd1 vccd1 vccd1 _09475_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08425_ _13864_/Q vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12874__A _12917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08356_ _09153_/B _08976_/A _09058_/B _08623_/A vssd1 vssd1 vccd1 vccd1 _08360_/A
+ sky130_fd_sc_hd__a22oi_1
X_07307_ _07307_/A _07307_/B _07307_/C vssd1 vssd1 vccd1 vccd1 _07319_/A sky130_fd_sc_hd__or3_1
X_08287_ _09596_/A _08287_/B _08287_/C vssd1 vssd1 vccd1 vccd1 _08376_/A sky130_fd_sc_hd__or3_1
XFILLER_109_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14365__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ _07258_/S vssd1 vssd1 vccd1 vccd1 _07252_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_106_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11002__B _11002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07169_ _14102_/Q _07167_/X _07168_/X vssd1 vssd1 vccd1 vccd1 _07169_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10180_ _10180_/A _10180_/B vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12114__A _13731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10631__B_N _10644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13870_ _13946_/CLK _13870_/D _12271_/Y vssd1 vssd1 vccd1 vccd1 _13870_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_74_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12821_ hold37/A _12772_/X _12803_/A _14148_/Q _12809_/A vssd1 vssd1 vccd1 vccd1
+ _12821_/X sky130_fd_sc_hd__a221o_1
XFILLER_41_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _12752_/A vssd1 vssd1 vccd1 vccd1 _12752_/Y sky130_fd_sc_hd__inv_2
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _13761_/Q _11703_/B vssd1 vssd1 vccd1 vccd1 _11920_/C sky130_fd_sc_hd__or2_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12696_/A _12683_/B vssd1 vssd1 vccd1 vccd1 _12684_/A sky130_fd_sc_hd__and2_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _14452_/CLK _14422_/D vssd1 vssd1 vccd1 vccd1 _14422_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12224__B1 _13193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ _11634_/A _11634_/B _11634_/C vssd1 vssd1 vccd1 vccd1 _11634_/X sky130_fd_sc_hd__or3_1
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14353_ _14464_/CLK _14353_/D vssd1 vssd1 vccd1 vccd1 _14353_/Q sky130_fd_sc_hd__dfxtp_1
X_11565_ _11545_/Y _11627_/A _11626_/B vssd1 vssd1 vccd1 vccd1 _11623_/A sky130_fd_sc_hd__o21a_2
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _14422_/Q _13284_/X _13303_/X _13299_/X vssd1 vssd1 vccd1 vccd1 _13304_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10516_ _09750_/Y _10512_/X _10515_/Y vssd1 vssd1 vccd1 vccd1 _10516_/Y sky130_fd_sc_hd__a21oi_4
X_14284_ _14284_/CLK _14284_/D _13146_/Y vssd1 vssd1 vccd1 vccd1 _14284_/Q sky130_fd_sc_hd__dfrtp_4
X_11496_ _08815_/B _11486_/X _11494_/X _11495_/X vssd1 vssd1 vccd1 vccd1 _13868_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12527__A1 _08896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13235_ _14440_/Q _13201_/X _13204_/X _14392_/Q vssd1 vssd1 vccd1 vccd1 _13235_/X
+ sky130_fd_sc_hd__a22o_1
X_10447_ _10493_/A _10447_/B vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10538__B1 _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ _13178_/A vssd1 vssd1 vccd1 vccd1 _13171_/A sky130_fd_sc_hd__buf_2
X_10378_ _10378_/A _10378_/B _10378_/C vssd1 vssd1 vccd1 vccd1 _10564_/B sky130_fd_sc_hd__and3_1
XANTENNA__11750__A2 hold16/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ _12146_/A vssd1 vssd1 vccd1 vccd1 _12117_/X sky130_fd_sc_hd__clkbuf_2
X_13097_ _13106_/A _13097_/B vssd1 vssd1 vccd1 vccd1 _13098_/A sky130_fd_sc_hd__and2_1
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12048_ _13428_/A vssd1 vssd1 vccd1 vccd1 _12536_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13999_ _14396_/CLK _13999_/D vssd1 vssd1 vccd1 vccd1 _13999_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12463__B1 _12462_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14388__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08210_ _09762_/A _09800_/A _09963_/B _08249_/A vssd1 vssd1 vccd1 vccd1 _08211_/B
+ sky130_fd_sc_hd__a22o_1
X_09190_ _09049_/A _09188_/X _09187_/X _09189_/X vssd1 vssd1 vccd1 vccd1 _09190_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_92_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12766__A1 _14149_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12766__B2 _14133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08141_ _08141_/A _08203_/C vssd1 vssd1 vccd1 vccd1 _08205_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08434__A2 _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _08150_/A _08150_/B _08071_/X vssd1 vssd1 vccd1 vccd1 _08073_/B sky130_fd_sc_hd__a21bo_1
XFILLER_88_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13715__A0 input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07023_ _07023_/A vssd1 vssd1 vccd1 vccd1 _14307_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09508__A _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08974_ _09041_/A _08974_/B vssd1 vssd1 vccd1 vccd1 _09029_/A sky130_fd_sc_hd__xnor2_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09147__B1 _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07925_ _14023_/Q vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__buf_2
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11773__A input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13464__S _13467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07856_ _07872_/A _07873_/A _07855_/Y vssd1 vssd1 vccd1 vccd1 _07869_/A sky130_fd_sc_hd__o21ai_1
XFILLER_60_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09243__A _09319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07787_ _07806_/B vssd1 vssd1 vccd1 vccd1 _10664_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_83_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13246__A2 _13336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ _09518_/Y _09519_/X _09454_/Y _09470_/X vssd1 vssd1 vccd1 vccd1 _09527_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09457_ _09457_/A _09457_/B _13874_/Q _09457_/D vssd1 vssd1 vccd1 vccd1 _09459_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_12_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08408_ _09749_/B _08240_/X _08239_/X _08193_/A vssd1 vssd1 vccd1 vccd1 _08409_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09388_ _09388_/A _09388_/B vssd1 vssd1 vccd1 vccd1 _09423_/B sky130_fd_sc_hd__xnor2_2
X_08339_ _08336_/A _08337_/Y _08194_/X _08338_/Y vssd1 vssd1 vccd1 vccd1 _09751_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12109__A _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ _11350_/A _11350_/B vssd1 vssd1 vccd1 vccd1 _11351_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12509__A1 _12209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10301_ _10048_/A _10279_/B _10282_/A vssd1 vssd1 vccd1 vccd1 _10302_/B sky130_fd_sc_hd__a21oi_2
XFILLER_119_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11948__A _11971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ _11338_/A _11342_/A _11339_/A vssd1 vssd1 vccd1 vccd1 _11336_/C sky130_fd_sc_hd__o21bai_1
XFILLER_106_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13020_ _13022_/A vssd1 vssd1 vccd1 vccd1 _13020_/Y sky130_fd_sc_hd__inv_2
X_10232_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10233_/B sky130_fd_sc_hd__xor2_1
XFILLER_106_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09925__A2 _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10163_ _10164_/A _10164_/B vssd1 vssd1 vccd1 vccd1 _10182_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input37_A io_wbs_adr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10094_ _10333_/B _10101_/A vssd1 vssd1 vccd1 vccd1 _10095_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11496__A1 _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13922_ _13927_/CLK _13922_/D _12335_/Y vssd1 vssd1 vccd1 vccd1 _13922_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_48_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09153__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13853_ _13892_/CLK _13853_/D _12248_/Y vssd1 vssd1 vccd1 vccd1 _13853_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13237__A2 _13236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ _14157_/Q _12801_/X _12803_/X _14141_/Q _12791_/X vssd1 vssd1 vccd1 vccd1
+ _12804_/X sky130_fd_sc_hd__a221o_2
X_10996_ _10999_/B _11000_/A _11220_/A vssd1 vssd1 vccd1 vccd1 _10997_/B sky130_fd_sc_hd__a21o_1
X_13784_ _13809_/CLK _13784_/D vssd1 vssd1 vccd1 vccd1 _13784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12735_ _12753_/A vssd1 vssd1 vccd1 vccd1 _12740_/A sky130_fd_sc_hd__buf_2
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12678_/A _12666_/B vssd1 vssd1 vccd1 vccd1 _12667_/A sky130_fd_sc_hd__and2_1
X_14405_ _14451_/CLK _14405_/D vssd1 vssd1 vccd1 vccd1 _14405_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11617_ _11617_/A vssd1 vssd1 vccd1 vccd1 _13850_/D sky130_fd_sc_hd__clkbuf_1
X_12597_ _12924_/A _14032_/Q _12600_/S vssd1 vssd1 vccd1 vccd1 _12598_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11420__A1 _11056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07120__B _07134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14336_ _14400_/CLK _14336_/D vssd1 vssd1 vccd1 vccd1 _14336_/Q sky130_fd_sc_hd__dfxtp_1
X_11548_ _14044_/Q _13956_/Q vssd1 vssd1 vccd1 vccd1 _11548_/X sky130_fd_sc_hd__or2_1
XFILLER_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13549__S _13559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14267_ _14275_/CLK _14267_/D _13126_/Y vssd1 vssd1 vccd1 vccd1 _14267_/Q sky130_fd_sc_hd__dfrtp_4
X_11479_ _11471_/A _11478_/X _10686_/X vssd1 vssd1 vccd1 vccd1 _11479_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13218_ _13245_/A vssd1 vssd1 vccd1 vccd1 _13218_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11184__A0 _11142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ _14198_/CLK _14198_/D _12989_/Y vssd1 vssd1 vccd1 vccd1 _14198_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__08232__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13152_/A vssd1 vssd1 vccd1 vccd1 _13149_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07710_ _07765_/S vssd1 vssd1 vccd1 vccd1 _07730_/S sky130_fd_sc_hd__buf_2
X_08690_ _08967_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _08964_/B sky130_fd_sc_hd__xnor2_2
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07641_ _07669_/A _07670_/A _07640_/Y vssd1 vssd1 vccd1 vccd1 _07667_/A sky130_fd_sc_hd__o21a_2
XFILLER_66_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06902__A2 _06873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09998__A _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07572_ _07572_/A vssd1 vssd1 vccd1 vccd1 _14096_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10002__A _10420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09311_ _09349_/A _09543_/C vssd1 vssd1 vccd1 vccd1 _09313_/B sky130_fd_sc_hd__and2_1
XANTENNA__09852__A1 _10127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09242_ _09242_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09173_ _09173_/A _09173_/B _09173_/C vssd1 vssd1 vccd1 vccd1 _09175_/A sky130_fd_sc_hd__and3_1
XFILLER_119_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07615__A0 _14076_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08124_ _08124_/A _08124_/B vssd1 vssd1 vccd1 vccd1 _08144_/B sky130_fd_sc_hd__and2_1
XANTENNA__11411__A1 _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08055_ _14022_/Q vssd1 vssd1 vccd1 vccd1 _09472_/B sky130_fd_sc_hd__clkbuf_2
X_07006_ _07006_/A vssd1 vssd1 vccd1 vccd1 _14309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_32_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_89_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07981__A _14019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08957_ _08957_/A _08957_/B vssd1 vssd1 vccd1 vccd1 _08957_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08796__B _08796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14468__180 vssd1 vssd1 vccd1 vccd1 _14468__180/HI io_oeb[0] sky130_fd_sc_hd__conb_1
X_07908_ _14027_/Q _13973_/Q vssd1 vssd1 vccd1 vccd1 _07909_/B sky130_fd_sc_hd__nand2_1
X_08888_ _08978_/B vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_99_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07839_ _07840_/A _07839_/B _07909_/A _07839_/D vssd1 vssd1 vccd1 vccd1 _07840_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13219__A2 _13336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10850_ _11100_/A vssd1 vssd1 vccd1 vccd1 _10851_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_60_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09509_ _09510_/B _09510_/C _08098_/X vssd1 vssd1 vccd1 vccd1 _09511_/B sky130_fd_sc_hd__a21bo_1
XFILLER_24_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _13930_/Q _10788_/B vssd1 vssd1 vccd1 vccd1 _10889_/B sky130_fd_sc_hd__and2_1
XFILLER_40_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12909_/A _08946_/A _12520_/S vssd1 vssd1 vccd1 vccd1 _12521_/B sky130_fd_sc_hd__mux2_1
XFILLER_40_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08317__A _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07221__A _07258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12451_ _12473_/A vssd1 vssd1 vccd1 vccd1 _12451_/X sky130_fd_sc_hd__clkbuf_2
X_11402_ _13879_/Q _11392_/X _11396_/X _11401_/X vssd1 vssd1 vccd1 vccd1 _13879_/D
+ sky130_fd_sc_hd__a22o_1
X_12382_ _12384_/A vssd1 vssd1 vccd1 vccd1 _12382_/Y sky130_fd_sc_hd__inv_2
X_14121_ _14239_/CLK _14121_/D vssd1 vssd1 vccd1 vccd1 _14121_/Q sky130_fd_sc_hd__dfxtp_1
X_11333_ _11333_/A _11333_/B _11333_/C vssd1 vssd1 vccd1 vccd1 _11334_/B sky130_fd_sc_hd__nand3_1
XFILLER_4_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14052_ _14367_/CLK _14052_/D vssd1 vssd1 vccd1 vccd1 _14052_/Q sky130_fd_sc_hd__dfxtp_2
X_11264_ _11264_/A _11264_/B _11264_/C vssd1 vssd1 vccd1 vccd1 _11268_/A sky130_fd_sc_hd__or3_1
XFILLER_106_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13003_ _13003_/A vssd1 vssd1 vccd1 vccd1 _13003_/Y sky130_fd_sc_hd__inv_2
X_10215_ _10215_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__nand2_1
XFILLER_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11195_ _10650_/A _11172_/X _11143_/A vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__o21ai_2
XFILLER_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10146_ _10146_/A _10144_/A vssd1 vssd1 vccd1 vccd1 _10146_/X sky130_fd_sc_hd__or2b_1
XFILLER_39_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output143_A _11825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11469__A1 _11082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10078_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12302__A _12304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13905_ _13905_/CLK _13905_/D _12314_/Y vssd1 vssd1 vccd1 vccd1 _13905_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_78_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07542__C1 _14192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ _14259_/CLK _13836_/D vssd1 vssd1 vccd1 vccd1 _13836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10979_ _10651_/A _10951_/B _10920_/A vssd1 vssd1 vccd1 vccd1 _11008_/A sky130_fd_sc_hd__o21ai_2
X_13767_ _13820_/CLK _13767_/D _11959_/Y vssd1 vssd1 vccd1 vccd1 _13767_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06954__B _14283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13950_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12718_ _12721_/A vssd1 vssd1 vccd1 vccd1 _12718_/Y sky130_fd_sc_hd__inv_2
X_13698_ input74/X _14453_/Q _13704_/S vssd1 vssd1 vccd1 vccd1 _13699_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12649_ _12649_/A vssd1 vssd1 vccd1 vccd1 _14045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06970__A _06970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07073__A1 _14268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14319_ _14322_/CLK _14319_/D _13189_/Y vssd1 vssd1 vccd1 vccd1 _14319_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09058__A _09234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _10186_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09966_/C sky130_fd_sc_hd__nand2_1
XFILLER_97_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08811_ _08811_/A _08811_/B _08811_/C vssd1 vssd1 vccd1 vccd1 _08811_/Y sky130_fd_sc_hd__nand3_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09791_ _10367_/A vssd1 vssd1 vccd1 vccd1 _10346_/A sky130_fd_sc_hd__clkbuf_2
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _08742_/A _08803_/A vssd1 vssd1 vccd1 vccd1 _08743_/B sky130_fd_sc_hd__nor2_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_io_wbs_clk clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14410_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08673_ _08670_/X _08669_/X _08668_/X _08970_/A vssd1 vssd1 vccd1 vccd1 _08971_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07624_ _14129_/Q _14064_/Q vssd1 vssd1 vccd1 vccd1 _07626_/A sky130_fd_sc_hd__nand2_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07555_ _07555_/A vssd1 vssd1 vccd1 vccd1 _14104_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08628__A2 _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07486_ _14076_/Q _11746_/S _07460_/A _13876_/Q _07471_/X vssd1 vssd1 vccd1 vccd1
+ _07486_/X sky130_fd_sc_hd__a221o_1
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09225_ _09225_/A _09225_/B _09225_/C vssd1 vssd1 vccd1 vccd1 _09227_/A sky130_fd_sc_hd__and3_1
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13385__A1 _14363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09156_ _09156_/A _09156_/B vssd1 vssd1 vccd1 vccd1 _09158_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07976__A _14020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08107_ _14013_/Q vssd1 vssd1 vccd1 vccd1 _08750_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09087_ _09087_/A _09087_/B _09087_/C vssd1 vssd1 vccd1 vccd1 _09090_/A sky130_fd_sc_hd__nand3_1
XFILLER_107_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08038_ _08580_/A _08555_/B _09508_/C vssd1 vssd1 vccd1 vccd1 _08039_/B sky130_fd_sc_hd__o21ai_1
XFILLER_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11010__B _11010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10000_ _10000_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _10000_/Y sky130_fd_sc_hd__nor2_2
XFILLER_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09989_ _10269_/A _10269_/B vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__xnor2_2
XFILLER_118_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13218__A _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12122__A input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07119__A2 _07085_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11951_ _11953_/A vssd1 vssd1 vccd1 vccd1 _11951_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10902_ _13929_/Q _10901_/X _10902_/S vssd1 vssd1 vccd1 vccd1 _10903_/A sky130_fd_sc_hd__mux2_1
X_11882_ _11882_/A vssd1 vssd1 vccd1 vccd1 _11882_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13621_ input85/X _14431_/Q _13628_/S vssd1 vssd1 vccd1 vccd1 _13622_/B sky130_fd_sc_hd__mux2_1
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13073__A0 _12515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ _10831_/X _10828_/C _10832_/Y _10675_/X _13942_/Q vssd1 vssd1 vccd1 vccd1
+ _13942_/D sky130_fd_sc_hd__a32o_1
XFILLER_83_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13552_ input95/X _14411_/Q _13559_/S vssd1 vssd1 vccd1 vccd1 _13553_/B sky130_fd_sc_hd__mux2_1
X_10764_ _13933_/Q _10797_/B vssd1 vssd1 vccd1 vccd1 _10873_/B sky130_fd_sc_hd__and2_1
XANTENNA__14449__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ _14056_/Q _12442_/X _12435_/X vssd1 vssd1 vccd1 vccd1 _12503_/X sky130_fd_sc_hd__a21o_1
X_13483_ _12911_/A _13475_/S _13482_/Y vssd1 vssd1 vccd1 vccd1 _14391_/D sky130_fd_sc_hd__o21a_1
X_10695_ _11020_/A vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__buf_2
XFILLER_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12434_ _13209_/A _13111_/C vssd1 vssd1 vccd1 vccd1 _12450_/A sky130_fd_sc_hd__nand2_1
X_12365_ _12366_/A vssd1 vssd1 vccd1 vccd1 _12365_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14104_ _14104_/CLK _14104_/D _12755_/Y vssd1 vssd1 vccd1 vccd1 _14104_/Q sky130_fd_sc_hd__dfrtp_4
X_11316_ _11119_/X _11312_/B _11315_/Y _10851_/B _11302_/A vssd1 vssd1 vccd1 vccd1
+ _13908_/D sky130_fd_sc_hd__a32o_1
XFILLER_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12296_/Y sky130_fd_sc_hd__inv_2
X_14035_ _14367_/CLK _14035_/D vssd1 vssd1 vccd1 vccd1 _14035_/Q sky130_fd_sc_hd__dfxtp_4
X_11247_ _13898_/Q vssd1 vssd1 vccd1 vccd1 _11273_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11178_ _11256_/A _11262_/C _11258_/A vssd1 vssd1 vccd1 vccd1 _11252_/B sky130_fd_sc_hd__and3_1
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10129_ _10307_/B _10129_/B vssd1 vssd1 vccd1 vccd1 _10129_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09341__A _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13819_ _13820_/CLK _13819_/D vssd1 vssd1 vccd1 vccd1 _13819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10487__A _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07340_ _14220_/Q _14222_/Q _07360_/S vssd1 vssd1 vccd1 vccd1 _07340_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12811__B1 _12810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07271_ _14178_/Q _14177_/Q _07520_/B vssd1 vssd1 vccd1 vccd1 _07312_/A sky130_fd_sc_hd__or3_2
X_09010_ _09010_/A _08627_/B vssd1 vssd1 vccd1 vccd1 _09071_/A sky130_fd_sc_hd__or2b_1
XFILLER_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12207__A _12216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09912_ _09912_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__xnor2_4
XFILLER_99_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09843_ _09843_/A _09863_/A vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__or2_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08420__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06986_ _14405_/Q _06985_/Y _06970_/X vssd1 vssd1 vccd1 vccd1 _06986_/X sky130_fd_sc_hd__a21o_1
X_09774_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09779_/A sky130_fd_sc_hd__xnor2_1
X_08725_ _08966_/A _10009_/A _08734_/B _08724_/Y vssd1 vssd1 vccd1 vccd1 _08779_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_73_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _08656_/A _08656_/B _08656_/C vssd1 vssd1 vccd1 vccd1 _08665_/A sky130_fd_sc_hd__nand3_2
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _14080_/Q input27/X _07615_/S vssd1 vssd1 vccd1 vccd1 _07608_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _08587_/A _08587_/B vssd1 vssd1 vccd1 vccd1 _08643_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07538_ _07543_/B _07538_/B vssd1 vssd1 vccd1 vccd1 _07538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07469_ _14196_/Q _14198_/Q _07469_/S vssd1 vssd1 vccd1 vccd1 _07470_/B sky130_fd_sc_hd__mux2_1
X_09208_ _08623_/B _08629_/A _09882_/A _08623_/A vssd1 vssd1 vccd1 vccd1 _09209_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_10_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ _10498_/C _10480_/B _10480_/C vssd1 vssd1 vccd1 vccd1 _10520_/A sky130_fd_sc_hd__nand3_1
XANTENNA__11908__A2 _11906_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07037__A1 _14305_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ _09137_/A _09137_/C _09137_/B vssd1 vssd1 vccd1 vccd1 _09140_/C sky130_fd_sc_hd__a21o_1
XFILLER_68_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12117__A _12146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12150_ input66/X vssd1 vssd1 vccd1 vccd1 _12904_/A sky130_fd_sc_hd__buf_6
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11101_ _10831_/X _11097_/C _11099_/Y _11100_/X _11079_/A vssd1 vssd1 vccd1 vccd1
+ _13924_/D sky130_fd_sc_hd__a32o_1
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13647__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _12081_/A _12081_/B vssd1 vssd1 vccd1 vccd1 _12082_/A sky130_fd_sc_hd__and2_1
X_11032_ _11032_/A vssd1 vssd1 vccd1 vccd1 _11052_/A sky130_fd_sc_hd__inv_2
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09145__B _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12983_ _12985_/A vssd1 vssd1 vccd1 vccd1 _12983_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11844__A1 _14340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ _12223_/A vssd1 vssd1 vccd1 vccd1 _11935_/A sky130_fd_sc_hd__buf_4
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11844__B2 _13799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11865_/A vssd1 vssd1 vccd1 vccd1 _11865_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _13607_/A _13604_/B vssd1 vssd1 vccd1 vccd1 _13605_/A sky130_fd_sc_hd__and2_1
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10816_ _10840_/A _10815_/X vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__or2b_1
X_11796_ _12440_/A vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13535_ input88/X _14406_/Q _13542_/S vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__mux2_1
XFILLER_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10747_ _13936_/Q _10806_/B vssd1 vssd1 vccd1 vccd1 _10858_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13411__A _13411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10678_ _10944_/S vssd1 vssd1 vccd1 vccd1 _10679_/A sky130_fd_sc_hd__buf_2
XANTENNA__09017__A2 _08925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13466_ _13466_/A vssd1 vssd1 vccd1 vccd1 _14386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12417_ _13010_/A vssd1 vssd1 vccd1 vccd1 _12722_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_2_2_0_io_wbs_clk_A clkbuf_2_3_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_86_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13397_ _13409_/A _13397_/B vssd1 vssd1 vccd1 vccd1 _13398_/A sky130_fd_sc_hd__and2_1
X_12348_ _12348_/A vssd1 vssd1 vccd1 vccd1 _12353_/A sky130_fd_sc_hd__buf_2
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12279_ _12279_/A vssd1 vssd1 vccd1 vccd1 _12279_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14018_ _14020_/CLK _14018_/D vssd1 vssd1 vccd1 vccd1 _14018_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09336__A _09336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07200__A1 _14093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09055__B _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08894__B _08941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08510_ _08823_/A _09361_/D _09092_/D _08595_/A vssd1 vssd1 vccd1 vccd1 _08693_/C
+ sky130_fd_sc_hd__a22oi_2
X_09490_ _09152_/A _09848_/A _09433_/B _09431_/X vssd1 vssd1 vccd1 vccd1 _09496_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_63_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08441_ _08750_/B vssd1 vssd1 vccd1 vccd1 _09508_/B sky130_fd_sc_hd__buf_4
XFILLER_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08372_ _09234_/B vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__buf_4
XFILLER_17_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12796__C1 _12216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07323_ _07363_/A vssd1 vssd1 vccd1 vccd1 _07323_/X sky130_fd_sc_hd__buf_2
XFILLER_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07254_ _07254_/A vssd1 vssd1 vccd1 vccd1 _14262_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08415__A _09044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07019__A1 _14275_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ _07185_/A vssd1 vssd1 vccd1 vccd1 _07185_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13467__S _13467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08150__A _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ _09826_/A _09826_/B vssd1 vssd1 vccd1 vccd1 _09926_/B sky130_fd_sc_hd__and2_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09757_ _09757_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__xnor2_1
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06969_ _14457_/Q _14281_/Q vssd1 vssd1 vccd1 vccd1 _06969_/Y sky130_fd_sc_hd__nand2_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _08709_/A _08708_/B _08708_/C vssd1 vssd1 vccd1 vccd1 _08760_/A sky130_fd_sc_hd__nand3_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09687_/A _09687_/C _09687_/B vssd1 vssd1 vccd1 vccd1 _09688_/X sky130_fd_sc_hd__o21a_1
XFILLER_64_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08639_/A _08639_/B _08639_/C vssd1 vssd1 vccd1 vccd1 _08641_/A sky130_fd_sc_hd__and3_1
XFILLER_14_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11016__A _11244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11650_/A _11650_/B vssd1 vssd1 vccd1 vccd1 _11651_/A sky130_fd_sc_hd__nor2_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10601_ _10644_/B _09117_/Y _10632_/A vssd1 vssd1 vccd1 vccd1 _10627_/A sky130_fd_sc_hd__a21oi_2
X_11581_ _11591_/A _11592_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11587_/C sky130_fd_sc_hd__a21boi_1
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13320_ _13341_/A vssd1 vssd1 vccd1 vccd1 _13320_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10532_ _10528_/X _10524_/B _10530_/Y _10531_/Y _10520_/B vssd1 vssd1 vccd1 vccd1
+ _10532_/X sky130_fd_sc_hd__a32o_1
XFILLER_7_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13251_ _14443_/Q _13250_/X _13245_/X _14395_/Q vssd1 vssd1 vccd1 vccd1 _13251_/X
+ sky130_fd_sc_hd__a22o_1
X_10463_ _10436_/B _09766_/A _10463_/S vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12202_ _12200_/X _12202_/B _12202_/C vssd1 vssd1 vccd1 vccd1 _12202_/Y sky130_fd_sc_hd__nand3b_1
X_13182_ _13183_/A vssd1 vssd1 vccd1 vccd1 _13182_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input67_A io_wbs_datwr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ _10394_/A _10394_/B vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__xor2_1
XFILLER_11_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12133_ _12146_/A vssd1 vssd1 vccd1 vccd1 _12133_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08698__C _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12064_ _13800_/Q _12059_/X _12060_/X hold17/A vssd1 vssd1 vccd1 vccd1 _12065_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11015_ _13918_/Q vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_78_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12966_ _12966_/A vssd1 vssd1 vccd1 vccd1 _12966_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11817__B2 _14114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07404__A _11746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11917_ _13821_/Q _13762_/Q _11920_/C vssd1 vssd1 vccd1 vccd1 _11917_/X sky130_fd_sc_hd__o21ba_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12490__A1 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _14147_/Q _12885_/X _12896_/X _12892_/X vssd1 vssd1 vccd1 vccd1 _14147_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12490__B2 _14052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11848_ _11848_/A vssd1 vssd1 vccd1 vccd1 _11848_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14017__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09238__A2 _09127_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12778__C1 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11779_ _12193_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12192_/A sky130_fd_sc_hd__and2_1
XFILLER_53_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13518_ _13518_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13519_/A sky130_fd_sc_hd__and2_1
X_13449_ _13461_/A _13449_/B vssd1 vssd1 vccd1 vccd1 _13450_/A sky130_fd_sc_hd__and2_1
XFILLER_86_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08990_ _08989_/A _08989_/B _08989_/C vssd1 vssd1 vccd1 vccd1 _08991_/C sky130_fd_sc_hd__a21o_1
XFILLER_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07941_ _09424_/B vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__buf_4
XFILLER_69_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_37_io_wbs_clk_A clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07872_ _07872_/A _07855_/Y vssd1 vssd1 vccd1 vccd1 _07873_/B sky130_fd_sc_hd__or2b_1
XFILLER_60_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09611_ _09708_/A _09612_/A _09708_/C vssd1 vssd1 vccd1 vccd1 _09611_/X sky130_fd_sc_hd__and3_1
XFILLER_110_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09542_ _09481_/B _09483_/B _09481_/A vssd1 vssd1 vccd1 vccd1 _09548_/A sky130_fd_sc_hd__o21ba_1
XFILLER_110_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09473_ _14021_/Q _09473_/B vssd1 vssd1 vccd1 vccd1 _09475_/B sky130_fd_sc_hd__and2_1
X_08424_ _09881_/B vssd1 vssd1 vccd1 vccd1 _09152_/B sky130_fd_sc_hd__buf_2
XFILLER_12_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08355_ _09286_/A vssd1 vssd1 vccd1 vccd1 _08623_/A sky130_fd_sc_hd__clkbuf_4
X_07306_ _07306_/A vssd1 vssd1 vccd1 vccd1 _14225_/D sky130_fd_sc_hd__clkbuf_1
X_08286_ _08716_/A _10000_/A _08208_/C _08632_/A vssd1 vssd1 vccd1 vccd1 _08287_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07237_ _07237_/A vssd1 vssd1 vccd1 vccd1 _14267_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07984__A _08012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ _07186_/A vssd1 vssd1 vccd1 vccd1 _07168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07099_ _07090_/X _07098_/X _14361_/Q vssd1 vssd1 vccd1 vccd1 _07100_/S sky130_fd_sc_hd__o21a_1
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09809_ _10123_/A vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06923__B1 _06877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13988__RESET_B _12419_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ _14122_/Q _12771_/X _12819_/X _12817_/X vssd1 vssd1 vccd1 vccd1 _14122_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12130__A input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12472__A1 _08716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12751_ _12752_/A vssd1 vssd1 vccd1 vccd1 _12751_/Y sky130_fd_sc_hd__inv_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13660__S _13670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11702_ _13760_/Q _11914_/B vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__or2_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12682_ _12681_/X _14053_/Q _12685_/S vssd1 vssd1 vccd1 vccd1 _12683_/B sky130_fd_sc_hd__mux2_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _14452_/CLK _14421_/D vssd1 vssd1 vccd1 vccd1 _14421_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11633_/A vssd1 vssd1 vccd1 vccd1 _13846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14352_ _14354_/CLK _14352_/D vssd1 vssd1 vccd1 vccd1 _14352_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12775__A2 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11564_ _14047_/Q _13959_/Q vssd1 vssd1 vccd1 vccd1 _11626_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08055__A _14022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13303_ _14374_/Q _13215_/A _13294_/X _14454_/Q vssd1 vssd1 vccd1 vccd1 _13303_/X
+ sky130_fd_sc_hd__a22o_1
X_10515_ _10614_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10515_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11495_ _11010_/B _11489_/X _11475_/X _11288_/A _11490_/X vssd1 vssd1 vccd1 vccd1
+ _11495_/X sky130_fd_sc_hd__o221a_1
XFILLER_100_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14283_ _14283_/CLK _14283_/D _13145_/Y vssd1 vssd1 vccd1 vccd1 _14283_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13234_ _14327_/Q _13196_/X _13233_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _14327_/D
+ sky130_fd_sc_hd__o211a_1
X_10446_ _10446_/A _10446_/B vssd1 vssd1 vccd1 vccd1 _10447_/B sky130_fd_sc_hd__nor2_1
XANTENNA_output173_A _14298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13165_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13165_/Y sky130_fd_sc_hd__inv_2
X_10377_ _10377_/A _10377_/B vssd1 vssd1 vccd1 vccd1 _10378_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12305__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12116_ _13811_/Q _12095_/X _12112_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _13811_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13488__A0 _12645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13096_ _12641_/X hold20/A _13096_/S vssd1 vssd1 vccd1 vccd1 _13097_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12047_ _13609_/A vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08903__A1 _09044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13998_ _14442_/CLK _13998_/D vssd1 vssd1 vccd1 vccd1 _13998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12949_ _12950_/A vssd1 vssd1 vccd1 vccd1 _12949_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13660__A0 input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06973__A _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08891__C _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12215__A1 _11990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08140_ _08140_/A _08140_/B vssd1 vssd1 vccd1 vccd1 _08203_/C sky130_fd_sc_hd__nor2_1
XFILLER_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08071_ _08547_/A _08284_/C _09834_/A _08573_/A vssd1 vssd1 vccd1 vccd1 _08071_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07300__C _14166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07022_ _07019_/X _14307_/Q _07022_/S vssd1 vssd1 vccd1 vccd1 _07023_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12923__C1 _12920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__B _09508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13479__A0 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ _08973_/A _08973_/B vssd1 vssd1 vccd1 vccd1 _08974_/B sky130_fd_sc_hd__xor2_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_07924_ _09788_/A vssd1 vssd1 vccd1 vccd1 _07924_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09524__A _09584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ _14036_/Q _13982_/Q vssd1 vssd1 vccd1 vccd1 _07855_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07786_ _07786_/A vssd1 vssd1 vccd1 vccd1 _11452_/B sky130_fd_sc_hd__buf_2
XFILLER_72_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09525_ _09629_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09527_/B sky130_fd_sc_hd__xor2_1
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07979__A _14020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ _09388_/A _09386_/X _09387_/A vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__a21o_1
XFILLER_101_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08407_ _09751_/C _08407_/B _08407_/C vssd1 vssd1 vccd1 vccd1 _10524_/A sky130_fd_sc_hd__or3_2
XFILLER_24_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09387_ _09387_/A _09386_/X vssd1 vssd1 vccd1 vccd1 _09388_/B sky130_fd_sc_hd__or2b_1
XFILLER_71_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08338_ _08194_/A _08194_/B _08194_/C vssd1 vssd1 vccd1 vccd1 _08338_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ _09634_/A _08270_/B vssd1 vssd1 vccd1 vccd1 _08271_/A sky130_fd_sc_hd__or2_1
X_10300_ _10278_/A _10278_/B _10273_/X vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__a21o_1
X_11280_ _11336_/B _11280_/B vssd1 vssd1 vccd1 vccd1 _11339_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08603__A _09132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _10194_/A _10200_/A _10195_/B _10195_/A vssd1 vssd1 vccd1 vccd1 _10231_/Y
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_69_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10162_ _10162_/A _10162_/B vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10093_ _10083_/A _10083_/B _10092_/X vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13921_ _13927_/CLK _13921_/D _12334_/Y vssd1 vssd1 vccd1 vccd1 _13921_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11175__S _11175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13852_ _13892_/CLK _13852_/D _12247_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09153__B _09153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12803_ _12803_/A vssd1 vssd1 vccd1 vccd1 _12803_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13783_ _14258_/CLK _13783_/D vssd1 vssd1 vccd1 vccd1 _13783_/Q sky130_fd_sc_hd__dfxtp_1
X_10995_ _13923_/Q vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13988_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12734_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12734_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12664_/X _14049_/Q _12665_/S vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__mux2_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _14440_/CLK _14404_/D vssd1 vssd1 vccd1 vccd1 _14404_/Q sky130_fd_sc_hd__dfxtp_1
X_11616_ _13850_/Q _11614_/Y _11632_/S vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__A2_N _08658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ _12637_/A vssd1 vssd1 vccd1 vccd1 _12615_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14335_ _14335_/CLK _14335_/D vssd1 vssd1 vccd1 vccd1 _14335_/Q sky130_fd_sc_hd__dfxtp_1
X_11547_ _14045_/Q _13957_/Q vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14266_ _14365_/CLK _14266_/D _13125_/Y vssd1 vssd1 vccd1 vccd1 _14266_/Q sky130_fd_sc_hd__dfrtp_2
X_11478_ _11478_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__and2_1
XANTENNA__11708__B1 hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13217_ _13637_/A vssd1 vssd1 vccd1 vccd1 _13336_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_48_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10429_ _10429_/A vssd1 vssd1 vccd1 vccd1 _10429_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14197_ _14198_/CLK _14197_/D _12988_/Y vssd1 vssd1 vccd1 vccd1 _14197_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _13152_/A vssd1 vssd1 vccd1 vccd1 _13148_/Y sky130_fd_sc_hd__inv_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13079_ _13079_/A _13079_/B vssd1 vssd1 vccd1 vccd1 _13105_/S sky130_fd_sc_hd__or2_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_io_wbs_clk clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14335_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07640_ _14131_/Q _14066_/Q vssd1 vssd1 vccd1 vccd1 _07640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07560__A0 _14101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07571_ _14096_/Q input13/X _07571_/S vssd1 vssd1 vccd1 vccd1 _07572_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09310_ _09508_/A _09508_/B _09792_/B _09553_/D vssd1 vssd1 vccd1 vccd1 _09313_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_34_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09241_ _09241_/A _09241_/B _09545_/D _09241_/D vssd1 vssd1 vccd1 vccd1 _09242_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07949__D _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09172_ _09171_/A _09171_/C _09171_/B vssd1 vssd1 vccd1 vccd1 _09173_/C sky130_fd_sc_hd__a21o_1
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _08076_/B _08076_/C _08076_/A vssd1 vssd1 vccd1 vccd1 _08160_/B sky130_fd_sc_hd__a21oi_1
XFILLER_119_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08054_ _08054_/A _08054_/B vssd1 vssd1 vccd1 vccd1 _08076_/C sky130_fd_sc_hd__nand2_1
XFILLER_31_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08423__A _13865_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07005_ _07002_/X _14309_/Q _07005_/S vssd1 vssd1 vccd1 vccd1 _07006_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08040__A1 _08716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08956_ _08952_/X _08954_/Y _08924_/B _08924_/A _08955_/X vssd1 vssd1 vccd1 vccd1
+ _08956_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_9_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07907_ _13951_/D _07921_/C _07840_/B _07905_/X _07906_/X vssd1 vssd1 vccd1 vccd1
+ _13974_/D sky130_fd_sc_hd__a41o_1
X_08887_ _08887_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _08887_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_99_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07838_ _14027_/Q _13973_/Q _07909_/C vssd1 vssd1 vccd1 vccd1 _07839_/D sky130_fd_sc_hd__a21o_1
XFILLER_99_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13624__A0 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ _07203_/A _14226_/Q _07769_/S vssd1 vssd1 vccd1 vccd1 _07769_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13504__A _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ _09508_/A _09508_/B _09508_/C _09545_/D vssd1 vssd1 vccd1 vccd1 _09510_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_13_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10780_ _10780_/A _10780_/B vssd1 vssd1 vccd1 vccd1 _10788_/B sky130_fd_sc_hd__xnor2_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09373_/B _09373_/C _09373_/A vssd1 vssd1 vccd1 vccd1 _09440_/C sky130_fd_sc_hd__a21bo_1
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08317__B _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12450_ _12450_/A vssd1 vssd1 vccd1 vccd1 _12473_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11401_ hold30/X _11403_/B vssd1 vssd1 vccd1 vccd1 _11401_/X sky130_fd_sc_hd__or2_1
X_12381_ _12384_/A vssd1 vssd1 vccd1 vccd1 _12381_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14120_ _14163_/CLK _14120_/D vssd1 vssd1 vccd1 vccd1 _14120_/Q sky130_fd_sc_hd__dfxtp_1
X_11332_ _11288_/A _11319_/X _11331_/Y _11322_/X vssd1 vssd1 vccd1 vccd1 _13903_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14228__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14051_ _14367_/CLK _14051_/D vssd1 vssd1 vccd1 vccd1 _14051_/Q sky130_fd_sc_hd__dfxtp_1
X_11263_ _11264_/A _11264_/B _11264_/C vssd1 vssd1 vccd1 vccd1 _11350_/A sky130_fd_sc_hd__nor3_1
XFILLER_107_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13002_ _13003_/A vssd1 vssd1 vccd1 vccd1 _13002_/Y sky130_fd_sc_hd__inv_2
X_10214_ _10214_/A _10214_/B vssd1 vssd1 vccd1 vccd1 _10214_/Y sky130_fd_sc_hd__nand2_1
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11194_ _10650_/A _11164_/X _11143_/A vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__o21ai_4
XFILLER_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10145_ _10151_/B vssd1 vssd1 vccd1 vccd1 _10145_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09164__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10076_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13904_ _13949_/CLK _13904_/D _12313_/Y vssd1 vssd1 vccd1 vccd1 _13904_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10677__B1 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13835_ _14441_/CLK _13835_/D vssd1 vssd1 vccd1 vccd1 _13835_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13615__A0 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13766_ _13825_/CLK _13766_/D _11958_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10978_ _10650_/A _10943_/X _10920_/A vssd1 vssd1 vccd1 vccd1 _11012_/A sky130_fd_sc_hd__o21ai_2
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12717_ _12721_/A vssd1 vssd1 vccd1 vccd1 _12717_/Y sky130_fd_sc_hd__inv_2
X_13697_ _13731_/A vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07131__B _14279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12648_ _12656_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _12649_/A sky130_fd_sc_hd__and2_1
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12579_ input91/X vssd1 vssd1 vccd1 vccd1 _12579_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14318_ _14322_/CLK _14318_/D _13188_/Y vssd1 vssd1 vccd1 vccd1 _14318_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__10601__B1 _10632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14249_ _14250_/CLK _14249_/D vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfxtp_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _08810_/A _08815_/C vssd1 vssd1 vccd1 vccd1 _08811_/C sky130_fd_sc_hd__xnor2_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _13969_/Q _07924_/X _09783_/X _09789_/Y vssd1 vssd1 vccd1 vccd1 _13969_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09074__A _09297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08741_ _08779_/A _08779_/B _08740_/Y vssd1 vssd1 vccd1 vccd1 _09038_/B sky130_fd_sc_hd__o21ai_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10668__B1 _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ _08672_/A vssd1 vssd1 vccd1 vccd1 _08675_/D sky130_fd_sc_hd__inv_2
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07623_ _14130_/Q _14065_/Q vssd1 vssd1 vccd1 vccd1 _07671_/B sky130_fd_sc_hd__or2_1
XFILLER_4_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13606__A0 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07554_ _14104_/Q input21/X _07560_/S vssd1 vssd1 vccd1 vccd1 _07555_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07485_ _07348_/A _07483_/X _07484_/X _07373_/A _14194_/Q vssd1 vssd1 vccd1 vccd1
+ _14194_/D sky130_fd_sc_hd__a32o_1
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09224_ _09223_/A _09223_/C _09223_/B vssd1 vssd1 vccd1 vccd1 _09225_/C sky130_fd_sc_hd__a21o_1
XFILLER_50_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09155_ _09155_/A _09155_/B vssd1 vssd1 vccd1 vccd1 _09156_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12593__A0 _12922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08106_ _14014_/Q vssd1 vssd1 vccd1 vccd1 _08595_/A sky130_fd_sc_hd__buf_2
X_09086_ _09472_/B _09941_/A _09941_/B _09472_/A vssd1 vssd1 vccd1 vccd1 _09087_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08037_ _08097_/B vssd1 vssd1 vccd1 vccd1 _09508_/C sky130_fd_sc_hd__buf_2
XFILLER_66_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07992__A _09800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09988_ _10268_/A _10268_/B vssd1 vssd1 vccd1 vccd1 _10269_/B sky130_fd_sc_hd__xor2_2
XFILLER_89_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08939_ _08939_/A _08939_/B vssd1 vssd1 vccd1 vccd1 _08940_/B sky130_fd_sc_hd__and2_1
XFILLER_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11950_ _11953_/A vssd1 vssd1 vccd1 vccd1 _11950_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07524__B1 _07528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09712__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ _10836_/S _10894_/B _10899_/Y _10900_/X vssd1 vssd1 vccd1 vccd1 _10901_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ hold40/X _11872_/X _11879_/X _11880_/Y _11874_/X vssd1 vssd1 vccd1 vccd1
+ _13749_/D sky130_fd_sc_hd__o221a_1
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11453__S _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13620_ _13620_/A vssd1 vssd1 vccd1 vccd1 _14430_/D sky130_fd_sc_hd__clkbuf_1
X_10832_ _10832_/A _10832_/B vssd1 vssd1 vccd1 vccd1 _10832_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13551_ _13551_/A vssd1 vssd1 vccd1 vccd1 _14410_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10763_ _11020_/A _10773_/A _10763_/S vssd1 vssd1 vccd1 vccd1 _10797_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12502_ _14004_/Q _12460_/A _12501_/X _12498_/X vssd1 vssd1 vccd1 vccd1 _14004_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13482_ _06880_/Y _13475_/S _11935_/A vssd1 vssd1 vccd1 vccd1 _13482_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_input97_A io_wbs_datwr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10694_ _11252_/A vssd1 vssd1 vccd1 vccd1 _11020_/A sky130_fd_sc_hd__buf_2
X_12433_ _12624_/A _12952_/B vssd1 vssd1 vccd1 vccd1 _13111_/C sky130_fd_sc_hd__nor2_2
XFILLER_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _12366_/A vssd1 vssd1 vccd1 vccd1 _12364_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14103_ _14107_/CLK _14103_/D _12754_/Y vssd1 vssd1 vccd1 vccd1 _14103_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_114_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11315_ _11315_/A _11315_/B _11315_/C vssd1 vssd1 vccd1 vccd1 _11315_/Y sky130_fd_sc_hd__nand3_1
X_12295_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12295_/Y sky130_fd_sc_hd__inv_2
X_14034_ _14367_/CLK _14034_/D vssd1 vssd1 vccd1 vccd1 _14034_/Q sky130_fd_sc_hd__dfxtp_4
X_11246_ _11276_/A _11276_/B vssd1 vssd1 vccd1 vccd1 _11338_/A sky130_fd_sc_hd__and2_1
XFILLER_84_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11177_ _10769_/A _11172_/X _11173_/X _10744_/X _11176_/X vssd1 vssd1 vccd1 vccd1
+ _11258_/A sky130_fd_sc_hd__a221oi_4
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10128_ _10307_/B _10129_/B vssd1 vssd1 vccd1 vccd1 _10135_/B sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_4_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14217_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_76_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10059_ _10059_/A _10080_/A vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07515__A0 hold34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13144__A _13146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13818_ _13825_/CLK _13818_/D vssd1 vssd1 vccd1 vccd1 _13818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08238__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13749_ _14335_/CLK _13749_/D _11937_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09060__C _09060_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07270_ _14176_/Q _14175_/Q _07534_/A vssd1 vssd1 vccd1 vccd1 _07520_/B sky130_fd_sc_hd__or3_1
XFILLER_31_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12575__A0 _12909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09911_ _10124_/B _10157_/A vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_0_io_wbs_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_59_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _09842_/A _09857_/B vssd1 vssd1 vccd1 vccd1 _10127_/A sky130_fd_sc_hd__xnor2_4
XFILLER_101_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12223__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__xnor2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _14437_/Q _14261_/Q vssd1 vssd1 vccd1 vccd1 _06985_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08724_ _08723_/B _08729_/B _08722_/B vssd1 vssd1 vccd1 vccd1 _08724_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _08654_/B _08654_/C _08654_/A vssd1 vssd1 vccd1 vccd1 _08656_/C sky130_fd_sc_hd__o21ai_1
XFILLER_82_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07606_ _14256_/Q vssd1 vssd1 vccd1 vccd1 _07615_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _08586_/A _08585_/X vssd1 vssd1 vccd1 vccd1 _08587_/B sky130_fd_sc_hd__or2b_1
XFILLER_23_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08148__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07537_ _14173_/Q _07541_/A vssd1 vssd1 vccd1 vccd1 _07538_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07809__A1 _07784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07987__A _09553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ _07452_/X _07466_/X _07467_/X _07462_/X _14198_/Q vssd1 vssd1 vccd1 vccd1
+ _14198_/D sky130_fd_sc_hd__a32o_1
X_09207_ _09286_/A _09286_/B _09207_/C _09869_/A vssd1 vssd1 vccd1 vccd1 _09209_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_44_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_33_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07399_ _07399_/A vssd1 vssd1 vccd1 vccd1 _07399_/X sky130_fd_sc_hd__buf_2
X_09138_ _09081_/A _09081_/C _09081_/B vssd1 vssd1 vccd1 vccd1 _09140_/B sky130_fd_sc_hd__a21bo_1
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09069_ _08991_/B _08993_/B _09119_/A _09068_/Y vssd1 vssd1 vccd1 vccd1 _09119_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_68_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11100_ _11100_/A vssd1 vssd1 vccd1 vccd1 _11100_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12080_ _13805_/Q _12000_/A _12021_/A _13821_/Q vssd1 vssd1 vccd1 vccd1 _12081_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _13914_/Q vssd1 vssd1 vccd1 vccd1 _11032_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12133__A _12146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12982_ _12985_/A vssd1 vssd1 vccd1 vccd1 _12982_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input12_A dout1[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14416__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _13153_/A vssd1 vssd1 vccd1 vccd1 _12223_/A sky130_fd_sc_hd__buf_4
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11864_ _14352_/Q _11864_/B vssd1 vssd1 vccd1 vccd1 _11865_/A sky130_fd_sc_hd__and2_1
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08058__A _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ input80/X _14426_/Q _13611_/S vssd1 vssd1 vccd1 vccd1 _13604_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _10705_/B _10727_/C _10727_/D _13939_/Q vssd1 vssd1 vccd1 vccd1 _10815_/X
+ sky130_fd_sc_hd__a31o_1
X_11795_ _11855_/A vssd1 vssd1 vccd1 vccd1 _11870_/B sky130_fd_sc_hd__buf_4
XFILLER_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13534_ _13534_/A vssd1 vssd1 vccd1 vccd1 _14405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08208__D _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10746_ _10746_/A _10746_/B vssd1 vssd1 vccd1 vccd1 _10806_/B sky130_fd_sc_hd__xor2_1
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13349__A2 _13216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13465_ _13485_/A _13465_/B vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__and2_1
X_10677_ _10669_/X _10670_/Y _10761_/C _10675_/X _11186_/S vssd1 vssd1 vccd1 vccd1
+ _13948_/D sky130_fd_sc_hd__a32o_1
XFILLER_12_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12416_ input98/X vssd1 vssd1 vccd1 vccd1 _13010_/A sky130_fd_sc_hd__buf_2
XFILLER_51_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ _12668_/X _14366_/Q _13408_/S vssd1 vssd1 vccd1 vccd1 _13397_/B sky130_fd_sc_hd__mux2_1
XFILLER_86_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12347_ _12347_/A vssd1 vssd1 vccd1 vccd1 _12347_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11866__B _11870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12278_ _12279_/A vssd1 vssd1 vccd1 vccd1 _12278_/Y sky130_fd_sc_hd__inv_2
X_14017_ _14020_/CLK _14017_/D vssd1 vssd1 vccd1 vccd1 _14017_/Q sky130_fd_sc_hd__dfxtp_2
X_11229_ _11229_/A _11229_/B vssd1 vssd1 vccd1 vccd1 _11288_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__11532__A1 _08937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11882__A _11882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08440_ _08982_/A _08794_/B vssd1 vssd1 vccd1 vccd1 _08503_/B sky130_fd_sc_hd__and2_1
XFILLER_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _08842_/A _09786_/A _09595_/B _08370_/X vssd1 vssd1 vccd1 vccd1 _08385_/A
+ sky130_fd_sc_hd__a31o_2
XANTENNA__11599__A1 _11598_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07322_ _13836_/Q vssd1 vssd1 vccd1 vccd1 _07363_/A sky130_fd_sc_hd__buf_2
XANTENNA__09661__B1 _09414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10945__B _13895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07253_ _14262_/Q _07252_/X _07253_/S vssd1 vssd1 vccd1 vccd1 _07254_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12218__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07184_ _07184_/A vssd1 vssd1 vccd1 vccd1 _14282_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09964__A1 _08980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11523__A1 _11032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input4_A dout1[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _10037_/A vssd1 vssd1 vccd1 vccd1 _10271_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09756_ _09769_/A _08255_/B _09755_/X vssd1 vssd1 vccd1 vccd1 _09757_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06886__A _13778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ _06968_/A vssd1 vssd1 vccd1 vccd1 _06968_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08707_ _08707_/A _08707_/B vssd1 vssd1 vccd1 vccd1 _08708_/C sky130_fd_sc_hd__xnor2_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09687_ _09687_/A _09687_/B _09687_/C vssd1 vssd1 vccd1 vccd1 _09687_/Y sky130_fd_sc_hd__nor3_4
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06899_ _06899_/A vssd1 vssd1 vccd1 vccd1 _14323_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _08998_/B _08636_/C _08636_/A vssd1 vssd1 vccd1 vccd1 _08639_/C sky130_fd_sc_hd__a21o_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08569_ _08863_/D vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__buf_4
XFILLER_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10600_ _10597_/X _10599_/X _13958_/Q _10545_/X vssd1 vssd1 vccd1 vccd1 _13958_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_11580_ _14055_/Q _13967_/Q vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10531_ _10482_/Y _10458_/X _10461_/X _10462_/X _10528_/X vssd1 vssd1 vccd1 vccd1
+ _10531_/Y sky130_fd_sc_hd__a41oi_1
XFILLER_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12128__A input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11032__A _11032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13250_ _13637_/A vssd1 vssd1 vccd1 vccd1 _13250_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10462_ _10450_/B _10456_/A _10450_/A vssd1 vssd1 vccd1 vccd1 _10462_/X sky130_fd_sc_hd__o21ba_1
X_12201_ _12201_/A _12205_/B _13835_/Q vssd1 vssd1 vccd1 vccd1 _12202_/B sky130_fd_sc_hd__or3b_1
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12562__S _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ _13183_/A vssd1 vssd1 vccd1 vccd1 _13181_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11762__A_N input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ _10393_/A _10413_/A vssd1 vssd1 vccd1 vccd1 _10404_/C sky130_fd_sc_hd__nand2_1
X_12132_ hold17/A _12117_/X _12130_/X _12131_/X vssd1 vssd1 vccd1 vccd1 _13816_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12063_ _12063_/A vssd1 vssd1 vccd1 vccd1 _13799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11014_ _11064_/B _11014_/B vssd1 vssd1 vccd1 vccd1 _11111_/B sky130_fd_sc_hd__and2b_1
XFILLER_93_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07194__A1 _14095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06941__A1 _14285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12965_ _12966_/A vssd1 vssd1 vccd1 vccd1 _12965_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ hold5/X _11916_/B vssd1 vssd1 vccd1 vccd1 _13760_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _12940_/A _12896_/B vssd1 vssd1 vccd1 vccd1 _12896_/X sky130_fd_sc_hd__or2_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _11870_/B vssd1 vssd1 vccd1 vccd1 _11847_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08446__A1 _09508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08446__B2 _08445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11778_ _12951_/B vssd1 vssd1 vccd1 vccd1 _12193_/B sky130_fd_sc_hd__inv_2
XFILLER_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07420__A _14227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11450__A0 _11142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13517_ _12561_/X _14402_/Q _13522_/S vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__mux2_1
X_10729_ _10729_/A vssd1 vssd1 vccd1 vccd1 _10730_/B sky130_fd_sc_hd__buf_2
XANTENNA__12038__A _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13448_ input83/X _14381_/Q _13460_/S vssd1 vssd1 vccd1 vccd1 _13449_/B sky130_fd_sc_hd__mux2_1
XFILLER_103_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13379_ _12645_/X _14361_/Q _13391_/S vssd1 vssd1 vccd1 vccd1 _13380_/B sky130_fd_sc_hd__mux2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08251__A _08251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07940_ _14022_/Q vssd1 vssd1 vccd1 vccd1 _09424_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11505__A1 _10215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_opt_2_0_io_wbs_clk clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14008_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07871_ _07871_/A vssd1 vssd1 vccd1 vccd1 _13983_/D sky130_fd_sc_hd__clkbuf_1
X_09610_ _09675_/A _09608_/Y _09586_/B _09586_/Y vssd1 vssd1 vccd1 vccd1 _09708_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09541_ _09541_/A _09541_/B vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11762__D input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09472_ _09472_/A _09472_/B _09844_/A _09844_/B vssd1 vssd1 vccd1 vccd1 _09475_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__08685__A1 _08683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08685__B2 _08767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09810__A _13867_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08423_ _13865_/Q vssd1 vssd1 vccd1 vccd1 _09881_/B sky130_fd_sc_hd__buf_2
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13332__A _13332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ _08353_/A _08353_/B _08353_/C vssd1 vssd1 vccd1 vccd1 _08363_/B sky130_fd_sc_hd__a21o_1
X_07305_ _07301_/Y _14225_/Q _07305_/S vssd1 vssd1 vccd1 vccd1 _07306_/A sky130_fd_sc_hd__mux2_1
X_08285_ _09001_/B vssd1 vssd1 vccd1 vccd1 _08716_/A sky130_fd_sc_hd__buf_6
XFILLER_20_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07236_ _14267_/Q _07235_/X _07236_/S vssd1 vssd1 vccd1 vccd1 _07237_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__C1 _09397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07167_ _07185_/A vssd1 vssd1 vccd1 vccd1 _07167_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07984__B _08573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07098_ _14409_/Q _07098_/B _14441_/Q vssd1 vssd1 vccd1 vccd1 _07098_/X sky130_fd_sc_hd__and3b_1
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13829__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07176__A1 _14100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _08794_/B _09806_/X _09807_/X vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__a21oi_4
XFILLER_28_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09739_ _09739_/A _09739_/B _09739_/C vssd1 vssd1 vccd1 vccd1 _09742_/B sky130_fd_sc_hd__and3_1
XFILLER_28_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11027__A _11056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12750_ _12752_/A vssd1 vssd1 vccd1 vccd1 _12750_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _13759_/Q _11911_/B vssd1 vssd1 vccd1 vccd1 _11914_/B sky130_fd_sc_hd__or2_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ input70/X vssd1 vssd1 vccd1 vccd1 _12681_/X sky130_fd_sc_hd__buf_4
XFILLER_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14452_/CLK _14420_/D vssd1 vssd1 vccd1 vccd1 _14420_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ hold19/A _11631_/Y _11632_/S vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14351_ _14354_/CLK _14351_/D vssd1 vssd1 vccd1 vccd1 _14351_/Q sky130_fd_sc_hd__dfxtp_1
X_11563_ _11546_/Y _11631_/A _11630_/B vssd1 vssd1 vccd1 vccd1 _11627_/A sky130_fd_sc_hd__o21a_2
XANTENNA__07100__A1 _14297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ _14341_/Q _13289_/X _13300_/X _13301_/X vssd1 vssd1 vccd1 vccd1 _14341_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ _10644_/A vssd1 vssd1 vccd1 vccd1 _10614_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14282_ _14283_/CLK _14282_/D _13144_/Y vssd1 vssd1 vccd1 vccd1 _14282_/Q sky130_fd_sc_hd__dfrtp_4
X_11494_ _11487_/A _11493_/X _11472_/X vssd1 vssd1 vccd1 vccd1 _11494_/X sky130_fd_sc_hd__a21o_1
X_13233_ _14359_/Q _13215_/X _13232_/X _13222_/X vssd1 vssd1 vccd1 vccd1 _13233_/X
+ sky130_fd_sc_hd__a211o_1
X_10445_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__nor2_1
XFILLER_100_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13164_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13164_/Y sky130_fd_sc_hd__inv_2
X_10376_ _10376_/A _10375_/X vssd1 vssd1 vccd1 vccd1 _10378_/B sky130_fd_sc_hd__or2b_1
XANTENNA_output166_A _14293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _12203_/A vssd1 vssd1 vccd1 vccd1 _12115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13488__A1 _14393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13095_ _13095_/A vssd1 vssd1 vccd1 vccd1 _14249_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12046_ _12046_/A vssd1 vssd1 vccd1 vccd1 _13609_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_43_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14427_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08903__A2 _10215_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13997_ _14440_/CLK _13997_/D vssd1 vssd1 vccd1 vccd1 _13997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07134__B _07134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12948_ _12950_/A vssd1 vssd1 vccd1 vccd1 _12948_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _12920_/A vssd1 vssd1 vccd1 vccd1 _12879_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08891__D _08925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08070_ _08126_/A _08284_/C _08070_/C vssd1 vssd1 vccd1 vccd1 _08150_/B sky130_fd_sc_hd__and3_1
XFILLER_105_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07021_ _07012_/X _07020_/X _14371_/Q vssd1 vssd1 vccd1 vccd1 _07022_/S sky130_fd_sc_hd__o21a_1
XFILLER_115_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ _08664_/A _08663_/A _08663_/B vssd1 vssd1 vccd1 vccd1 _08973_/B sky130_fd_sc_hd__o21ba_1
XFILLER_69_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07923_ _11452_/A _10664_/B _11452_/B vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__nand3b_4
XFILLER_116_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07158__A1 _14105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13327__A _13526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07854_ _07876_/A _07877_/A _07876_/B vssd1 vssd1 vccd1 vccd1 _07873_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__06905__A1 _14322_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07785_ _10655_/A vssd1 vssd1 vccd1 vccd1 _11452_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09524_ _09584_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09455_ _09455_/A _09626_/A vssd1 vssd1 vccd1 vccd1 _09468_/A sky130_fd_sc_hd__and2_1
XFILLER_101_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08406_ _08406_/A _09735_/A vssd1 vssd1 vccd1 vccd1 _08407_/C sky130_fd_sc_hd__nor2_1
XFILLER_51_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09386_ _09385_/A _09385_/C _09385_/B vssd1 vssd1 vccd1 vccd1 _09386_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10217__A1 _10067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ _08337_/A vssd1 vssd1 vccd1 vccd1 _08337_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08268_ _08245_/A _08225_/B _08224_/A vssd1 vssd1 vccd1 vccd1 _08270_/B sky130_fd_sc_hd__a21oi_1
X_07219_ _14272_/Q _07218_/X _07219_/S vssd1 vssd1 vccd1 vccd1 _07220_/A sky130_fd_sc_hd__mux2_1
X_08199_ _08243_/B _08199_/B vssd1 vssd1 vccd1 vccd1 _08201_/B sky130_fd_sc_hd__nand2_1
X_10230_ _10271_/B _10228_/X _10229_/X vssd1 vssd1 vccd1 vccd1 _10236_/B sky130_fd_sc_hd__o21a_1
X_10161_ _10175_/B _10176_/B _10160_/Y vssd1 vssd1 vccd1 vccd1 _10164_/A sky130_fd_sc_hd__a21o_1
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _10092_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__or2_1
XFILLER_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12142__A1 _13820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13920_ _13920_/CLK _13920_/D _12333_/Y vssd1 vssd1 vccd1 vccd1 _13920_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12141__A input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13851_ _13892_/CLK _13851_/D _12245_/Y vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfrtp_1
XFILLER_75_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09153__C _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12802_ _13202_/B _12196_/C _12828_/A vssd1 vssd1 vccd1 vccd1 _12803_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__11980__A _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13782_ _14451_/CLK _13782_/D _11981_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Q sky130_fd_sc_hd__dfrtp_1
X_10994_ _11079_/A _11079_/B vssd1 vssd1 vccd1 vccd1 _11097_/B sky130_fd_sc_hd__nand2_1
XFILLER_76_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12733_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ input97/X vssd1 vssd1 vccd1 vccd1 _12664_/X sky130_fd_sc_hd__buf_4
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14451_/CLK _14403_/D vssd1 vssd1 vccd1 vccd1 _14403_/Q sky130_fd_sc_hd__dfxtp_1
X_11615_ _11615_/A vssd1 vssd1 vccd1 vccd1 _11632_/S sky130_fd_sc_hd__clkbuf_2
X_12595_ _12595_/A vssd1 vssd1 vccd1 vccd1 _14031_/D sky130_fd_sc_hd__clkbuf_1
X_14334_ _14400_/CLK _14334_/D vssd1 vssd1 vccd1 vccd1 _14334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11546_ _14046_/Q _13958_/Q vssd1 vssd1 vccd1 vccd1 _11546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14265_ _14365_/CLK _14265_/D _13124_/Y vssd1 vssd1 vccd1 vccd1 _14265_/Q sky130_fd_sc_hd__dfrtp_2
X_11477_ _10486_/S _11455_/X _11473_/X _11476_/X vssd1 vssd1 vccd1 vccd1 _13872_/D
+ sky130_fd_sc_hd__a22o_1
X_13216_ _13526_/A vssd1 vssd1 vccd1 vccd1 _13216_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ _10443_/S _10428_/B vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__xnor2_1
X_14196_ _14224_/CLK _14196_/D _12987_/Y vssd1 vssd1 vccd1 vccd1 _14196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13147_/A vssd1 vssd1 vccd1 vccd1 _13152_/A sky130_fd_sc_hd__buf_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _10360_/A _10360_/B _10360_/C vssd1 vssd1 vccd1 vccd1 _10361_/A sky130_fd_sc_hd__o21a_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09129__A2 _09060_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13078_/A vssd1 vssd1 vccd1 vccd1 _14245_/D sky130_fd_sc_hd__clkbuf_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12029_ _13791_/Q _12020_/X _12021_/X hold24/A vssd1 vssd1 vccd1 vccd1 _12030_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07560__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07570_ _07570_/A vssd1 vssd1 vccd1 vccd1 _14097_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09360__A _09360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09240_ _09053_/B _08070_/C _09822_/A _09053_/A vssd1 vssd1 vccd1 vccd1 _09242_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09171_ _09171_/A _09171_/B _09171_/C vssd1 vssd1 vccd1 vccd1 _09173_/B sky130_fd_sc_hd__nand3_2
XANTENNA__13610__A _13680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08122_ _08122_/A _08122_/B _08122_/C vssd1 vssd1 vccd1 vccd1 _08122_/X sky130_fd_sc_hd__or3_2
XFILLER_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_49_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08053_ _08053_/A _08005_/A vssd1 vssd1 vccd1 vccd1 _08076_/B sky130_fd_sc_hd__or2b_1
X_07004_ _06973_/X _07003_/X _14373_/Q vssd1 vssd1 vccd1 vccd1 _07005_/S sky130_fd_sc_hd__o21a_1
XFILLER_116_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07039__B _14272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_io_wbs_clk io_wbs_clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_io_wbs_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08955_ _08935_/A _08935_/B _08952_/X _08954_/Y _08932_/A vssd1 vssd1 vccd1 vccd1
+ _08955_/X sky130_fd_sc_hd__a221o_1
XFILLER_5_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07906_ _13974_/Q _07919_/S vssd1 vssd1 vccd1 vccd1 _07906_/X sky130_fd_sc_hd__and2_1
XANTENNA__08796__D _09200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08886_ _08887_/A _08887_/B _08885_/A vssd1 vssd1 vccd1 vccd1 _08960_/B sky130_fd_sc_hd__o21ai_1
XFILLER_111_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07837_ _07914_/A _07915_/A _07836_/Y vssd1 vssd1 vccd1 vccd1 _07909_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__12896__A _12940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07768_ _13987_/Q _07786_/A _13988_/Q vssd1 vssd1 vccd1 vccd1 _11362_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__06894__A _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09507_ _08791_/B _08097_/B _09821_/B _08791_/A vssd1 vssd1 vccd1 vccd1 _09510_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07699_ _07700_/A _07700_/B _07658_/X _07698_/X vssd1 vssd1 vccd1 vccd1 _07699_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09437_/A _09437_/C _09437_/B vssd1 vssd1 vccd1 vccd1 _09440_/B sky130_fd_sc_hd__a21o_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13388__A0 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09369_ _09286_/B _09217_/D _09843_/A _09479_/A vssd1 vssd1 vccd1 vccd1 _09369_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13520__A _13609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ _13880_/Q _11392_/X _11396_/X _11399_/X vssd1 vssd1 vccd1 vccd1 _13880_/D
+ sky130_fd_sc_hd__a22o_1
X_12380_ _12384_/A vssd1 vssd1 vccd1 vccd1 _12380_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08614__A _08905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _11331_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11331_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14050_ _14367_/CLK _14050_/D vssd1 vssd1 vccd1 vccd1 _14050_/Q sky130_fd_sc_hd__dfxtp_1
X_11262_ _11262_/A _11355_/B _11262_/C vssd1 vssd1 vccd1 vccd1 _11264_/C sky130_fd_sc_hd__nor3_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13001_ _13003_/A vssd1 vssd1 vccd1 vccd1 _13001_/Y sky130_fd_sc_hd__inv_2
X_10213_ _10213_/A _10213_/B _10213_/C vssd1 vssd1 vccd1 vccd1 _10213_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__09764__C1 _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11193_ _11236_/B _11237_/A _11233_/A vssd1 vssd1 vccd1 vccd1 _11228_/B sky130_fd_sc_hd__and3_1
XANTENNA_input42_A io_wbs_adr[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _10144_/A _10146_/A vssd1 vssd1 vccd1 vccd1 _10151_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11186__S _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10075_ _10071_/X _10099_/B _10074_/X vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__a21oi_1
XFILLER_47_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_51_io_wbs_clk_A clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13903_ _13905_/CLK _13903_/D _12312_/Y vssd1 vssd1 vccd1 vccd1 _13903_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__10677__A1 _10669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10677__B2 _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13834_ _14259_/CLK _13834_/D vssd1 vssd1 vccd1 vccd1 _13834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13765_ _13825_/CLK _13765_/D _11957_/Y vssd1 vssd1 vccd1 vccd1 _13765_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _11016_/B _11017_/A vssd1 vssd1 vccd1 vccd1 _11011_/B sky130_fd_sc_hd__nor2_1
XFILLER_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12716_ _12722_/A vssd1 vssd1 vccd1 vccd1 _12721_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13696_ _13696_/A vssd1 vssd1 vccd1 vccd1 _14452_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13379__A0 _12645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12647_ _12645_/X _14045_/Q _12665_/S vssd1 vssd1 vccd1 vccd1 _12648_/B sky130_fd_sc_hd__mux2_1
XFILLER_87_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13430__A _13447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12578_ _12637_/A vssd1 vssd1 vccd1 vccd1 _12594_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10601__A1 _10644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11529_ _11529_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14317_ _14322_/CLK _14317_/D _13187_/Y vssd1 vssd1 vccd1 vccd1 _14317_/Q sky130_fd_sc_hd__dfrtp_4
X_14248_ _14250_/CLK _14248_/D vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11885__A _11920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14179_ _14179_/CLK _14179_/D _12965_/Y vssd1 vssd1 vccd1 vccd1 _14179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07230__A0 _14269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _08740_/A _08740_/B vssd1 vssd1 vccd1 vccd1 _08740_/Y sky130_fd_sc_hd__nand2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09074__B _09074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10668__A1 _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08671_ _08970_/A _08668_/X _08669_/X _08670_/X vssd1 vssd1 vccd1 vccd1 _08672_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07622_ _14131_/Q _14066_/Q vssd1 vssd1 vccd1 vccd1 _07669_/A sky130_fd_sc_hd__nor2_1
XFILLER_81_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07553_ _07553_/A vssd1 vssd1 vccd1 vccd1 _14105_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11125__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07390__B_N _07363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07484_ _14077_/Q _11746_/S _07460_/A _13877_/Q _07471_/X vssd1 vssd1 vccd1 vccd1
+ _07484_/X sky130_fd_sc_hd__a221o_1
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08137__C _08621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09223_ _09223_/A _09223_/B _09223_/C vssd1 vssd1 vccd1 vccd1 _09225_/B sky130_fd_sc_hd__nand3_1
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07049__B1 _07048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ _08573_/B _08449_/C _09011_/B _08012_/A vssd1 vssd1 vccd1 vccd1 _09155_/B
+ sky130_fd_sc_hd__a22oi_1
X_08105_ _09234_/A vssd1 vssd1 vccd1 vccd1 _08435_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12593__A1 _14031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09085_ _09362_/A _09085_/B vssd1 vssd1 vccd1 vccd1 _09087_/B sky130_fd_sc_hd__and2_1
X_08036_ _08579_/A vssd1 vssd1 vccd1 vccd1 _08555_/B sky130_fd_sc_hd__clkbuf_2
Xinput90 io_wbs_datwr[31] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13542__A0 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08549__B1 _08783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11795__A _11855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09987_ _09900_/A _09985_/X _09986_/X vssd1 vssd1 vccd1 vccd1 _10268_/B sky130_fd_sc_hd__o21ai_2
XFILLER_67_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08938_ _14008_/Q _08941_/B _08941_/C vssd1 vssd1 vccd1 vccd1 _08949_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08869_ _08869_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08897_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10900_ _13971_/Q _10900_/B vssd1 vssd1 vccd1 vccd1 _10900_/X sky130_fd_sc_hd__and2_1
XANTENNA__13058__C1 _13053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ _11883_/B vssd1 vssd1 vccd1 vccd1 _11880_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10831_ _11119_/A vssd1 vssd1 vccd1 vccd1 _10831_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13550_ _13556_/A _13550_/B vssd1 vssd1 vccd1 vccd1 _13551_/A sky130_fd_sc_hd__and2_1
XFILLER_73_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10762_ _10757_/X _10735_/X _10761_/X _10748_/X vssd1 vssd1 vccd1 vccd1 _10763_/S
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12501_ _14039_/Q _12485_/X _12500_/X _12473_/A vssd1 vssd1 vccd1 vccd1 _12501_/X
+ sky130_fd_sc_hd__a211o_1
X_13481_ _13481_/A vssd1 vssd1 vccd1 vccd1 _14390_/D sky130_fd_sc_hd__clkbuf_1
X_10693_ _11262_/A vssd1 vssd1 vccd1 vccd1 _11252_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13250__A _13637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12432_ _08966_/A _12486_/A _12485_/A _14024_/Q _12431_/X vssd1 vssd1 vccd1 vccd1
+ _12432_/X sky130_fd_sc_hd__a221o_1
XFILLER_8_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _12366_/A vssd1 vssd1 vccd1 vccd1 _12363_/Y sky130_fd_sc_hd__inv_2
X_14102_ _14102_/CLK _14102_/D _12752_/Y vssd1 vssd1 vccd1 vccd1 _14102_/Q sky130_fd_sc_hd__dfrtp_2
X_11314_ _07784_/X _11312_/X _11313_/Y _10904_/X _11457_/A vssd1 vssd1 vccd1 vccd1
+ _13909_/D sky130_fd_sc_hd__o32a_1
XFILLER_5_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12294_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12294_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14033_ _14367_/CLK _14033_/D vssd1 vssd1 vccd1 vccd1 _14033_/Q sky130_fd_sc_hd__dfxtp_4
X_11245_ _11245_/A _11245_/B vssd1 vssd1 vccd1 vccd1 _11276_/B sky130_fd_sc_hd__xnor2_2
XFILLER_45_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09752__A2 _10524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ _10722_/B _11174_/X _11175_/X _10730_/B vssd1 vssd1 vccd1 vccd1 _11176_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10127_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10307_/B sky130_fd_sc_hd__xnor2_4
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10058_ _10065_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__nor2_1
XFILLER_76_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08519__A _08980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13817_ _13820_/CLK _13817_/D vssd1 vssd1 vccd1 vccd1 _13817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13748_ _14335_/CLK _13748_/D _11936_/Y vssd1 vssd1 vccd1 vccd1 _13748_/Q sky130_fd_sc_hd__dfrtp_1
X_13679_ _13679_/A vssd1 vssd1 vccd1 vccd1 _14447_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13160__A _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12575__A1 _14026_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09910_ _09975_/B vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__buf_2
XFILLER_63_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09085__A _09362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09841_ _09968_/A _10463_/S vssd1 vssd1 vccd1 vccd1 _09959_/A sky130_fd_sc_hd__xnor2_2
XFILLER_113_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09772_ _09772_/A _09772_/B vssd1 vssd1 vccd1 vccd1 _09773_/B sky130_fd_sc_hd__xnor2_1
XFILLER_112_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ _06984_/A vssd1 vssd1 vccd1 vccd1 _14312_/D sky130_fd_sc_hd__clkbuf_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08723_/A _08723_/B _08723_/C vssd1 vssd1 vccd1 vccd1 _08729_/B sky130_fd_sc_hd__nand3_1
XFILLER_113_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08654_ _08654_/A _08654_/B _08654_/C vssd1 vssd1 vccd1 vccd1 _08656_/B sky130_fd_sc_hd__or3_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08429__A _13864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07605_ _07605_/A vssd1 vssd1 vccd1 vccd1 _14081_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _08637_/B _08584_/C _08584_/A vssd1 vssd1 vccd1 vccd1 _08585_/X sky130_fd_sc_hd__a21o_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07536_ _14172_/Q _14171_/Q vssd1 vssd1 vccd1 vccd1 _07541_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07809__A2 _11510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07467_ _14081_/Q _07459_/X _07460_/X _13881_/Q _07444_/X vssd1 vssd1 vccd1 vccd1
+ _07467_/X sky130_fd_sc_hd__a221o_1
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14368__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09206_ _09553_/C _09206_/B vssd1 vssd1 vccd1 vccd1 _09210_/A sky130_fd_sc_hd__nand2_2
XFILLER_72_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07398_ _14210_/Q _07373_/X _07375_/X _07397_/X vssd1 vssd1 vccd1 vccd1 _14210_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08164__A _09590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12566__A1 _12942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09137_ _09137_/A _09137_/B _09137_/C vssd1 vssd1 vccd1 vccd1 _09140_/A sky130_fd_sc_hd__nand3_1
XFILLER_5_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09068_ _09067_/B _09067_/C _09067_/A vssd1 vssd1 vccd1 vccd1 _09068_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_118_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08019_ _08020_/B _08078_/B _08131_/A vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09552__A1_N _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11030_ _11054_/A _11054_/B vssd1 vssd1 vccd1 vccd1 _11122_/B sky130_fd_sc_hd__and2_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07745__A1 _14155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11829__B1 _11823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ _12985_/A vssd1 vssd1 vccd1 vccd1 _12981_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13245__A _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11932_ input98/X vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__buf_4
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11863_ _11863_/A vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _13602_/A vssd1 vssd1 vccd1 vccd1 _14425_/D sky130_fd_sc_hd__clkbuf_1
X_10814_ _10853_/B _10853_/C _10853_/A vssd1 vssd1 vccd1 vccd1 _10846_/C sky130_fd_sc_hd__o21ai_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11794_ _13194_/A vssd1 vssd1 vccd1 vccd1 _11855_/A sky130_fd_sc_hd__clkbuf_4
X_13533_ _13539_/A _13533_/B vssd1 vssd1 vccd1 vccd1 _13534_/A sky130_fd_sc_hd__and2_1
XFILLER_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ _11184_/S _10730_/A _10744_/X _10730_/B vssd1 vssd1 vccd1 vccd1 _10746_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13464_ input89/X _14386_/Q _13467_/S vssd1 vssd1 vccd1 vccd1 _13465_/B sky130_fd_sc_hd__mux2_1
XFILLER_40_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10676_ _10676_/A vssd1 vssd1 vccd1 vccd1 _11186_/S sky130_fd_sc_hd__buf_2
XFILLER_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12415_ _12415_/A vssd1 vssd1 vccd1 vccd1 _12415_/Y sky130_fd_sc_hd__inv_2
X_13395_ _13467_/S vssd1 vssd1 vccd1 vccd1 _13408_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12346_ _12347_/A vssd1 vssd1 vccd1 vccd1 _12346_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11780__A2 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10543__S _10585_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ _12279_/A vssd1 vssd1 vccd1 vccd1 _12277_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12324__A _12348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14016_ _14020_/CLK _14016_/D vssd1 vssd1 vccd1 vccd1 _14016_/Q sky130_fd_sc_hd__dfxtp_1
X_11228_ _11228_/A _11228_/B vssd1 vssd1 vccd1 vccd1 _11229_/B sky130_fd_sc_hd__nor2_2
XFILLER_96_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10966__S1 _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ _13911_/Q _13912_/Q _13913_/Q _13914_/Q _11171_/S _10721_/C vssd1 vssd1 vccd1
+ vccd1 _11159_/X sky130_fd_sc_hd__mux4_1
XFILLER_1_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13285__A2 _13315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08249__A _08249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _09378_/A _08579_/A _13874_/Q _09457_/D vssd1 vssd1 vccd1 vccd1 _08370_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_90_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12796__A1 _14114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07321_ _07376_/A vssd1 vssd1 vccd1 vccd1 _07321_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09661__A1 _10613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07252_ _14078_/Q _13878_/Q _07252_/S vssd1 vssd1 vccd1 vccd1 _07252_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07183_ _14282_/Q _07182_/X _07183_/S vssd1 vssd1 vccd1 vccd1 _07184_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09964__A2 _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12234__A _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07047__B _14271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _09824_/A _09824_/B vssd1 vssd1 vccd1 vccd1 _10037_/A sky130_fd_sc_hd__xnor2_4
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09543__A _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06967_ _06967_/A vssd1 vssd1 vccd1 vccd1 _14314_/D sky130_fd_sc_hd__clkbuf_1
X_09755_ _09755_/A _09755_/B vssd1 vssd1 vccd1 vccd1 _09755_/X sky130_fd_sc_hd__and2_2
XANTENNA__13276__A2 _13236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08706_ _08706_/A _08706_/B vssd1 vssd1 vccd1 vccd1 _08707_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09686_ _09678_/X _09677_/Y _09676_/Y _09676_/B vssd1 vssd1 vccd1 vccd1 _09687_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06898_ _06879_/X _14323_/Q _06898_/S vssd1 vssd1 vccd1 vccd1 _06899_/A sky130_fd_sc_hd__mux2_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _08637_/A _08637_/B vssd1 vssd1 vccd1 vccd1 _08639_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _08568_/A _08562_/B vssd1 vssd1 vccd1 vccd1 _08619_/A sky130_fd_sc_hd__or2b_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12787__A1 _14153_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07519_ _07519_/A vssd1 vssd1 vccd1 vccd1 _07519_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08499_ _08560_/B _08499_/B vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__nor2_1
XFILLER_11_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07112__C1 _14359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10530_ _10530_/A _10530_/B vssd1 vssd1 vccd1 vccd1 _10530_/Y sky130_fd_sc_hd__nand2_4
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _10461_/A _10546_/C vssd1 vssd1 vccd1 vccd1 _10461_/X sky130_fd_sc_hd__or2_1
XFILLER_13_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12200_ _07323_/X _12201_/A _12205_/B _13838_/Q vssd1 vssd1 vccd1 vccd1 _12200_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13180_ _13183_/A vssd1 vssd1 vccd1 vccd1 _13180_/Y sky130_fd_sc_hd__inv_2
X_10392_ _10392_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10413_/A sky130_fd_sc_hd__nor2_2
XFILLER_108_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12131_ _12203_/A vssd1 vssd1 vccd1 vccd1 _12131_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12144__A _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12062_ _12065_/A _12062_/B vssd1 vssd1 vccd1 vccd1 _12063_/A sky130_fd_sc_hd__and2_1
XANTENNA__07238__A _07258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11013_ _13919_/Q vssd1 vssd1 vccd1 vccd1 _11014_/B sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_33_io_wbs_clk clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13963_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_81_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13267__A2 _13236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12964_ _12966_/A vssd1 vssd1 vccd1 vccd1 _12964_/Y sky130_fd_sc_hd__inv_2
XFILLER_73_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11915_ _13820_/Q _11882_/A _11914_/Y _11703_/B vssd1 vssd1 vccd1 vccd1 _11916_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output111_A _11745_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _14146_/Q _12885_/X _12894_/X _12892_/X vssd1 vssd1 vccd1 vccd1 _14146_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12227__B1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _14341_/Q _11833_/X _11848_/A _13800_/Q _11845_/X vssd1 vssd1 vccd1 vccd1
+ _11846_/X sky130_fd_sc_hd__a221o_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _13206_/A vssd1 vssd1 vccd1 vccd1 _13194_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10765__C _11186_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ _10758_/A _10950_/S _07798_/A vssd1 vssd1 vccd1 vccd1 _10729_/A sky130_fd_sc_hd__nor3b_1
X_13516_ _13516_/A vssd1 vssd1 vccd1 vccd1 _14401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11450__A1 _11087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10659_ _11322_/A vssd1 vssd1 vccd1 vccd1 _11108_/A sky130_fd_sc_hd__buf_4
X_13447_ _13447_/A vssd1 vssd1 vccd1 vccd1 _13460_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_16_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_72_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14239_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09628__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ _13467_/S vssd1 vssd1 vccd1 vccd1 _13391_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12329_ _12329_/A vssd1 vssd1 vccd1 vccd1 _12329_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07709__A1 hold3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07870_ _07869_/Y _13983_/Q _07874_/S vssd1 vssd1 vccd1 vccd1 _07871_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11910__C1 hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09540_ _09540_/A _09540_/B _09540_/C vssd1 vssd1 vccd1 vccd1 _09540_/Y sky130_fd_sc_hd__nand3_1
XFILLER_3_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10302__A _10302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08134__B2 _08249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09471_ _09471_/A _09471_/B _09471_/C vssd1 vssd1 vccd1 vccd1 _09471_/Y sky130_fd_sc_hd__nand3_1
XFILLER_110_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08685__A2 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08422_ _09457_/B vssd1 vssd1 vccd1 vccd1 _08449_/B sky130_fd_sc_hd__buf_2
XFILLER_63_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09810__B _13866_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _08353_/A _08353_/B _08353_/C vssd1 vssd1 vccd1 vccd1 _08366_/B sky130_fd_sc_hd__nand3_2
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07304_ _07274_/A _07312_/A _07491_/A _07307_/A vssd1 vssd1 vccd1 vccd1 _07305_/S
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11441__A1 _11079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ _08632_/A _09001_/B _08284_/C _09834_/A vssd1 vssd1 vccd1 vccd1 _08287_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__13718__A0 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07235_ _14083_/Q _13883_/Q _07235_/S vssd1 vssd1 vccd1 vccd1 _07235_/X sky130_fd_sc_hd__mux2_2
XFILLER_30_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09398__B1 _09396_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ _07166_/A vssd1 vssd1 vccd1 vccd1 _14287_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07097_ _14265_/Q _07085_/X _07096_/X _14361_/Q vssd1 vssd1 vccd1 vccd1 _07097_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07324__B_N _07323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09273__A _09273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09807_ _09807_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _09807_/X sky130_fd_sc_hd__and2_2
XFILLER_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07999_ _07997_/X _07999_/B vssd1 vssd1 vccd1 vccd1 _08003_/A sky130_fd_sc_hd__and2b_1
XFILLER_87_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09738_ _09704_/X _09706_/Y _09739_/C _09737_/X vssd1 vssd1 vccd1 vccd1 _10540_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_56_io_wbs_clk_A clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_39_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09669_ _08298_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__and2b_1
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _13758_/Q _13757_/Q _11906_/B vssd1 vssd1 vccd1 vccd1 _11911_/B sky130_fd_sc_hd__or3_1
XANTENNA__13523__A _13539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12680_ _13072_/A vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11631_/A _11631_/B vssd1 vssd1 vccd1 vccd1 _11631_/Y sky130_fd_sc_hd__xnor2_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12139__A input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14350_ _14354_/CLK _14350_/D vssd1 vssd1 vccd1 vccd1 _14350_/Q sky130_fd_sc_hd__dfxtp_1
X_11562_ _14046_/Q _13958_/Q vssd1 vssd1 vccd1 vccd1 _11630_/B sky130_fd_sc_hd__nand2_1
X_13301_ _13343_/A vssd1 vssd1 vccd1 vccd1 _13301_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10513_ _10528_/A vssd1 vssd1 vccd1 vccd1 _10644_/A sky130_fd_sc_hd__buf_2
X_14281_ _14281_/CLK _14281_/D _13143_/Y vssd1 vssd1 vccd1 vccd1 _14281_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11978__A _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11493_ _11493_/A _11493_/B vssd1 vssd1 vccd1 vccd1 _11493_/X sky130_fd_sc_hd__or2_1
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13232_ _14407_/Q _13230_/X _13231_/X vssd1 vssd1 vccd1 vccd1 _13232_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input72_A io_wbs_datwr[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10446_/A sky130_fd_sc_hd__and2_1
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13163_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13163_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08061__B1 _09233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10375_ _10323_/B _10588_/A _10374_/Y vssd1 vssd1 vccd1 vccd1 _10375_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12114_ _13731_/A vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13094_ _13106_/A _13094_/B vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__and2_1
XFILLER_46_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10106__B _10106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output159_A _14314_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ _12045_/A vssd1 vssd1 vccd1 vccd1 _13795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13996_ _14442_/CLK _13996_/D vssd1 vssd1 vccd1 vccd1 _13996_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12947_ _12950_/A vssd1 vssd1 vccd1 vccd1 _12947_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12922_/A _12883_/B vssd1 vssd1 vccd1 vccd1 _12878_/X sky130_fd_sc_hd__or2_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11829_ _13999_/Q _11797_/X _11823_/X _13793_/Q _11828_/X vssd1 vssd1 vccd1 vccd1
+ _11829_/X sky130_fd_sc_hd__a221o_2
XFILLER_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12049__A _12536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11423__A1 _11058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07150__B _14259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07020_ _14419_/Q _07020_/B _14451_/Q vssd1 vssd1 vccd1 vccd1 _07020_/X sky130_fd_sc_hd__and3b_1
XANTENNA__12923__A1 _14156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08971_ _08971_/A _08971_/B vssd1 vssd1 vccd1 vccd1 _08973_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07922_ _13970_/Q _07922_/B vssd1 vssd1 vccd1 vccd1 _13970_/D sky130_fd_sc_hd__xnor2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07606__A _14256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07853_ _14035_/Q _13981_/Q vssd1 vssd1 vccd1 vccd1 _07876_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07497__B_N _07452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07784_ _11322_/A vssd1 vssd1 vccd1 vccd1 _07784_/X sky130_fd_sc_hd__buf_2
XFILLER_83_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09523_ _09468_/A _09468_/B _09522_/Y vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09821__A _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09855__A1 _09482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13343__A _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ _09423_/A _09423_/Y _09452_/X _09453_/Y vssd1 vssd1 vccd1 vccd1 _09454_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_101_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08437__A _13865_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08405_ _08402_/X _08403_/X _08406_/A _08404_/Y vssd1 vssd1 vccd1 vccd1 _09735_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09385_ _09385_/A _09385_/B _09385_/C vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__and3_1
XFILLER_101_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12611__A0 _12610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _08336_/A _08336_/B _08336_/C vssd1 vssd1 vccd1 vccd1 _08337_/A sky130_fd_sc_hd__or3_1
X_08267_ _08403_/A vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__buf_2
X_07218_ _14088_/Q hold35/A _07218_/S vssd1 vssd1 vccd1 vccd1 _07218_/X sky130_fd_sc_hd__mux2_2
XFILLER_119_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08198_ _08198_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08199_/B sky130_fd_sc_hd__or2_1
XANTENNA__12914__A1 _14153_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ _11663_/B vssd1 vssd1 vccd1 vccd1 _14259_/D sky130_fd_sc_hd__clkinv_4
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10160_ _10172_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10091_ _10091_/A _10091_/B vssd1 vssd1 vccd1 vccd1 _10333_/B sky130_fd_sc_hd__xnor2_4
XFILLER_86_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11038__A _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13850_ _14198_/CLK _13850_/D _12244_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12801_ _12801_/A vssd1 vssd1 vccd1 vccd1 _12801_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09731__A _09777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10993_ _10993_/A _10993_/B vssd1 vssd1 vccd1 vccd1 _11079_/B sky130_fd_sc_hd__xnor2_1
X_13781_ _14348_/CLK _13781_/D _11980_/Y vssd1 vssd1 vccd1 vccd1 _13781_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12850__A0 _12650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12732_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08347__A _13868_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12663_/A vssd1 vssd1 vccd1 vccd1 _14048_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14402_ _14451_/CLK _14402_/D vssd1 vssd1 vccd1 vccd1 _14402_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07609__A0 _14079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11614_ _11614_/A _11614_/B vssd1 vssd1 vccd1 vccd1 _11614_/Y sky130_fd_sc_hd__xnor2_4
X_12594_ _12594_/A _12594_/B vssd1 vssd1 vccd1 vccd1 _12595_/A sky130_fd_sc_hd__and2_1
XFILLER_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14333_ _14396_/CLK _14333_/D vssd1 vssd1 vccd1 vccd1 _14333_/Q sky130_fd_sc_hd__dfxtp_1
X_11545_ _14047_/Q _13959_/Q vssd1 vssd1 vccd1 vccd1 _11545_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11476_ _11079_/A _11460_/X _11475_/X _11300_/A _11461_/X vssd1 vssd1 vccd1 vccd1
+ _11476_/X sky130_fd_sc_hd__o221a_1
X_14264_ _14281_/CLK _14264_/D _13121_/Y vssd1 vssd1 vccd1 vccd1 _14264_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08513__C _09200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12905__A1 _14149_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ _13215_/A vssd1 vssd1 vccd1 vccd1 _13215_/X sky130_fd_sc_hd__buf_2
X_10427_ _09766_/A _10430_/S _10426_/X vssd1 vssd1 vccd1 vccd1 _10428_/B sky130_fd_sc_hd__a21o_1
X_14195_ _14224_/CLK _14195_/D _12985_/Y vssd1 vssd1 vccd1 vccd1 _14195_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09782__B1 _09781_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09906__A _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13146_ _13146_/A vssd1 vssd1 vccd1 vccd1 _13146_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10358_ _10358_/A _10381_/A vssd1 vssd1 vccd1 vccd1 _10360_/C sky130_fd_sc_hd__xnor2_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _13089_/A _13077_/B vssd1 vssd1 vccd1 vccd1 _13078_/A sky130_fd_sc_hd__and2_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _10290_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _10289_/Y sky130_fd_sc_hd__nor2_1
X_12028_ _12216_/A vssd1 vssd1 vccd1 vccd1 _12044_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14101__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09641__A _09641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13979_ _14107_/CLK _13979_/D _12406_/Y vssd1 vssd1 vccd1 vccd1 _13979_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ _09216_/A _09168_/C _09168_/B vssd1 vssd1 vccd1 vccd1 _09171_/C sky130_fd_sc_hd__o21ai_1
XFILLER_30_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08121_ _08389_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _08122_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07076__A1 _14300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09088__A _09088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ _08325_/A _08325_/B _08325_/C vssd1 vssd1 vccd1 vccd1 _08052_/Y sky130_fd_sc_hd__nand3_1
X_07003_ _14421_/Q _07020_/B _14453_/Q vssd1 vssd1 vccd1 vccd1 _07003_/X sky130_fd_sc_hd__and3b_1
XANTENNA__10907__B1 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08954_ _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _08954_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07336__A _07363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07905_ _07840_/A _07839_/B _07909_/A _07839_/D vssd1 vssd1 vccd1 vccd1 _07905_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08885_ _08885_/A _08885_/B vssd1 vssd1 vccd1 vccd1 _08887_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07836_ _14026_/Q _13972_/Q vssd1 vssd1 vccd1 vccd1 _07836_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13085__A0 _13084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__A _14020_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07767_ _13986_/Q vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09506_ _08098_/X _09459_/C _09459_/B vssd1 vssd1 vccd1 vccd1 _09511_/A sky130_fd_sc_hd__o21bai_1
XFILLER_24_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07698_ _07661_/X _07697_/X _07657_/Y _14144_/Q vssd1 vssd1 vccd1 vccd1 _07698_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _09437_/A _09437_/B _09437_/C vssd1 vssd1 vccd1 vccd1 _09440_/A sky130_fd_sc_hd__nand3_1
XANTENNA__11305__B _11305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13388__A1 _14364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09482_/A _09842_/A vssd1 vssd1 vccd1 vccd1 _09371_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08319_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _08322_/C sky130_fd_sc_hd__nand2_1
X_09299_ _09377_/A _09299_/B _09299_/C vssd1 vssd1 vccd1 vccd1 _09302_/A sky130_fd_sc_hd__or3_1
XANTENNA__12417__A _13010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08614__B _08658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11330_/A _11330_/B _11334_/A vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__and3_1
X_14475__187 vssd1 vssd1 vccd1 vccd1 _14475__187/HI io_oeb[7] sky130_fd_sc_hd__conb_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11261_ _11262_/A _11355_/B _11262_/C vssd1 vssd1 vccd1 vccd1 _11264_/B sky130_fd_sc_hd__o21a_1
X_10212_ _10214_/A _10214_/B vssd1 vssd1 vccd1 vccd1 _10213_/C sky130_fd_sc_hd__or2_1
XFILLER_97_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13000_ _13003_/A vssd1 vssd1 vccd1 vccd1 _13000_/Y sky130_fd_sc_hd__inv_2
X_11192_ _10650_/A _11158_/X _11143_/A vssd1 vssd1 vccd1 vccd1 _11233_/A sky130_fd_sc_hd__o21ai_4
XFILLER_106_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10143_ _10143_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10074_ _10098_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10074_/X sky130_fd_sc_hd__and2_1
XANTENNA_input35_A io_wbs_adr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13902_ _13905_/CLK _13902_/D _12310_/Y vssd1 vssd1 vccd1 vccd1 _13902_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13076__A0 _12641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13833_ _14441_/CLK _13833_/D vssd1 vssd1 vccd1 vccd1 _13833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09819__A1 _09233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13764_ _13825_/CLK _13764_/D _11956_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Q sky130_fd_sc_hd__dfrtp_1
X_10976_ _10918_/A _10917_/X _10964_/X _10735_/X _10975_/X vssd1 vssd1 vccd1 vccd1
+ _11017_/A sky130_fd_sc_hd__o221a_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12715_ _12715_/A vssd1 vssd1 vccd1 vccd1 _12715_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13695_ _13695_/A _13695_/B vssd1 vssd1 vccd1 vccd1 _13696_/A sky130_fd_sc_hd__and2_1
X_12646_ _12695_/S vssd1 vssd1 vccd1 vccd1 _12665_/S sky130_fd_sc_hd__buf_2
XFILLER_106_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07058__A1 _14270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12577_ _12577_/A vssd1 vssd1 vccd1 vccd1 _14026_/D sky130_fd_sc_hd__clkbuf_1
X_14316_ _14453_/CLK _14316_/D _13186_/Y vssd1 vssd1 vccd1 vccd1 _14316_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11528_ _08944_/D _11510_/X _11526_/X _11527_/X vssd1 vssd1 vccd1 vccd1 _13861_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14247_ _14250_/CLK _14247_/D vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dfxtp_1
X_11459_ _11467_/A _13945_/Q vssd1 vssd1 vccd1 vccd1 _11513_/A sky130_fd_sc_hd__or2_1
XFILLER_113_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14178_ _14256_/CLK _14178_/D _12964_/Y vssd1 vssd1 vccd1 vccd1 _14178_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07230__A1 _07229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13147_/A vssd1 vssd1 vccd1 vccd1 _13134_/A sky130_fd_sc_hd__buf_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09507__B1 _09821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08670_ _08670_/A _08670_/B vssd1 vssd1 vccd1 vccd1 _08670_/X sky130_fd_sc_hd__and2_1
XFILLER_94_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07621_ _14132_/Q _14067_/Q vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07552_ _14105_/Q input22/X _07560_/S vssd1 vssd1 vccd1 vccd1 _07553_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_7_0_io_wbs_clk_A clkbuf_3_7_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07483_ _07483_/A _07483_/B vssd1 vssd1 vccd1 vccd1 _07483_/X sky130_fd_sc_hd__or2_1
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ _09295_/A _09220_/C _09220_/B vssd1 vssd1 vccd1 vccd1 _09223_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__08137__D _10000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08715__A _09084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _09153_/A _09153_/B _09807_/A _09361_/D vssd1 vssd1 vccd1 vccd1 _09155_/A
+ sky130_fd_sc_hd__and4_1
X_08104_ _08789_/A vssd1 vssd1 vccd1 vccd1 _09234_/A sky130_fd_sc_hd__buf_2
XFILLER_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09084_ _09084_/A _09084_/B _09084_/C _09084_/D vssd1 vssd1 vccd1 vccd1 _09087_/A
+ sky130_fd_sc_hd__nand4_2
X_08035_ _14016_/Q vssd1 vssd1 vccd1 vccd1 _08579_/A sky130_fd_sc_hd__clkbuf_2
Xinput80 io_wbs_datwr[22] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__buf_2
Xinput91 io_wbs_datwr[3] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__buf_4
XFILLER_116_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08549__A1 _08571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08549__B2 _08128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09986_ _09986_/A _09986_/B vssd1 vssd1 vccd1 vccd1 _09986_/X sky130_fd_sc_hd__or2_1
XFILLER_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08937_ _08946_/A _08937_/B _08937_/C _10156_/A vssd1 vssd1 vccd1 vccd1 _08941_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_112_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12502__C1 _12498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08868_ _08896_/A _08925_/C _10057_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08869_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_85_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ _14034_/Q _13980_/Q vssd1 vssd1 vccd1 vccd1 _07819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08799_ _08799_/A _08799_/B _08799_/C vssd1 vssd1 vccd1 vccd1 _08820_/A sky130_fd_sc_hd__nand3_1
XFILLER_44_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10830_ _10669_/X _10828_/Y _10829_/X _10675_/X _13943_/Q vssd1 vssd1 vccd1 vccd1
+ _13943_/D sky130_fd_sc_hd__a32o_1
XFILLER_60_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10761_ _10918_/A _10761_/B _10761_/C vssd1 vssd1 vccd1 vccd1 _10761_/X sky130_fd_sc_hd__or3_1
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12500_ _10547_/A _12486_/X _12476_/A _14055_/Q vssd1 vssd1 vccd1 vccd1 _12500_/X
+ sky130_fd_sc_hd__a22o_1
X_10692_ _13944_/Q vssd1 vssd1 vccd1 vccd1 _11262_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13480_ _13485_/A _13480_/B vssd1 vssd1 vccd1 vccd1 _13481_/A sky130_fd_sc_hd__and2_1
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12431_ _14040_/Q _13200_/B _12425_/B vssd1 vssd1 vccd1 vccd1 _12431_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__12147__A _12147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ _12366_/A vssd1 vssd1 vccd1 vccd1 _12362_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14101_ _14102_/CLK _14101_/D _12751_/Y vssd1 vssd1 vccd1 vccd1 _14101_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11986__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11313_ _11312_/A _11312_/B _11312_/C vssd1 vssd1 vccd1 vccd1 _11313_/Y sky130_fd_sc_hd__a21oi_1
X_12293_ _12317_/A vssd1 vssd1 vccd1 vccd1 _12298_/A sky130_fd_sc_hd__buf_2
XFILLER_5_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11244_ _11244_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11245_/B sky130_fd_sc_hd__nand2_1
X_14032_ _14054_/CLK _14032_/D vssd1 vssd1 vccd1 vccd1 _14032_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_10_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09201__A2 _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11175_ _13915_/Q _13916_/Q _11175_/S vssd1 vssd1 vccd1 vccd1 _11175_/X sky130_fd_sc_hd__mux2_1
X_10126_ _10126_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _10127_/B sky130_fd_sc_hd__xor2_2
XFILLER_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output141_A _11819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10057_ _10057_/A vssd1 vssd1 vccd1 vccd1 _10065_/A sky130_fd_sc_hd__inv_2
XFILLER_36_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08519__B _08815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13816_ _13826_/CLK _13816_/D vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13747_ _14335_/CLK _13747_/D _11931_/X vssd1 vssd1 vccd1 vccd1 _13747_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10959_ _13900_/Q _13901_/Q _13902_/Q _13903_/Q _11175_/S _10676_/A vssd1 vssd1 vccd1
+ vccd1 _10959_/X sky130_fd_sc_hd__mux4_2
XFILLER_17_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13678_ _13678_/A _13678_/B vssd1 vssd1 vccd1 vccd1 _13679_/A sky130_fd_sc_hd__and2_1
XFILLER_19_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12629_ _12629_/A vssd1 vssd1 vccd1 vccd1 _14040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08270__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09840_ _09969_/A _09968_/B vssd1 vssd1 vccd1 vccd1 _10463_/S sky130_fd_sc_hd__nand2_4
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09771_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09772_/B sky130_fd_sc_hd__xor2_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _06980_/X _14312_/Q _06983_/S vssd1 vssd1 vccd1 vccd1 _06984_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08722_ _08722_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _08734_/B sky130_fd_sc_hd__xnor2_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08653_ _08449_/B _09804_/A _09000_/B _08983_/A vssd1 vssd1 vccd1 vccd1 _08654_/C
+ sky130_fd_sc_hd__a22oi_4
XFILLER_96_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07604_ _14081_/Q input28/X _07604_/S vssd1 vssd1 vccd1 vccd1 _07605_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08584_ _08584_/A _08637_/B _08584_/C vssd1 vssd1 vccd1 vccd1 _08586_/A sky130_fd_sc_hd__and3_1
XFILLER_54_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12799__C1 _12216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07535_ _14182_/Q _07526_/X _07533_/X _07534_/Y _07519_/X vssd1 vssd1 vccd1 vccd1
+ _14174_/D sky130_fd_sc_hd__o221a_1
X_07466_ _07483_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _07466_/X sky130_fd_sc_hd__or2_1
XFILLER_50_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09205_ _09205_/A _09205_/B _09205_/C vssd1 vssd1 vccd1 vccd1 _09212_/A sky130_fd_sc_hd__nand3_1
XFILLER_10_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07397_ _07376_/X _07395_/X _07396_/X _07379_/X vssd1 vssd1 vccd1 vccd1 _07397_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09136_ _09130_/A _09130_/B _09130_/C vssd1 vssd1 vccd1 vccd1 _09137_/C sky130_fd_sc_hd__a21o_1
XFILLER_108_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09067_ _09067_/A _09067_/B _09067_/C vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__and3_1
XFILLER_118_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08018_ _09434_/A _08284_/C vssd1 vssd1 vccd1 vccd1 _08131_/A sky130_fd_sc_hd__nand2_2
XFILLER_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08180__A _09336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13947_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__10215__A _10215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09969_ _09969_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _09970_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13526__A _13526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12980_ _13004_/A vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11931_ _12216_/A vssd1 vssd1 vccd1 vccd1 _11931_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _14351_/Q _11864_/B vssd1 vssd1 vccd1 vccd1 _11863_/A sky130_fd_sc_hd__and2_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _13607_/A _13601_/B vssd1 vssd1 vccd1 vccd1 _13602_/A sky130_fd_sc_hd__and2_1
XFILLER_26_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13451__A0 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10813_ _10846_/B _10813_/B vssd1 vssd1 vccd1 vccd1 _10853_/A sky130_fd_sc_hd__and2_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _11848_/A vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13532_ _13084_/X _14405_/Q _13542_/S vssd1 vssd1 vccd1 vccd1 _13533_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10744_ _10744_/A vssd1 vssd1 vccd1 vccd1 _10744_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13463_ _13504_/A vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__clkbuf_4
X_10675_ _11100_/A vssd1 vssd1 vccd1 vccd1 _10675_/X sky130_fd_sc_hd__buf_2
XFILLER_40_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12414_ _12415_/A vssd1 vssd1 vccd1 vccd1 _12414_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_62_io_wbs_clk clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14363_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_12_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13394_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13409_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_63_io_wbs_clk_A clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12345_ _12347_/A vssd1 vssd1 vccd1 vccd1 _12345_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12276_ _12279_/A vssd1 vssd1 vccd1 vccd1 _12276_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14015_ _14020_/CLK _14015_/D vssd1 vssd1 vccd1 vccd1 _14015_/Q sky130_fd_sc_hd__dfxtp_1
X_11227_ _13903_/Q vssd1 vssd1 vccd1 vccd1 _11288_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08933__A1 _08896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11158_ _11149_/B _11146_/X _11158_/S vssd1 vssd1 vccd1 vccd1 _11158_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10109_ _10053_/A _10053_/B _10108_/X vssd1 vssd1 vccd1 vccd1 _10116_/A sky130_fd_sc_hd__a21o_1
XFILLER_49_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11089_ _11308_/A _11089_/B vssd1 vssd1 vccd1 vccd1 _11090_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12493__A1 _09762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12493__B2 _14053_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08249__B _09999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09646__C1 _09404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07320_ _13893_/Q _13836_/Q _07464_/A _07263_/A vssd1 vssd1 vccd1 vccd1 _07376_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_32_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07251_ _07251_/A vssd1 vssd1 vccd1 vccd1 _14263_/D sky130_fd_sc_hd__clkbuf_1
X_07182_ _14098_/Q _07167_/X _07168_/X vssd1 vssd1 vccd1 vccd1 _07182_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07424__A1 _07399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12515__A input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09824__A _09824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _10151_/A _09826_/B vssd1 vssd1 vccd1 vccd1 _09926_/A sky130_fd_sc_hd__nor2_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _08245_/A _08245_/B _08244_/A vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__a21o_1
X_06966_ _06963_/X _14314_/Q _06966_/S vssd1 vssd1 vccd1 vccd1 _06967_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12250__A _12251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08705_ _09132_/A _09132_/B _09206_/B _09873_/A vssd1 vssd1 vccd1 vccd1 _08706_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_100_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13681__A0 _12610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ _09685_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__xnor2_2
X_06897_ _06894_/X _06896_/X _14365_/Q vssd1 vssd1 vccd1 vccd1 _06898_/S sky130_fd_sc_hd__o21a_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14335__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _08636_/A _08998_/B _08636_/C vssd1 vssd1 vccd1 vccd1 _08639_/A sky130_fd_sc_hd__nand3_1
XANTENNA__07063__B _14260_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08567_ _08567_/A _08731_/A vssd1 vssd1 vccd1 vccd1 _08613_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07518_ _07518_/A vssd1 vssd1 vccd1 vccd1 _14179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08498_ _09000_/A _08893_/A _08560_/A _08490_/Y vssd1 vssd1 vccd1 vccd1 _08499_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07449_ _07458_/A _07449_/B vssd1 vssd1 vccd1 vccd1 _07449_/X sky130_fd_sc_hd__or2_1
XFILLER_109_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_io_wbs_clk clkbuf_2_3_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_io_wbs_clk/A
+ sky130_fd_sc_hd__clkbuf_2
X_10460_ _10412_/A _10417_/A _10459_/X vssd1 vssd1 vccd1 vccd1 _10546_/C sky130_fd_sc_hd__a21o_1
XFILLER_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07415__A1 _14208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09119_ _09119_/A _09119_/B vssd1 vssd1 vccd1 vccd1 _09191_/A sky130_fd_sc_hd__nor2_2
X_10391_ _10391_/A _10391_/B _10391_/C vssd1 vssd1 vccd1 vccd1 _10392_/B sky130_fd_sc_hd__and3_1
XANTENNA__12425__A _14007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08622__B _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12130_ input74/X _12130_/B vssd1 vssd1 vccd1 vccd1 _12130_/X sky130_fd_sc_hd__or2_1
XFILLER_11_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12061_ _13799_/Q _12059_/X _12060_/X _13815_/Q vssd1 vssd1 vccd1 vccd1 _12062_/B
+ sky130_fd_sc_hd__a22o_1
X_11012_ _11012_/A _11012_/B vssd1 vssd1 vccd1 vccd1 _11064_/B sky130_fd_sc_hd__xor2_1
XFILLER_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12160__A _12911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12963_ _12966_/A vssd1 vssd1 vccd1 vccd1 _12963_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10486__A0 _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11914_ _13760_/Q _11914_/B vssd1 vssd1 vccd1 vccd1 _11914_/Y sky130_fd_sc_hd__nand2_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12894_ _12938_/A _12896_/B vssd1 vssd1 vccd1 vccd1 _12894_/X sky130_fd_sc_hd__or2_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _14006_/Q _11845_/B vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__and2_1
XFILLER_60_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _12193_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _13206_/A sky130_fd_sc_hd__nor2_4
XANTENNA__07103__B1 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09643__A2 _09404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13515_ _13518_/A _13515_/B vssd1 vssd1 vccd1 vccd1 _13516_/A sky130_fd_sc_hd__and2_1
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10727_ _13939_/Q _10727_/B _10727_/C _10727_/D vssd1 vssd1 vccd1 vccd1 _10840_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13446_ _13504_/A vssd1 vssd1 vccd1 vccd1 _13461_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10658_ _10652_/X _07804_/B _10657_/X vssd1 vssd1 vccd1 vccd1 _13950_/D sky130_fd_sc_hd__o21a_1
XFILLER_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13377_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13392_/A sky130_fd_sc_hd__clkbuf_1
X_10589_ _10589_/A _10589_/B vssd1 vssd1 vccd1 vccd1 _10589_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_103_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12328_ _12329_/A vssd1 vssd1 vccd1 vccd1 _12328_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10961__A1 _10722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12259_ _12259_/A vssd1 vssd1 vccd1 vccd1 _12259_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09644__A _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13166__A _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14358__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12466__A1 _08983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08134__A2 _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09470_ _09454_/Y _09470_/B _09470_/C _09470_/D vssd1 vssd1 vccd1 vccd1 _09470_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08421_ _08750_/B vssd1 vssd1 vccd1 vccd1 _09457_/B sky130_fd_sc_hd__buf_2
XFILLER_63_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08352_ _09555_/B _09555_/C _09555_/A vssd1 vssd1 vccd1 vccd1 _08353_/C sky130_fd_sc_hd__a21bo_1
XFILLER_20_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07303_ _07471_/A vssd1 vssd1 vccd1 vccd1 _07491_/A sky130_fd_sc_hd__clkbuf_2
X_08283_ _09543_/B vssd1 vssd1 vccd1 vccd1 _09001_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07234_ _07234_/A vssd1 vssd1 vccd1 vccd1 _14268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07165_ _14287_/Q _07164_/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07166_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07096_ _14409_/Q _07095_/Y _07087_/X vssd1 vssd1 vccd1 vccd1 _07096_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06908__B1 _06877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09806_ _09806_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _09806_/X sky130_fd_sc_hd__or2_2
XANTENNA__09273__B _09273_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07998_ _09084_/B _08976_/A _09058_/B _09084_/A vssd1 vssd1 vccd1 vccd1 _07999_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09737_ _09739_/B _09732_/X _09731_/Y _09697_/A vssd1 vssd1 vccd1 vccd1 _09737_/X
+ sky130_fd_sc_hd__a211o_1
X_06949_ _07027_/A vssd1 vssd1 vccd1 vccd1 _06981_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09668_ _10576_/A _09655_/B _09664_/X _09666_/X _09667_/Y vssd1 vssd1 vccd1 vccd1
+ _10557_/C sky130_fd_sc_hd__o311a_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07802__A _11175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _08619_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__and2_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _08366_/B _08363_/B _08363_/C vssd1 vssd1 vccd1 vccd1 _09601_/B sky130_fd_sc_hd__a21o_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07521__B _07521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11546_/Y _11630_/B vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__and2b_1
XFILLER_11_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09625__A2 _09396_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ _11634_/B _11634_/C _11634_/A vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__o21ba_1
XFILLER_7_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13300_ _14421_/Q _13284_/X _13298_/X _13299_/X vssd1 vssd1 vccd1 vccd1 _13300_/X
+ sky130_fd_sc_hd__a211o_1
X_10512_ _08412_/Y _10524_/B _09751_/Y vssd1 vssd1 vccd1 vccd1 _10512_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10640__B1 _09788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14280_ _14281_/CLK _14280_/D _13142_/Y vssd1 vssd1 vccd1 vccd1 _14280_/Q sky130_fd_sc_hd__dfrtp_4
X_11492_ _08767_/B _11486_/X _11488_/Y _11491_/X vssd1 vssd1 vccd1 vccd1 _13869_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13231_ _14439_/Q _13336_/A _13218_/X _14391_/Q vssd1 vssd1 vccd1 vccd1 _13231_/X
+ sky130_fd_sc_hd__a22o_1
X_10443_ _10428_/B _10367_/A _10443_/S vssd1 vssd1 vccd1 vccd1 _10445_/B sky130_fd_sc_hd__mux2_1
XFILLER_40_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input65_A io_wbs_cyc vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13162_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08061__A1 _08251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _10374_/A _10374_/B _10374_/C vssd1 vssd1 vccd1 vccd1 _10374_/Y sky130_fd_sc_hd__nand3_1
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12113_ _13609_/A vssd1 vssd1 vccd1 vccd1 _13731_/A sky130_fd_sc_hd__buf_4
XFILLER_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13093_ _12579_/X hold32/A _13096_/S vssd1 vssd1 vccd1 vccd1 _13094_/B sky130_fd_sc_hd__mux2_1
X_12044_ _12044_/A _12044_/B vssd1 vssd1 vccd1 vccd1 _12045_/A sky130_fd_sc_hd__and2_1
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11218__B _11297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13995_ _14441_/CLK _13995_/D vssd1 vssd1 vccd1 vccd1 _13995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13714__A _13731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12946_ _12950_/A vssd1 vssd1 vccd1 vccd1 _12946_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _14139_/Q _12872_/X _12876_/X _12866_/X vssd1 vssd1 vccd1 vccd1 _14139_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _14334_/Q _11855_/A _12254_/B _14118_/Q vssd1 vssd1 vccd1 vccd1 _11828_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11759_ input62/X input46/X _11759_/C _11759_/D vssd1 vssd1 vccd1 vccd1 _11774_/B
+ sky130_fd_sc_hd__or4_4
X_13429_ _13504_/A vssd1 vssd1 vccd1 vccd1 _13444_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08970_ _08970_/A vssd1 vssd1 vccd1 vccd1 _08971_/A sky130_fd_sc_hd__inv_2
XFILLER_103_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14180__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07921_ _14024_/Q _13951_/D _07921_/C vssd1 vssd1 vccd1 vccd1 _07922_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13748__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11895__C1 _11874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09552__B2 _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ _07819_/Y _07882_/A _07881_/B vssd1 vssd1 vccd1 vccd1 _07877_/A sky130_fd_sc_hd__o21ai_1
XFILLER_84_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07563__A0 _14100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput1 dout1[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
X_07783_ _10895_/B vssd1 vssd1 vccd1 vccd1 _11322_/A sky130_fd_sc_hd__clkbuf_4
X_09522_ _09522_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09522_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09821__B _09821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09453_ _09471_/A _09471_/C _09471_/B vssd1 vssd1 vccd1 vccd1 _09453_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08404_ _08337_/A _08400_/Y _09729_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _08404_/Y
+ sky130_fd_sc_hd__a211oi_1
X_09384_ _09441_/A _09382_/B _09382_/C vssd1 vssd1 vccd1 vccd1 _09385_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__07618__A1 _14256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08335_ _08343_/B _08335_/B vssd1 vssd1 vccd1 vccd1 _08336_/C sky130_fd_sc_hd__or2_1
XFILLER_71_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12611__A1 _14036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08266_ _08266_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08273_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07217_ _07217_/A vssd1 vssd1 vccd1 vccd1 _14273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08197_ _08198_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08243_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07148_ _13774_/Q _13772_/Q vssd1 vssd1 vccd1 vccd1 _11663_/B sky130_fd_sc_hd__or2b_4
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09240__B1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07079_ _14411_/Q _07078_/Y _07048_/X vssd1 vssd1 vccd1 vccd1 _07079_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12703__A _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10090_ _10090_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _10091_/B sky130_fd_sc_hd__xor2_2
XFILLER_102_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11319__A _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07554__A0 _14104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12800_ _12800_/A vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13780_ _14427_/CLK _13780_/D _11979_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Q sky130_fd_sc_hd__dfrtp_1
X_10992_ _13924_/Q vssd1 vssd1 vccd1 vccd1 _11079_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12731_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11054__A _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12678_/A _12662_/B vssd1 vssd1 vccd1 vccd1 _12663_/A sky130_fd_sc_hd__and2_1
XFILLER_43_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09059__B1 _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14451_/CLK _14401_/D vssd1 vssd1 vccd1 vccd1 _14401_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11543_/Y _11613_/B vssd1 vssd1 vccd1 vccd1 _11614_/B sky130_fd_sc_hd__and2b_1
XFILLER_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12593_ _12922_/A _14031_/Q _12600_/S vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__mux2_1
X_14332_ _14396_/CLK _14332_/D vssd1 vssd1 vccd1 vccd1 _14332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11544_ _14048_/Q _13960_/Q vssd1 vssd1 vccd1 vccd1 _11544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _14365_/CLK _14263_/D _13120_/Y vssd1 vssd1 vccd1 vccd1 _14263_/Q sky130_fd_sc_hd__dfrtp_2
X_11475_ _11499_/A vssd1 vssd1 vccd1 vccd1 _11475_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11169__A1 _10912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13214_ _13328_/A vssd1 vssd1 vccd1 vccd1 _13215_/A sky130_fd_sc_hd__clkbuf_2
X_10426_ _10399_/B _10426_/B vssd1 vssd1 vccd1 vccd1 _10426_/X sky130_fd_sc_hd__and2b_1
X_14194_ _14224_/CLK _14194_/D _12984_/Y vssd1 vssd1 vccd1 vccd1 _14194_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_output171_A _14296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _13146_/A vssd1 vssd1 vccd1 vccd1 _13145_/Y sky130_fd_sc_hd__inv_2
X_10357_ _10331_/A _10395_/A _09926_/A vssd1 vssd1 vccd1 vccd1 _10381_/A sky130_fd_sc_hd__o21ba_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13076_ _12641_/X hold21/A _13076_/S vssd1 vssd1 vccd1 vccd1 _13077_/B sky130_fd_sc_hd__mux2_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _10288_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10315_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09534__A1 _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12027_ _12027_/A vssd1 vssd1 vccd1 vccd1 _13790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09922__A _10091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13618__A0 input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13978_ _14107_/CLK _13978_/D _12405_/Y vssd1 vssd1 vccd1 vccd1 _13978_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12929_ _12942_/B vssd1 vssd1 vccd1 vccd1 _12940_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08120_ _08120_/A _08120_/B vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__nor2_1
X_08051_ _08119_/C _08051_/B vssd1 vssd1 vccd1 vccd1 _08325_/C sky130_fd_sc_hd__and2_1
XANTENNA__09088__B _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07002_ _14277_/Q _06968_/X _07001_/X _14373_/Q vssd1 vssd1 vccd1 vccd1 _07002_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12523__A _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07617__A hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _08953_/A _08953_/B vssd1 vssd1 vccd1 vccd1 _08954_/B sky130_fd_sc_hd__and2_1
X_07904_ _07904_/A vssd1 vssd1 vccd1 vccd1 _13951_/D sky130_fd_sc_hd__clkbuf_2
X_08884_ _08883_/A _08883_/C _08883_/B vssd1 vssd1 vccd1 vccd1 _08885_/B sky130_fd_sc_hd__o21ai_1
XFILLER_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07835_ _07918_/A _07918_/B _07834_/A vssd1 vssd1 vccd1 vccd1 _07915_/A sky130_fd_sc_hd__o21a_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09551__B _14019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ _07766_/A vssd1 vssd1 vccd1 vccd1 _14060_/D sky130_fd_sc_hd__clkbuf_1
X_09505_ _09450_/A _09448_/X _09449_/A vssd1 vssd1 vccd1 vccd1 _09515_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__11096__B1 _11092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07697_ _14143_/Q _07727_/A _07732_/A _14142_/Q _07696_/X vssd1 vssd1 vccd1 vccd1
+ _07697_/X sky130_fd_sc_hd__a221o_1
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07071__B _14268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09430_/A _09430_/B _09430_/C vssd1 vssd1 vccd1 vccd1 _09437_/C sky130_fd_sc_hd__a21o_1
XFILLER_53_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09367_/A _09367_/B _09367_/C vssd1 vssd1 vccd1 vccd1 _09373_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09279__A _09362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ _08318_/A _08318_/B vssd1 vssd1 vccd1 vccd1 _08364_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08183__A _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09298_ _09217_/B _09817_/B _09479_/D _09165_/A vssd1 vssd1 vccd1 vccd1 _09299_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08249_ _08249_/A _09999_/B vssd1 vssd1 vccd1 vccd1 _08253_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11260_ _13895_/Q vssd1 vssd1 vccd1 vccd1 _11264_/A sky130_fd_sc_hd__inv_2
XANTENNA__12899__A1 _14148_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10211_ _10211_/A _10211_/B vssd1 vssd1 vccd1 vccd1 _10214_/B sky130_fd_sc_hd__xnor2_1
XFILLER_107_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_68_io_wbs_clk_A clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09764__A1 _09188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ _11142_/A _11141_/X _11190_/X vssd1 vssd1 vccd1 vccd1 _11237_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__08630__B _10215_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ _10166_/A _10166_/B _10141_/X vssd1 vssd1 vccd1 vccd1 _10144_/A sky130_fd_sc_hd__a21bo_1
XFILLER_43_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10073_ _10330_/B _10073_/B vssd1 vssd1 vccd1 vccd1 _10099_/B sky130_fd_sc_hd__xnor2_2
XFILLER_48_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12520__A0 _12909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13901_ _13905_/CLK _13901_/D _12309_/Y vssd1 vssd1 vccd1 vccd1 _13901_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input28_A dout1[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ _14164_/CLK _13832_/D vssd1 vssd1 vccd1 vccd1 _13832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08358__A _14019_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13763_ _13825_/CLK _13763_/D _11955_/Y vssd1 vssd1 vccd1 vccd1 _13763_/Q sky130_fd_sc_hd__dfrtp_1
X_10975_ _10975_/A _10975_/B vssd1 vssd1 vccd1 vccd1 _10975_/X sky130_fd_sc_hd__or2_1
XFILLER_44_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _12715_/A vssd1 vssd1 vccd1 vccd1 _12714_/Y sky130_fd_sc_hd__inv_2
X_13694_ input73/X _14452_/Q _13704_/S vssd1 vssd1 vccd1 vccd1 _13695_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12645_ input93/X vssd1 vssd1 vccd1 vccd1 _12645_/X sky130_fd_sc_hd__buf_4
XFILLER_62_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12587__A0 _12917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12576_ _12576_/A _12576_/B vssd1 vssd1 vccd1 vccd1 _12577_/A sky130_fd_sc_hd__and2_1
XFILLER_8_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14315_ _14457_/CLK _14315_/D _13185_/Y vssd1 vssd1 vccd1 vccd1 _14315_/Q sky130_fd_sc_hd__dfrtp_4
X_11527_ _11038_/A _11513_/X _11499_/A _11269_/A _11514_/X vssd1 vssd1 vccd1 vccd1
+ _11527_/X sky130_fd_sc_hd__o221a_1
XFILLER_102_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14246_ _14250_/CLK _14246_/D vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_2
XFILLER_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11458_ _11533_/S _11457_/Y _11467_/A vssd1 vssd1 vccd1 vccd1 _11458_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10409_ _10493_/A _10413_/B _10413_/A vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__mux2_1
X_14177_ _14179_/CLK _14177_/D _12963_/Y vssd1 vssd1 vccd1 vccd1 _14177_/Q sky130_fd_sc_hd__dfrtp_1
X_11389_ _13884_/Q _11379_/X _11383_/X _11388_/X vssd1 vssd1 vccd1 vccd1 _13884_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13128_/A vssd1 vssd1 vccd1 vccd1 _13128_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07437__A _07464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09507__A1 _08791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09507__B2 _08791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ _13059_/A _13059_/B vssd1 vssd1 vccd1 vccd1 _13079_/B sky130_fd_sc_hd__nand2_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11314__A1 _07784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09652__A _09652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ _14069_/Q vssd1 vssd1 vccd1 vccd1 _07662_/A sky130_fd_sc_hd__inv_2
XFILLER_4_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_70_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_47_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07551_ _07595_/A vssd1 vssd1 vccd1 vccd1 _07560_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12814__B2 _14145_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07482_ _14193_/Q _14195_/Q _07482_/S vssd1 vssd1 vccd1 vccd1 _07483_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09221_ _09156_/A _09155_/B _09155_/A vssd1 vssd1 vccd1 vccd1 _09223_/B sky130_fd_sc_hd__o21bai_1
XFILLER_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13936__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11750__B1_N _07548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _09152_/A _09152_/B vssd1 vssd1 vccd1 vccd1 _09156_/A sky130_fd_sc_hd__nand2_1
X_08103_ _09508_/A _09233_/B _09508_/C vssd1 vssd1 vccd1 vccd1 _09535_/B sky130_fd_sc_hd__o21ai_1
X_09083_ _09083_/A _09083_/B vssd1 vssd1 vccd1 vccd1 _09144_/A sky130_fd_sc_hd__nor2_1
X_08034_ _09378_/A vssd1 vssd1 vccd1 vccd1 _08580_/A sky130_fd_sc_hd__clkbuf_4
Xinput70 io_wbs_datwr[13] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__clkbuf_1
Xinput81 io_wbs_datwr[23] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_2
XFILLER_66_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput92 io_wbs_datwr[4] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__buf_4
XANTENNA__08549__A2 _09943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14031_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__12253__A _12259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09985_ _09986_/A _09986_/B vssd1 vssd1 vccd1 vccd1 _09985_/X sky130_fd_sc_hd__and2_1
XFILLER_66_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08936_ _08936_/A vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__buf_4
XANTENNA__07509__A0 hold20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06980__A1 _14280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08867_ _08867_/A vssd1 vssd1 vccd1 vccd1 _08896_/A sky130_fd_sc_hd__buf_4
XANTENNA__13084__A input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07818_ _14035_/Q _13981_/Q vssd1 vssd1 vccd1 vccd1 _07876_/A sky130_fd_sc_hd__or2_1
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08798_ _08798_/A _08798_/B vssd1 vssd1 vccd1 vccd1 _08820_/C sky130_fd_sc_hd__xnor2_1
XFILLER_57_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08178__A _08944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07749_ _07673_/B _07723_/X _07724_/X vssd1 vssd1 vccd1 vccd1 _07749_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10760_ _10765_/A vssd1 vssd1 vccd1 vccd1 _10918_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09419_ _09416_/Y _09417_/X _09263_/X _09415_/Y vssd1 vssd1 vccd1 vccd1 _09420_/B
+ sky130_fd_sc_hd__o211a_1
X_10691_ _10691_/A vssd1 vssd1 vccd1 vccd1 _13945_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12569__A0 _12218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12430_ _12440_/B vssd1 vssd1 vccd1 vccd1 _13200_/B sky130_fd_sc_hd__buf_4
XFILLER_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_io_wbs_clk clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13826_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12361_ _12379_/A vssd1 vssd1 vccd1 vccd1 _12366_/A sky130_fd_sc_hd__buf_4
X_14100_ _14102_/CLK _14100_/D _12750_/Y vssd1 vssd1 vccd1 vccd1 _14100_/Q sky130_fd_sc_hd__dfrtp_2
X_11312_ _11312_/A _11312_/B _11312_/C vssd1 vssd1 vccd1 vccd1 _11312_/X sky130_fd_sc_hd__and3_1
XFILLER_14_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12292_ _12385_/A vssd1 vssd1 vccd1 vccd1 _12317_/A sky130_fd_sc_hd__buf_2
XFILLER_10_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14031_ _14031_/CLK _14031_/D vssd1 vssd1 vccd1 vccd1 _14031_/Q sky130_fd_sc_hd__dfxtp_4
X_11243_ _13899_/Q vssd1 vssd1 vccd1 vccd1 _11276_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12163__A input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11174_ _11038_/A _11032_/A _11175_/S vssd1 vssd1 vccd1 vccd1 _11174_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14241__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10125_ _10122_/Y _10123_/Y _10124_/Y vssd1 vssd1 vccd1 vccd1 _10283_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__13297__A1 _14340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09472__A _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ _10123_/A _10056_/B vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__xor2_1
XFILLER_75_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08088__A _14011_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11226__B _11291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13815_ _13826_/CLK _13815_/D vssd1 vssd1 vccd1 vccd1 _13815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ _13746_/A vssd1 vssd1 vccd1 vccd1 _14467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10958_ _10957_/X _10923_/X _11158_/S vssd1 vssd1 vccd1 vccd1 _10958_/X sky130_fd_sc_hd__mux2_2
XFILLER_91_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13677_ _12673_/X _14447_/Q _13687_/S vssd1 vssd1 vccd1 vccd1 _13678_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10889_ _10889_/A _10889_/B _10889_/C vssd1 vssd1 vccd1 vccd1 _10889_/X sky130_fd_sc_hd__or3_1
X_12628_ _12635_/A _12628_/B vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__and2_1
XFILLER_8_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12559_ _12576_/A _12559_/B vssd1 vssd1 vccd1 vccd1 _12560_/A sky130_fd_sc_hd__and2_1
XFILLER_89_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14229_ _14256_/CLK _14229_/D _13027_/Y vssd1 vssd1 vccd1 vccd1 _14229_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07167__A _07185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10305__B _10305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09770_/A _09770_/B vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__xnor2_1
XFILLER_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13288__A1 _14338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06982_ _06973_/X _06981_/X _14376_/Q vssd1 vssd1 vccd1 vccd1 _06983_/S sky130_fd_sc_hd__o21a_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08530_/A _08529_/A _08529_/B vssd1 vssd1 vccd1 vccd1 _08722_/B sky130_fd_sc_hd__o21ba_1
XFILLER_100_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08652_ _09508_/A _09233_/B _09074_/B _09206_/B vssd1 vssd1 vccd1 vccd1 _08654_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_81_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07603_ _07603_/A vssd1 vssd1 vccd1 vccd1 _14082_/D sky130_fd_sc_hd__clkbuf_1
X_08583_ _08637_/A _08582_/C _08578_/Y vssd1 vssd1 vccd1 vccd1 _08584_/C sky130_fd_sc_hd__a21bo_1
XFILLER_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13632__A _13644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07534_ _07534_/A _07534_/B vssd1 vssd1 vccd1 vccd1 _07534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07630__A _14125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07465_ _14197_/Q _14199_/Q _07469_/S vssd1 vssd1 vccd1 vccd1 _07466_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12248__A _12251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09204_ _09148_/B _09148_/C _09148_/A vssd1 vssd1 vccd1 vccd1 _09205_/C sky130_fd_sc_hd__o21bai_1
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07396_ _14209_/Q _14211_/Q _07415_/S vssd1 vssd1 vccd1 vccd1 _07396_/X sky130_fd_sc_hd__mux2_1
X_09135_ _09135_/A _09135_/B vssd1 vssd1 vccd1 vccd1 _09137_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10991__A _11082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ _09065_/B _09065_/C _09065_/A vssd1 vssd1 vccd1 vccd1 _09067_/C sky130_fd_sc_hd__a21o_1
X_08017_ _09821_/A vssd1 vssd1 vccd1 vccd1 _08284_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_2_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10215__B _10215_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09968_ _09968_/A _09968_/B vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08919_ _08919_/A _08919_/B vssd1 vssd1 vccd1 vccd1 _08953_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09553__B_N _09594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09899_ _09986_/A _09986_/B vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__xor2_1
XFILLER_94_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11930_ _12933_/A vssd1 vssd1 vccd1 vccd1 _12216_/A sky130_fd_sc_hd__buf_2
XFILLER_40_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _11861_/A vssd1 vssd1 vccd1 vccd1 _11861_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ input79/X _14425_/Q _13611_/S vssd1 vssd1 vccd1 vccd1 _13601_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _13938_/Q _10812_/B vssd1 vssd1 vccd1 vccd1 _10813_/B sky130_fd_sc_hd__or2_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _11823_/A vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13531_ _13531_/A vssd1 vssd1 vccd1 vccd1 _14404_/D sky130_fd_sc_hd__clkbuf_1
X_10743_ _10743_/A vssd1 vssd1 vccd1 vccd1 _10744_/A sky130_fd_sc_hd__buf_2
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13462_ _13462_/A vssd1 vssd1 vccd1 vccd1 _14385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10674_ _10674_/A vssd1 vssd1 vccd1 vccd1 _10761_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA_input95_A io_wbs_datwr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12413_ _12415_/A vssd1 vssd1 vccd1 vccd1 _12413_/Y sky130_fd_sc_hd__inv_2
X_13393_ _13393_/A vssd1 vssd1 vccd1 vccd1 _14365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12344_ _12347_/A vssd1 vssd1 vccd1 vccd1 _12344_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12275_ _12279_/A vssd1 vssd1 vccd1 vccd1 _12275_/Y sky130_fd_sc_hd__inv_2
X_14014_ _14304_/CLK _14014_/D vssd1 vssd1 vccd1 vccd1 _14014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11226_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11324_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07197__A1 _14094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11157_ _10715_/A _11152_/X _11153_/X _10744_/X _11156_/X vssd1 vssd1 vccd1 vccd1
+ _11253_/A sky130_fd_sc_hd__a221oi_4
XFILLER_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06944__A1 _14317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10108_ _10052_/B _10351_/B vssd1 vssd1 vccd1 vccd1 _10108_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11088_ _10700_/X _10987_/A _10987_/B vssd1 vssd1 vccd1 vccd1 _11089_/B sky130_fd_sc_hd__o21a_1
XFILLER_23_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10039_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10039_/X sky130_fd_sc_hd__or2_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13729_ _13729_/A _13729_/B vssd1 vssd1 vccd1 vccd1 _13730_/A sky130_fd_sc_hd__and2_1
XFILLER_108_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07121__A1 _07090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09661__A3 _10613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07250_ _14263_/Q _07249_/X _07253_/S vssd1 vssd1 vccd1 vccd1 _07251_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14287__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07181_ _07181_/A vssd1 vssd1 vccd1 vccd1 _14283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11508__A1 _11058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09822_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09826_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13627__A _13680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09753_ _08280_/A _08280_/B _08277_/A vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__o21a_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06965_ _06934_/X _06964_/X _14378_/Q vssd1 vssd1 vccd1 vccd1 _06966_/S sky130_fd_sc_hd__o21a_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08704_ _09241_/B _09000_/B _09152_/B _09241_/A vssd1 vssd1 vccd1 vccd1 _08706_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09684_ _09684_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09685_/B sky130_fd_sc_hd__nor2_1
X_06896_ _14413_/Q _07085_/A _14445_/Q vssd1 vssd1 vccd1 vccd1 _06896_/X sky130_fd_sc_hd__and3b_1
XFILLER_67_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08635_ _08998_/A _08634_/C _08630_/Y vssd1 vssd1 vccd1 vccd1 _08636_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__09840__A _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08566_ _08566_/A _08566_/B _08566_/C vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__nand3_1
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08456__A _08980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07517_ hold27/X _14179_/Q _07517_/S vssd1 vssd1 vccd1 vccd1 _07518_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08497_ _09870_/A vssd1 vssd1 vccd1 vccd1 _08893_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__07112__A1 _14263_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07448_ _14200_/Q _14202_/Q _07469_/S vssd1 vssd1 vccd1 vccd1 _07449_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14283_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07379_ _07491_/A vssd1 vssd1 vccd1 vccd1 _07379_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _09118_/A vssd1 vssd1 vccd1 vccd1 _09118_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08191__A _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ _10391_/B _10391_/C _10391_/A vssd1 vssd1 vccd1 vccd1 _10392_/A sky130_fd_sc_hd__a21oi_1
X_09049_ _09049_/A _09049_/B vssd1 vssd1 vccd1 vccd1 _09188_/C sky130_fd_sc_hd__nor2_1
XFILLER_89_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ _12060_/A vssd1 vssd1 vccd1 vccd1 _12060_/X sky130_fd_sc_hd__buf_2
XFILLER_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07179__A1 _14099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11011_ _11240_/A _11011_/B vssd1 vssd1 vccd1 vccd1 _11012_/B sky130_fd_sc_hd__or2_1
XANTENNA__06926__A1 _06894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__A _12441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12962_ _12966_/A vssd1 vssd1 vccd1 vccd1 _12962_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input10_A dout1[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11913_ hold5/X _11913_/B vssd1 vssd1 vccd1 vccd1 _13759_/D sky130_fd_sc_hd__nor2_1
XANTENNA__10486__A1 _09188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _14145_/Q _12885_/X _12891_/X _12892_/X vssd1 vssd1 vccd1 vccd1 _14145_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11844_ _14340_/Q _11833_/X _11834_/X _13799_/Q _11843_/X vssd1 vssd1 vccd1 vccd1
+ _11844_/X sky130_fd_sc_hd__a221o_1
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _12762_/B input59/X _11767_/B vssd1 vssd1 vccd1 vccd1 _12951_/B sky130_fd_sc_hd__or3b_4
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _12681_/X _14401_/Q _13522_/S vssd1 vssd1 vccd1 vccd1 _13515_/B sky130_fd_sc_hd__mux2_1
X_10726_ _11216_/A _10748_/B vssd1 vssd1 vccd1 vccd1 _10727_/D sky130_fd_sc_hd__xnor2_1
XFILLER_16_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13445_ _13445_/A vssd1 vssd1 vccd1 vccd1 _14380_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10657_ _10826_/A _10705_/B _11110_/A _10652_/X vssd1 vssd1 vccd1 vccd1 _10657_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09197__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13376_ _13376_/A vssd1 vssd1 vccd1 vccd1 _14360_/D sky130_fd_sc_hd__clkbuf_1
X_10588_ _10588_/A _10588_/B vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__or2_1
X_12327_ _12329_/A vssd1 vssd1 vccd1 vccd1 _12327_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12258_ _12259_/A vssd1 vssd1 vccd1 vccd1 _12258_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13447__A _13447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ _11302_/A _11302_/B vssd1 vssd1 vccd1 vccd1 _11312_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12189_ _13209_/A vssd1 vssd1 vccd1 vccd1 _13037_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__06917__A1 _14288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09660__A _09660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08420_ _08595_/A vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__buf_6
XFILLER_52_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08351_ _09361_/A _09361_/B _09473_/B _09844_/A vssd1 vssd1 vccd1 vccd1 _09555_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_32_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07302_ _07312_/B vssd1 vssd1 vccd1 vccd1 _07471_/A sky130_fd_sc_hd__buf_2
X_08282_ _08580_/A vssd1 vssd1 vccd1 vccd1 _08632_/A sky130_fd_sc_hd__buf_6
XFILLER_20_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07233_ _14268_/Q _07232_/X _07236_/S vssd1 vssd1 vccd1 vccd1 _07234_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07164_ _14103_/Q _07140_/X _07143_/X vssd1 vssd1 vccd1 vccd1 _07164_/X sky130_fd_sc_hd__a21o_2
XFILLER_118_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07095_ _14441_/Q _14265_/Q vssd1 vssd1 vccd1 vccd1 _07095_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13357__A _13411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07355__A _14101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _10036_/B vssd1 vssd1 vccd1 vccd1 _10122_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_input2_A dout1[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07997_ _09084_/A _09084_/B _08976_/A _09058_/B vssd1 vssd1 vccd1 vccd1 _07997_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_86_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07074__B _07098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06948_ _14284_/Q _06929_/X _06947_/X _14380_/Q vssd1 vssd1 vccd1 vccd1 _06948_/X
+ sky130_fd_sc_hd__o211a_1
X_09736_ _09739_/B _09739_/C _09739_/A vssd1 vssd1 vccd1 vccd1 _09742_/A sky130_fd_sc_hd__a21oi_2
XFILLER_28_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09667_ _09667_/A vssd1 vssd1 vccd1 vccd1 _09667_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06879_ _14269_/Q _06873_/X _06878_/X _14365_/Q vssd1 vssd1 vccd1 vccd1 _06879_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_43_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13092__A _13411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ _08619_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _08618_/X sky130_fd_sc_hd__or2_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08186__A _09584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _09681_/A _09598_/B vssd1 vssd1 vccd1 vccd1 _09676_/A sky130_fd_sc_hd__xnor2_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07090__A _07090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08549_ _08571_/A _09943_/B _08783_/A _08128_/B vssd1 vssd1 vccd1 vccd1 _08550_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09086__B2 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11560_ _14045_/Q _13957_/Q vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__and2_1
XFILLER_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10511_ _10597_/A _10511_/B _10511_/C vssd1 vssd1 vccd1 vccd1 _10511_/X sky130_fd_sc_hd__and3_1
XANTENNA__10640__A1 _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ _11007_/B _11489_/X _11475_/X _11291_/A _11490_/X vssd1 vssd1 vccd1 vccd1
+ _11491_/X sky130_fd_sc_hd__o221a_1
XFILLER_52_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13230_ _13526_/A vssd1 vssd1 vccd1 vccd1 _13230_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10442_ _10472_/S _10471_/A vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__xnor2_1
XFILLER_100_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13161_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13161_/Y sky130_fd_sc_hd__inv_2
X_10373_ _10326_/A _10373_/B vssd1 vssd1 vccd1 vccd1 _10588_/A sky130_fd_sc_hd__and2b_1
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12112_ _12936_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12112_/X sky130_fd_sc_hd__or2_1
XANTENNA__11994__B _12952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input58_A io_wbs_adr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_46_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12043_ _13795_/Q _12038_/X _12039_/X _13811_/Q vssd1 vssd1 vccd1 vccd1 _12044_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_0_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_38_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13994_ _14442_/CLK _13994_/D vssd1 vssd1 vccd1 vccd1 _13994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12945_ _12973_/A vssd1 vssd1 vccd1 vccd1 _12950_/A sky130_fd_sc_hd__buf_2
XFILLER_80_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12919_/A _12883_/B vssd1 vssd1 vccd1 vccd1 _12876_/X sky130_fd_sc_hd__or2_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_75_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_2_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11234__B _11285_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _14333_/Q _11808_/X _11823_/X _13792_/Q _11826_/X vssd1 vssd1 vccd1 vccd1
+ _11827_/X sky130_fd_sc_hd__a221o_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07088__B1 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11758_ input45/X input48/X input47/X input50/X vssd1 vssd1 vccd1 vccd1 _11759_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_53_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08824__A _08983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ _10828_/B _10709_/B vssd1 vssd1 vccd1 vccd1 _10832_/A sky130_fd_sc_hd__nand2_1
X_11689_ _13765_/Q _13764_/Q _13763_/Q vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__or3_1
X_13428_ _13428_/A vssd1 vssd1 vccd1 vccd1 _13504_/A sky130_fd_sc_hd__clkbuf_4
X_13359_ _13359_/A _13525_/A vssd1 vssd1 vccd1 vccd1 _13447_/A sky130_fd_sc_hd__or2_4
XFILLER_115_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07920_ _07920_/A vssd1 vssd1 vccd1 vccd1 _13971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07851_ _14034_/Q _13980_/Q vssd1 vssd1 vccd1 vccd1 _07881_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07563__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 dout1[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_07782_ _10900_/B vssd1 vssd1 vccd1 vccd1 _10895_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09521_ _09527_/A vssd1 vssd1 vccd1 vccd1 _09521_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09452_ _09471_/A _09471_/B _09471_/C vssd1 vssd1 vccd1 vccd1 _09452_/X sky130_fd_sc_hd__and3_1
XFILLER_92_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08403_ _08403_/A _08403_/B vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__or2_1
XFILLER_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09383_ _09553_/C _09074_/B _09287_/X _09286_/X _09873_/A vssd1 vssd1 vccd1 vccd1
+ _09385_/B sky130_fd_sc_hd__a32o_1
XANTENNA__07079__B1 _07048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ _09336_/A _08334_/B vssd1 vssd1 vccd1 vccd1 _08335_/B sky130_fd_sc_hd__and2_1
XFILLER_36_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08265_ _08226_/A _08265_/B vssd1 vssd1 vccd1 vccd1 _08266_/B sky130_fd_sc_hd__and2b_1
XFILLER_119_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12256__A _12259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07216_ _14273_/Q _07215_/X _07219_/S vssd1 vssd1 vccd1 vccd1 _07217_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08196_ _08317_/A _09999_/A _08131_/B _08130_/A vssd1 vssd1 vccd1 vccd1 _08198_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13572__A0 _12681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07147_ _13951_/Q _07203_/A _07146_/Y _14058_/Q vssd1 vssd1 vccd1 vccd1 _07150_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07078_ _14443_/Q _14267_/Q vssd1 vssd1 vccd1 vccd1 _07078_/Y sky130_fd_sc_hd__nand2_1
XFILLER_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10620__B1_N _09273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07085__A _07085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07554__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09719_ _09715_/A _09715_/C _09715_/B vssd1 vssd1 vccd1 vccd1 _09720_/B sky130_fd_sc_hd__o21ai_1
XFILLER_56_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10991_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11083_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12734_/A vssd1 vssd1 vccd1 vccd1 _12730_/Y sky130_fd_sc_hd__inv_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12660_/X _14048_/Q _12665_/S vssd1 vssd1 vccd1 vccd1 _12662_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09059__A1 _09508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09059__B2 _08445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14400_ _14400_/CLK _14400_/D vssd1 vssd1 vccd1 vccd1 _14400_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11612_/A vssd1 vssd1 vccd1 vccd1 _13851_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12592_/A vssd1 vssd1 vccd1 vccd1 _14030_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14331_ _14396_/CLK _14331_/D vssd1 vssd1 vccd1 vccd1 _14331_/Q sky130_fd_sc_hd__dfxtp_1
X_11543_ _14050_/Q _13962_/Q vssd1 vssd1 vccd1 vccd1 _11543_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12166__A input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14262_ _14365_/CLK _14262_/D _13119_/Y vssd1 vssd1 vccd1 vccd1 _14262_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_52_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11474_ _11474_/A _11533_/S vssd1 vssd1 vccd1 vccd1 _11499_/A sky130_fd_sc_hd__nand2_2
XFILLER_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13563__A0 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13213_ _14324_/Q _13196_/X _13212_/X _13053_/X vssd1 vssd1 vccd1 vccd1 _14324_/D
+ sky130_fd_sc_hd__o211a_1
X_10425_ _10440_/A _10425_/B vssd1 vssd1 vccd1 vccd1 _10443_/S sky130_fd_sc_hd__xor2_2
X_14193_ _14224_/CLK _14193_/D _12983_/Y vssd1 vssd1 vccd1 vccd1 _14193_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13144_ _13146_/A vssd1 vssd1 vccd1 vccd1 _13144_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10356_ _10380_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10358_/A sky130_fd_sc_hd__xor2_2
XFILLER_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output164_A _14319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _13075_/A vssd1 vssd1 vccd1 vccd1 _14244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10287_ _10311_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10288_/B sky130_fd_sc_hd__xor2_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12026_ _12026_/A _12026_/B vssd1 vssd1 vccd1 vccd1 _12027_/A sky130_fd_sc_hd__and2_1
XFILLER_39_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12826__C1 _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13977_ _14107_/CLK _13977_/D _12403_/Y vssd1 vssd1 vccd1 vccd1 _13977_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12928_ _12928_/A vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10852__A1 _10845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12859_ _12898_/B vssd1 vssd1 vccd1 vccd1 _12870_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08554__A _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11801__B1 _11800_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ _08146_/A _08050_/B vssd1 vssd1 vccd1 vccd1 _08051_/B sky130_fd_sc_hd__nand2_1
X_07001_ _14421_/Q _07000_/Y _06970_/X vssd1 vssd1 vccd1 vccd1 _07001_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07233__A0 _14268_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08952_ _08935_/Y _08942_/Y _08948_/X _08951_/X vssd1 vssd1 vccd1 vccd1 _08952_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07903_ _07901_/Y _07902_/X _07890_/A _13975_/Q vssd1 vssd1 vccd1 vccd1 _13975_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_08883_ _08883_/A _08883_/B _08883_/C vssd1 vssd1 vccd1 vccd1 _08885_/A sky130_fd_sc_hd__or3_1
XFILLER_69_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13635__A _13644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _07834_/A _07834_/B vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07765_ _14060_/Q _07764_/X _07765_/S vssd1 vssd1 vccd1 vccd1 _07766_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _09514_/A _09465_/B _09464_/A vssd1 vssd1 vccd1 vccd1 _09516_/A sky130_fd_sc_hd__o21ai_2
X_07696_ _14141_/Q _07665_/Y _07732_/A _14142_/Q _07695_/X vssd1 vssd1 vccd1 vccd1
+ _07696_/X sky130_fd_sc_hd__o221a_1
XFILLER_25_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09435_ _09435_/A _09435_/B vssd1 vssd1 vccd1 vccd1 _09437_/B sky130_fd_sc_hd__xnor2_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10994__A _11079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ _09281_/B _09281_/C _09281_/A vssd1 vssd1 vccd1 vccd1 _09367_/C sky130_fd_sc_hd__a21bo_1
XFILLER_40_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_42_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14457_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_08317_ _08317_/A _09962_/B vssd1 vssd1 vccd1 vccd1 _08318_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09297_ _09297_/A _09818_/A vssd1 vssd1 vccd1 vccd1 _09299_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ _09762_/B _09786_/A _08211_/B _08208_/X vssd1 vssd1 vccd1 vccd1 _09755_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_119_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_1_0_0_io_wbs_clk_A clkbuf_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08179_ _09402_/A vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10210_ _10211_/A _10211_/B vssd1 vssd1 vccd1 vccd1 _10213_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07224__A0 _14271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11190_ _10735_/X _11151_/X _11153_/X _10975_/A vssd1 vssd1 vccd1 vccd1 _11190_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12195__B_N input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09764__A2 _09088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12433__B _12952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _10141_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10141_/X sky130_fd_sc_hd__or2b_1
XFILLER_106_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10072_ _09922_/Y _10033_/Y _10034_/Y vssd1 vssd1 vccd1 vccd1 _10330_/B sky130_fd_sc_hd__a21oi_2
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12520__A1 _08946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ _13905_/CLK _13900_/D _12308_/Y vssd1 vssd1 vccd1 vccd1 _13900_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__13545__A _13634_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10531__B1 _10528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13831_ _14258_/CLK _13831_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__14020__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10974_ _11020_/B _11021_/A vssd1 vssd1 vccd1 vccd1 _11016_/B sky130_fd_sc_hd__nand2_1
X_13762_ _13820_/CLK _13762_/D _11953_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ _12715_/A vssd1 vssd1 vccd1 vccd1 _12713_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13693_ _13693_/A vssd1 vssd1 vccd1 vccd1 _14451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12644_ _12644_/A vssd1 vssd1 vccd1 vccd1 _14044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12587__A1 _14029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12575_ _12909_/A _14026_/Q _12583_/S vssd1 vssd1 vccd1 vccd1 _12576_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08093__B _09319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14314_ _14453_/CLK _14314_/D _13183_/Y vssd1 vssd1 vccd1 vccd1 _14314_/Q sky130_fd_sc_hd__dfrtp_4
X_11526_ _11521_/A _11525_/Y _11464_/X vssd1 vssd1 vccd1 vccd1 _11526_/X sky130_fd_sc_hd__a21o_1
XFILLER_102_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14245_ _14250_/CLK _14245_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10843__S _10871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _11457_/A vssd1 vssd1 vccd1 vccd1 _11457_/Y sky130_fd_sc_hd__inv_2
X_10408_ _10407_/A _10414_/S _10361_/A vssd1 vssd1 vccd1 vccd1 _10413_/B sky130_fd_sc_hd__a21o_1
X_14176_ _14179_/CLK _14176_/D _12962_/Y vssd1 vssd1 vccd1 vccd1 _14176_/Q sky130_fd_sc_hd__dfrtp_1
X_11388_ hold28/X _11390_/B vssd1 vssd1 vccd1 vccd1 _11388_/X sky130_fd_sc_hd__or2_1
XFILLER_98_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13127_ _13128_/A vssd1 vssd1 vccd1 vccd1 _13127_/Y sky130_fd_sc_hd__inv_2
X_10339_ _10310_/A _10310_/B _10338_/Y vssd1 vssd1 vccd1 vccd1 _10347_/B sky130_fd_sc_hd__a21o_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _14239_/Q _13041_/A _13057_/X _13053_/X vssd1 vssd1 vccd1 vccd1 _14239_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09507__A2 _08097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12009_ _12009_/A vssd1 vssd1 vccd1 vccd1 _13785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07550_ _14256_/Q vssd1 vssd1 vccd1 vccd1 _07595_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07481_ _07348_/A _07479_/X _07480_/X _07462_/X _14195_/Q vssd1 vssd1 vccd1 vccd1
+ _14195_/D sky130_fd_sc_hd__a32o_1
XANTENNA__13190__A _13193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ _09295_/A _09220_/B _09220_/C vssd1 vssd1 vccd1 vccd1 _09223_/A sky130_fd_sc_hd__or3_2
XFILLER_22_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13224__C1 _13053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08284__A _08632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09151_ _09151_/A _09151_/B _09151_/C vssd1 vssd1 vccd1 vccd1 _09158_/A sky130_fd_sc_hd__nand3_1
XFILLER_33_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10319__A _10393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ _09348_/B vssd1 vssd1 vccd1 vccd1 _09233_/B sky130_fd_sc_hd__buf_2
X_09082_ _09081_/B _09081_/C _09081_/A vssd1 vssd1 vccd1 vccd1 _09083_/B sky130_fd_sc_hd__a21oi_1
X_08033_ _14017_/Q vssd1 vssd1 vccd1 vccd1 _09378_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput60 io_wbs_adr[5] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_2
Xinput71 io_wbs_datwr[14] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_2
Xinput82 io_wbs_datwr[24] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_2
Xinput93 io_wbs_datwr[5] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_4
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09984_ _09984_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _10268_/A sky130_fd_sc_hd__xnor2_2
XFILLER_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08935_ _08935_/A _08935_/B vssd1 vssd1 vccd1 vccd1 _08935_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08866_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08897_/A sky130_fd_sc_hd__xnor2_2
XFILLER_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07363__A _07363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07817_ _14036_/Q _13982_/Q vssd1 vssd1 vccd1 vccd1 _07872_/A sky130_fd_sc_hd__nor2_1
X_08797_ _08797_/A _08797_/B vssd1 vssd1 vccd1 vccd1 _08798_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08178__B _10302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07748_ _14154_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07748_/X sky130_fd_sc_hd__and2_1
XFILLER_77_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ _07679_/A _07679_/B vssd1 vssd1 vccd1 vccd1 _07687_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09418_ _09263_/X _09415_/Y _09416_/Y _09417_/X vssd1 vssd1 vccd1 vccd1 _09420_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_41_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10690_ _13984_/Q _11533_/S _10690_/S vssd1 vssd1 vccd1 vccd1 _10691_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12428__B _12900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12569__A1 _14024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09349_ _09349_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09351_/B sky130_fd_sc_hd__nand2_1
X_12360_ _12360_/A vssd1 vssd1 vccd1 vccd1 _12360_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11311_ _11305_/Y _11311_/B vssd1 vssd1 vccd1 vccd1 _11312_/C sky130_fd_sc_hd__and2b_1
X_12291_ _12291_/A vssd1 vssd1 vccd1 vccd1 _12291_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14030_ _14031_/CLK _14030_/D vssd1 vssd1 vccd1 vccd1 _14030_/Q sky130_fd_sc_hd__dfxtp_4
X_11242_ _11279_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11336_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11173_ _13917_/Q _13918_/Q _13919_/Q _13920_/Q _10967_/S _10676_/A vssd1 vssd1 vccd1
+ vccd1 _11173_/X sky130_fd_sc_hd__mux4_2
XFILLER_45_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10124_ _10214_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _10124_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_input40_A io_wbs_adr[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10055_ _10055_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _10112_/B sky130_fd_sc_hd__xnor2_2
XFILLER_57_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08211__A_N _08208_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_14_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_90_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13814_ _13826_/CLK _13814_/D vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13745_ _13745_/A _13745_/B vssd1 vssd1 vccd1 vccd1 _13746_/A sky130_fd_sc_hd__and2_1
X_10957_ _13904_/Q _13905_/Q _13906_/Q _13907_/Q _10946_/B _10954_/A vssd1 vssd1 vccd1
+ vccd1 _10957_/X sky130_fd_sc_hd__mux4_2
XFILLER_95_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10838__S _10871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__A1 _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ _13676_/A vssd1 vssd1 vccd1 vccd1 _14446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10888_ _10888_/A vssd1 vssd1 vccd1 vccd1 _13932_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11242__B _11279_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12627_ _12218_/X _14040_/Q _12642_/S vssd1 vssd1 vccd1 vccd1 _12628_/B sky130_fd_sc_hd__mux2_1
XFILLER_106_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12558_ _12938_/A _09762_/B _12562_/S vssd1 vssd1 vccd1 vccd1 _12559_/B sky130_fd_sc_hd__mux2_1
XFILLER_117_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ _10215_/B _11486_/X _11507_/Y _11508_/X vssd1 vssd1 vccd1 vccd1 _13865_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09647__B _09652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12489_ _14000_/Q _12481_/X _12488_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _14000_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14228_ _14256_/CLK _14228_/D _13026_/Y vssd1 vssd1 vccd1 vccd1 _14228_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__07739__A1 _14068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _14164_/CLK _14159_/D vssd1 vssd1 vccd1 vccd1 _14159_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _14424_/Q _06981_/B _14456_/Q vssd1 vssd1 vccd1 vccd1 _06981_/X sky130_fd_sc_hd__and3b_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _08723_/A _08723_/C _08723_/B vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__a21bo_1
XFILLER_79_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08651_ _08982_/A _09842_/A vssd1 vssd1 vccd1 vccd1 _08654_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07602_ _14082_/Q input29/X _07604_/S vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08582_ _08578_/Y _08637_/A _08582_/C vssd1 vssd1 vccd1 vccd1 _08637_/B sky130_fd_sc_hd__nand3b_1
XFILLER_19_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07533_ _14173_/Q _14172_/Q _14171_/Q _14174_/Q vssd1 vssd1 vccd1 vccd1 _07533_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07464_ _07464_/A vssd1 vssd1 vccd1 vccd1 _07483_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09203_ _08312_/A _09011_/B _09202_/A _09202_/C vssd1 vssd1 vccd1 vccd1 _09205_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07395_ _14093_/Q _07363_/A vssd1 vssd1 vccd1 vccd1 _07395_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09134_ _09134_/A _09834_/A vssd1 vssd1 vccd1 vccd1 _09135_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ _09065_/A _09065_/B _09065_/C vssd1 vssd1 vccd1 vccd1 _09067_/B sky130_fd_sc_hd__nand3_2
XFILLER_118_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08016_ _13875_/Q vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08927__B1 _08783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07327__B_N _07323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09967_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09970_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08918_ _08944_/C _08918_/B vssd1 vssd1 vccd1 vccd1 _08919_/B sky130_fd_sc_hd__nand2_1
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09898_ _10191_/A _09902_/B _09897_/X vssd1 vssd1 vccd1 vccd1 _09986_/B sky130_fd_sc_hd__a21oi_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08189__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08849_ _08849_/A _08849_/B _08849_/C vssd1 vssd1 vccd1 vccd1 _08883_/A sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_5_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _14350_/Q _11864_/B vssd1 vssd1 vccd1 vccd1 _11861_/A sky130_fd_sc_hd__and2_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07821__A _14032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10811_ _10858_/B _10858_/C _10858_/A vssd1 vssd1 vccd1 vccd1 _10853_/C sky130_fd_sc_hd__a21oi_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _11791_/A vssd1 vssd1 vccd1 vccd1 _11791_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12439__A _12486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13530_ _13539_/A _13530_/B vssd1 vssd1 vccd1 vccd1 _13531_/A sky130_fd_sc_hd__and2_1
X_10742_ _13950_/Q _13949_/Q vssd1 vssd1 vccd1 vccd1 _10743_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11462__B2 _11092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10673_ _10954_/A _11171_/S vssd1 vssd1 vccd1 vccd1 _10674_/A sky130_fd_sc_hd__or2_1
X_13461_ _13461_/A _13461_/B vssd1 vssd1 vccd1 vccd1 _13462_/A sky130_fd_sc_hd__and2_1
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09407__A1 _09404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12412_ _12415_/A vssd1 vssd1 vccd1 vccd1 _12412_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input88_A io_wbs_datwr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ _13392_/A _13392_/B vssd1 vssd1 vccd1 vccd1 _13393_/A sky130_fd_sc_hd__and2_1
XFILLER_51_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08652__A _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12343_ _12347_/A vssd1 vssd1 vccd1 vccd1 _12343_/Y sky130_fd_sc_hd__inv_2
X_12274_ _12286_/A vssd1 vssd1 vccd1 vccd1 _12279_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11225_ _11225_/A _11225_/B vssd1 vssd1 vccd1 vccd1 _11291_/B sky130_fd_sc_hd__xnor2_2
XFILLER_5_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14013_ _14304_/CLK _14013_/D vssd1 vssd1 vccd1 vccd1 _14013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11156_ _10722_/B _11154_/X _11155_/X _10730_/B vssd1 vssd1 vccd1 vccd1 _11156_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10107_ _10280_/B _10121_/B vssd1 vssd1 vccd1 vccd1 _10120_/B sky130_fd_sc_hd__nand2_1
XFILLER_110_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11087_ _11142_/B _11087_/B vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__xnor2_2
X_10038_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10067_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07495__C_N _07452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11989_ _12001_/B vssd1 vssd1 vccd1 vccd1 _11990_/B sky130_fd_sc_hd__buf_2
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13728_ input84/X _14462_/Q _13738_/S vssd1 vssd1 vccd1 vccd1 _13729_/B sky130_fd_sc_hd__mux2_1
XFILLER_56_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13659_ _13659_/A vssd1 vssd1 vccd1 vccd1 _14441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07180_ _14283_/Q _07179_/X _07183_/S vssd1 vssd1 vccd1 vccd1 _07181_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10010__A1_N _09895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09821_ _09821_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__xor2_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09752_ _08412_/Y _10524_/B _09750_/Y _09751_/Y vssd1 vssd1 vccd1 vccd1 _10515_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ _14426_/Q _06981_/B _14458_/Q vssd1 vssd1 vccd1 vccd1 _06964_/X sky130_fd_sc_hd__and3b_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _09134_/A _08703_/B vssd1 vssd1 vccd1 vccd1 _08707_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06895_ _07105_/A vssd1 vssd1 vccd1 vccd1 _07085_/A sky130_fd_sc_hd__clkbuf_4
X_09683_ _09683_/A _09683_/B _09683_/C vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__and3_1
XFILLER_39_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ _08630_/Y _08998_/A _08634_/C vssd1 vssd1 vccd1 vccd1 _08998_/B sky130_fd_sc_hd__nand3b_1
XFILLER_27_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08537_/A _08534_/C _08534_/A vssd1 vssd1 vccd1 vccd1 _08566_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12259__A _12259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08456__B _08767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ _07516_/A vssd1 vssd1 vccd1 vccd1 _14180_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11444__A1 _11082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08496_ _09865_/A vssd1 vssd1 vccd1 vccd1 _09870_/A sky130_fd_sc_hd__buf_4
XFILLER_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07112__A2 _07085_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07447_ _14227_/Q vssd1 vssd1 vccd1 vccd1 _07469_/S sky130_fd_sc_hd__clkbuf_2
X_07378_ _14213_/Q _14215_/Q _07387_/S vssd1 vssd1 vccd1 vccd1 _07378_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09117_ _10632_/B _10631_/A vssd1 vssd1 vccd1 vccd1 _09117_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09048_ _09048_/A _09048_/B _09048_/C vssd1 vssd1 vccd1 vccd1 _09049_/B sky130_fd_sc_hd__and3_1
XFILLER_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _11067_/B _11010_/B vssd1 vssd1 vccd1 vccd1 _11107_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11904__C1 _11874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07816__A _14037_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12961_ _12973_/A vssd1 vssd1 vccd1 vccd1 _12966_/A sky130_fd_sc_hd__buf_2
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09876__A1 _08494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11912_ _13819_/Q _11872_/A _11911_/Y _11914_/B vssd1 vssd1 vccd1 vccd1 _11913_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_73_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _12920_/A vssd1 vssd1 vccd1 vccd1 _12892_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _14005_/Q _11845_/B vssd1 vssd1 vccd1 vccd1 _11843_/X sky130_fd_sc_hd__and2_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12169__A input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11774_ _11774_/A _11774_/B _11774_/C vssd1 vssd1 vccd1 vccd1 _12762_/B sky130_fd_sc_hd__or3_2
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13513_/A vssd1 vssd1 vccd1 vccd1 _14400_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10725_ _10951_/A _11158_/S _10967_/S _10676_/A vssd1 vssd1 vccd1 vccd1 _10748_/B
+ sky130_fd_sc_hd__or4b_4
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13444_ _13444_/A _13444_/B vssd1 vssd1 vccd1 vccd1 _13445_/A sky130_fd_sc_hd__and2_1
X_10656_ _11100_/A vssd1 vssd1 vccd1 vccd1 _11110_/A sky130_fd_sc_hd__buf_2
X_13375_ _13375_/A _13375_/B vssd1 vssd1 vccd1 vccd1 _13376_/A sky130_fd_sc_hd__and2_1
X_10587_ _10587_/A _10598_/C vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__nor2_1
X_12326_ _12329_/A vssd1 vssd1 vccd1 vccd1 _12326_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12257_ _12259_/A vssd1 vssd1 vccd1 vccd1 _12257_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11208_ _11208_/A _11208_/B vssd1 vssd1 vccd1 vccd1 _11302_/B sky130_fd_sc_hd__xnor2_2
X_12188_ _12211_/A input65/X vssd1 vssd1 vccd1 vccd1 _13209_/A sky130_fd_sc_hd__and2b_2
XFILLER_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06917__A2 _06873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__A2 _11872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _11140_/B _11138_/X _11184_/S vssd1 vssd1 vccd1 vccd1 _11139_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09941__A _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11123__B1 _11100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09867__A1 _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13463__A _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09660__B _10604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14254__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08350_ _13866_/Q vssd1 vssd1 vccd1 vccd1 _09844_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07301_ _07313_/C vssd1 vssd1 vccd1 vccd1 _07301_/Y sky130_fd_sc_hd__inv_2
X_08281_ _09749_/B _09749_/C _09749_/A vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__o21ai_2
XFILLER_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11711__A _11920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07232_ _14084_/Q _13884_/Q _07235_/S vssd1 vssd1 vccd1 vccd1 _07232_/X sky130_fd_sc_hd__mux2_2
XFILLER_118_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07163_ _07163_/A vssd1 vssd1 vccd1 vccd1 _14288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ _07094_/A vssd1 vssd1 vccd1 vccd1 _14298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07030__A1 _14306_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09804_ _09804_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _10036_/B sky130_fd_sc_hd__xnor2_4
XFILLER_75_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07996_ _13870_/Q vssd1 vssd1 vccd1 vccd1 _09058_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09851__A _09895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _09735_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__or2_1
X_06947_ _14428_/Q _06946_/Y _06931_/X vssd1 vssd1 vccd1 vccd1 _06947_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09858__A1 _08703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09666_ _09666_/A _10576_/B vssd1 vssd1 vccd1 vccd1 _09666_/X sky130_fd_sc_hd__or2_1
XANTENNA__08467__A _08828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06878_ _14413_/Q _06874_/Y _06877_/X vssd1 vssd1 vccd1 vccd1 _06878_/X sky130_fd_sc_hd__a21o_1
X_08617_ _08617_/A _08738_/A vssd1 vssd1 vccd1 vccd1 _08964_/A sky130_fd_sc_hd__nand2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09680_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09598_/B sky130_fd_sc_hd__xnor2_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12614__A0 _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ _08824_/C vssd1 vssd1 vccd1 vccd1 _09943_/B sky130_fd_sc_hd__buf_2
XFILLER_70_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09086__A2 _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07097__A1 _14265_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08479_ _09493_/B _09905_/B _09941_/B _09493_/A vssd1 vssd1 vccd1 vccd1 _08479_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_11_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12717__A _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10510_ _10508_/B _10520_/B _10506_/Y _10508_/A vssd1 vssd1 vccd1 vccd1 _10511_/C
+ sky130_fd_sc_hd__a211o_1
X_11490_ _11534_/S vssd1 vssd1 vccd1 vccd1 _11490_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ _09968_/A _10443_/S _10440_/X vssd1 vssd1 vccd1 vccd1 _10471_/A sky130_fd_sc_hd__o21a_1
XFILLER_108_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13160_ _13178_/A vssd1 vssd1 vccd1 vccd1 _13165_/A sky130_fd_sc_hd__buf_2
X_10372_ _10598_/A _10598_/B _10327_/X _10376_/A vssd1 vssd1 vccd1 vccd1 _10564_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_3_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ input69/X vssd1 vssd1 vccd1 vccd1 _12936_/A sky130_fd_sc_hd__buf_4
X_13091_ _13428_/A vssd1 vssd1 vccd1 vccd1 _13411_/A sky130_fd_sc_hd__buf_4
XFILLER_2_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12042_ _12042_/A vssd1 vssd1 vccd1 vccd1 _13794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09849__A1 _08836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13993_ _14441_/CLK _13993_/D vssd1 vssd1 vccd1 vccd1 _13993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12853__A0 _12654_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ _13010_/A vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12875_ _14138_/Q _12872_/X _12874_/X _12866_/X vssd1 vssd1 vccd1 vccd1 _14138_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _13998_/Q _11845_/B _12254_/B _14117_/Q vssd1 vssd1 vccd1 vccd1 _11826_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11757_ input49/X input52/X input51/X vssd1 vssd1 vccd1 vccd1 _11759_/C sky130_fd_sc_hd__or3_2
XFILLER_57_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08824__B _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10708_ _13942_/Q _10708_/B vssd1 vssd1 vccd1 vccd1 _10709_/B sky130_fd_sc_hd__or2_1
X_11688_ _11682_/B _11661_/X _11687_/Y vssd1 vssd1 vccd1 vccd1 _13775_/D sky130_fd_sc_hd__o21a_1
X_13427_ _13427_/A vssd1 vssd1 vccd1 vccd1 _14375_/D sky130_fd_sc_hd__clkbuf_1
X_10639_ _10639_/A _10639_/B vssd1 vssd1 vccd1 vccd1 _10639_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _13358_/A _13358_/B vssd1 vssd1 vccd1 vccd1 _13525_/A sky130_fd_sc_hd__nand2_4
XFILLER_6_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ _12310_/A vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__inv_2
X_13289_ _13332_/A vssd1 vssd1 vccd1 vccd1 _13289_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12362__A _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10147__A1 _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07850_ _07885_/B _07886_/B _07885_/A vssd1 vssd1 vccd1 vccd1 _07882_/A sky130_fd_sc_hd__o21ba_1
XFILLER_112_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07781_ _13988_/Q _13987_/Q _07786_/A vssd1 vssd1 vccd1 vccd1 _10900_/B sky130_fd_sc_hd__or3b_2
Xinput3 dout1[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13193__A _13193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09520_ _09454_/Y _09470_/X _09518_/Y _09519_/X vssd1 vssd1 vccd1 vccd1 _09527_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_65_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09451_ _09440_/A _09440_/B _09440_/C vssd1 vssd1 vccd1 vccd1 _09471_/C sky130_fd_sc_hd__a21o_1
XFILLER_91_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08402_ _09712_/A _08402_/B vssd1 vssd1 vccd1 vccd1 _08402_/X sky130_fd_sc_hd__or2_1
XFILLER_40_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09382_ _09441_/A _09382_/B _09382_/C vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__or3_1
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13794__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08333_ _08122_/X _08331_/Y _08391_/A _08330_/Y vssd1 vssd1 vccd1 vccd1 _08336_/B
+ sky130_fd_sc_hd__a211oi_1
Xclkbuf_leaf_32_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13946_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08264_ _09771_/A _08264_/B vssd1 vssd1 vccd1 vccd1 _08266_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07215_ _14089_/Q hold39/A _07218_/S vssd1 vssd1 vccd1 vccd1 _07215_/X sky130_fd_sc_hd__mux2_2
X_08195_ _08195_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08221_/C sky130_fd_sc_hd__or2_1
XFILLER_119_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09846__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _12205_/A _07146_/B vssd1 vssd1 vccd1 vccd1 _07146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07077_ _07077_/A vssd1 vssd1 vccd1 vccd1 _14300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07539__C1 _14192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09581__A _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13088__A0 _12633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _14020_/Q vssd1 vssd1 vccd1 vccd1 _09286_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09718_ _09718_/A _09717_/X vssd1 vssd1 vccd1 vccd1 _09718_/X sky130_fd_sc_hd__or2b_1
Xclkbuf_leaf_71_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14149_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__07813__B _07921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _10990_/A _10990_/B vssd1 vssd1 vccd1 vccd1 _11082_/B sky130_fd_sc_hd__xnor2_1
XFILLER_71_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09649_ _09651_/A _09647_/X _09640_/X _09638_/B vssd1 vssd1 vccd1 vccd1 _09649_/Y
+ sky130_fd_sc_hd__o211ai_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ input96/X vssd1 vssd1 vccd1 vccd1 _12660_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09059__A2 _09218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08925__A _08925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ hold13/A _11610_/Y _11611_/S vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12591_ _12594_/A _12591_/B vssd1 vssd1 vccd1 vccd1 _12592_/A sky130_fd_sc_hd__and2_1
X_14330_ _14396_/CLK _14330_/D vssd1 vssd1 vccd1 vccd1 _14330_/Q sky130_fd_sc_hd__dfxtp_1
X_11542_ _14051_/Q _13963_/Q vssd1 vssd1 vccd1 vccd1 _11609_/A sky130_fd_sc_hd__or2_1
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ _14281_/CLK _14261_/D _13118_/Y vssd1 vssd1 vccd1 vccd1 _14261_/Q sky130_fd_sc_hd__dfrtp_4
X_11473_ _11466_/A _11471_/X _11472_/X vssd1 vssd1 vccd1 vccd1 _11473_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input70_A io_wbs_datwr[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13212_ _14404_/Q _13199_/X _13205_/X _13211_/X vssd1 vssd1 vccd1 vccd1 _13212_/X
+ sky130_fd_sc_hd__a211o_1
X_10424_ _10394_/A _10394_/B _10423_/X vssd1 vssd1 vccd1 vccd1 _10425_/B sky130_fd_sc_hd__a21bo_1
X_14192_ _14244_/CLK _14192_/D _12982_/Y vssd1 vssd1 vccd1 vccd1 _14192_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13278__A _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13143_ _13146_/A vssd1 vssd1 vccd1 vccd1 _13143_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12182__A _12952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10355_ _10332_/A _10332_/B _10354_/X vssd1 vssd1 vccd1 vccd1 _10380_/B sky130_fd_sc_hd__a21oi_1
XFILLER_98_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _13089_/A _13074_/B vssd1 vssd1 vccd1 vccd1 _13075_/A sky130_fd_sc_hd__and2_1
X_10286_ _09980_/A _09980_/B _10285_/X vssd1 vssd1 vccd1 vccd1 _10311_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_output157_A _14312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12025_ _13790_/Q _12020_/X _12021_/X _13830_/Q vssd1 vssd1 vccd1 vccd1 _12026_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09491__A _09491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13976_ _14107_/CLK _13976_/D _12402_/Y vssd1 vssd1 vccd1 vccd1 _13976_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12927_ _14158_/Q _12915_/X _12926_/X _12920_/X vssd1 vssd1 vccd1 vccd1 _14158_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14259__D _14259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12858_ _13042_/B _12900_/B vssd1 vssd1 vccd1 vccd1 _12898_/B sky130_fd_sc_hd__or2_2
XFILLER_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _11809_/A vssd1 vssd1 vccd1 vccd1 _11845_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _14112_/Q _12782_/X _12787_/X _12788_/X _12207_/X vssd1 vssd1 vccd1 vccd1
+ _14112_/D sky130_fd_sc_hd__o221a_1
XANTENNA__12357__A _12360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14459_ _14467_/CLK _14459_/D vssd1 vssd1 vccd1 vccd1 _14459_/Q sky130_fd_sc_hd__dfxtp_1
X_07000_ _14453_/Q _14277_/Q vssd1 vssd1 vccd1 vccd1 _07000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_21_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__08570__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07233__A1 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08951_ _08935_/Y _08942_/Y _08944_/X _08950_/Y vssd1 vssd1 vccd1 vccd1 _08951_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07902_ _07901_/A _07840_/A _07840_/B _07874_/S vssd1 vssd1 vccd1 vccd1 _07902_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_97_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08882_ _08849_/A _08849_/B _08849_/C vssd1 vssd1 vccd1 vccd1 _08883_/C sky130_fd_sc_hd__a21oi_1
XFILLER_111_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07833_ _14025_/Q _13971_/Q vssd1 vssd1 vccd1 vccd1 _07834_/B sky130_fd_sc_hd__or2_1
XFILLER_99_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07764_ _07763_/Y _14149_/Q _07764_/S vssd1 vssd1 vccd1 vccd1 _07764_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09503_ _09471_/A _09471_/Y _09501_/X _09502_/Y vssd1 vssd1 vccd1 vccd1 _09518_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07695_ _14141_/Q _07665_/Y _07668_/X _07694_/X vssd1 vssd1 vccd1 vccd1 _07695_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09434_ _09434_/A _09434_/B vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__nand2_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _09425_/A _09873_/A _09364_/A _09364_/C vssd1 vssd1 vccd1 vccd1 _09367_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10486__S _10486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08316_ _08316_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _08364_/A sky130_fd_sc_hd__xnor2_2
XFILLER_20_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09296_ _09378_/A _09378_/B _09817_/B _09296_/D vssd1 vssd1 vccd1 vccd1 _09377_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__07472__A1 _14080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ _09769_/A _08247_/B vssd1 vssd1 vccd1 vccd1 _08257_/C sky130_fd_sc_hd__nand2_1
XFILLER_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09576__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08480__A _13861_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _08944_/C _10302_/A vssd1 vssd1 vccd1 vccd1 _09402_/A sky130_fd_sc_hd__nand2_4
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07224__A1 _07222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ _07126_/X _14293_/Q _07129_/S vssd1 vssd1 vccd1 vccd1 _07130_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10515__A _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10140_ _10141_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10166_/B sky130_fd_sc_hd__xnor2_1
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput170 _14295_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[3] sky130_fd_sc_hd__buf_2
X_10071_ _10098_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10071_/X sky130_fd_sc_hd__or2_1
XFILLER_47_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07824__A _14031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13830_ _14335_/CLK _13830_/D vssd1 vssd1 vccd1 vccd1 _13830_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12808__B1 _12807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ _14354_/CLK _13761_/D _11952_/Y vssd1 vssd1 vccd1 vccd1 _13761_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10973_ _10918_/A _10924_/X _10972_/X vssd1 vssd1 vccd1 vccd1 _11021_/A sky130_fd_sc_hd__o21ai_1
XFILLER_44_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ _12715_/A vssd1 vssd1 vccd1 vccd1 _12712_/Y sky130_fd_sc_hd__inv_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _13695_/A _13692_/B vssd1 vssd1 vccd1 vccd1 _13693_/A sky130_fd_sc_hd__and2_1
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12643_ _12656_/A _12643_/B vssd1 vssd1 vccd1 vccd1 _12644_/A sky130_fd_sc_hd__and2_1
XFILLER_54_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12177__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12574_ _12574_/A vssd1 vssd1 vccd1 vccd1 _14025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14313_ _14453_/CLK _14313_/D _13182_/Y vssd1 vssd1 vccd1 vccd1 _14313_/Q sky130_fd_sc_hd__dfrtp_4
X_11525_ _11525_/A _11525_/B vssd1 vssd1 vccd1 vccd1 _11525_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14244_ _14244_/CLK _14244_/D vssd1 vssd1 vccd1 vccd1 _14244_/Q sky130_fd_sc_hd__dfxtp_1
X_11456_ _11465_/B _11447_/Y _11451_/A vssd1 vssd1 vccd1 vccd1 _11456_/X sky130_fd_sc_hd__o21a_1
XFILLER_109_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10407_ _10407_/A vssd1 vssd1 vccd1 vccd1 _10493_/A sky130_fd_sc_hd__clkbuf_2
X_14175_ _14179_/CLK _14175_/D _12960_/Y vssd1 vssd1 vccd1 vccd1 _14175_/Q sky130_fd_sc_hd__dfrtp_1
X_11387_ _13885_/Q _11379_/X _11383_/X _11386_/X vssd1 vssd1 vccd1 vccd1 _13885_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13126_ _13128_/A vssd1 vssd1 vccd1 vccd1 _13126_/Y sky130_fd_sc_hd__inv_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ _10338_/A _10338_/B vssd1 vssd1 vccd1 vccd1 _10338_/Y sky130_fd_sc_hd__nor2_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ hold18/A _13051_/X _13032_/X vssd1 vssd1 vccd1 vccd1 _13057_/X sky130_fd_sc_hd__a21o_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10269_ _10269_/A _10269_/B vssd1 vssd1 vccd1 vccd1 _10297_/B sky130_fd_sc_hd__nand2_1
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12008_ _12008_/A _12008_/B vssd1 vssd1 vccd1 vccd1 _12009_/A sky130_fd_sc_hd__and2_1
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13959_ _13963_/CLK _13959_/D _12381_/Y vssd1 vssd1 vccd1 vccd1 _13959_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07480_ _14078_/Q _07459_/X _07460_/X _13878_/Q _07471_/X vssd1 vssd1 vccd1 vccd1
+ _07480_/X sky130_fd_sc_hd__a221o_1
XFILLER_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10825__A2 _10705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13224__B1 _13223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12087__A input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08284__B _09001_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ _09087_/B _09087_/C _09087_/A vssd1 vssd1 vccd1 vccd1 _09151_/C sky130_fd_sc_hd__a21bo_1
XFILLER_33_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08101_ _14013_/Q vssd1 vssd1 vccd1 vccd1 _09348_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09081_ _09081_/A _09081_/B _09081_/C vssd1 vssd1 vccd1 vccd1 _09083_/A sky130_fd_sc_hd__and3_1
XFILLER_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08032_ _09443_/A _09543_/B _08097_/B vssd1 vssd1 vccd1 vccd1 _08039_/A sky130_fd_sc_hd__and3_1
Xinput50 io_wbs_adr[25] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_1
Xinput61 io_wbs_adr[6] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_2
Xinput72 io_wbs_datwr[15] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput83 io_wbs_datwr[25] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_2
Xinput94 io_wbs_datwr[6] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__clkbuf_4
XFILLER_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ _10290_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__xor2_1
XFILLER_103_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08934_ _08934_/A _08934_/B vssd1 vssd1 vccd1 vccd1 _08935_/B sky130_fd_sc_hd__and2_1
XANTENNA__13646__A _13680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07644__A _14068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08865_ _08980_/A _08899_/A vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07816_ _14037_/Q _13983_/Q vssd1 vssd1 vccd1 vccd1 _07868_/A sky130_fd_sc_hd__or2_1
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08796_ _08796_/A _08796_/B _09806_/A _09200_/B vssd1 vssd1 vccd1 vccd1 _08797_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_26_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07747_ _07747_/A vssd1 vssd1 vccd1 vccd1 _14066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10277__A0 _10302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09131__A1 _09241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__B2 _09241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07678_ _07628_/Y _07678_/B vssd1 vssd1 vccd1 vccd1 _07679_/B sky130_fd_sc_hd__and2b_1
XFILLER_25_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09417_ _09342_/Y _09343_/X _09340_/X _09341_/X vssd1 vssd1 vccd1 vccd1 _09417_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08890__B1 _09943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09348_ _09457_/A _09348_/B _09457_/D _13872_/Q vssd1 vssd1 vccd1 vccd1 _09351_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_32_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07445__A1 _14085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ _09362_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _09281_/B sky130_fd_sc_hd__and2_1
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _11087_/B _10845_/X _11309_/X _10826_/X vssd1 vssd1 vccd1 vccd1 _13910_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07819__A _14034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12290_ _12291_/A vssd1 vssd1 vccd1 vccd1 _12290_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11241_ _11241_/A _11241_/B vssd1 vssd1 vccd1 vccd1 _11279_/B sky130_fd_sc_hd__xnor2_2
XFILLER_4_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ _11140_/B _11169_/X _11170_/X _11171_/X _10953_/A _10916_/A vssd1 vssd1 vccd1
+ vccd1 _11172_/X sky130_fd_sc_hd__mux4_2
XFILLER_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10123_ _10123_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _10123_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ _10054_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10055_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input33_A io_wbs_adr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09472__C _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11076__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A1 _09074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13813_ _14335_/CLK _13813_/D vssd1 vssd1 vccd1 vccd1 _13813_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13454__A0 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13744_ input90/X _14467_/Q _13744_/S vssd1 vssd1 vccd1 vccd1 _13745_/B sky130_fd_sc_hd__mux2_1
XFILLER_56_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10956_ _10953_/X _10955_/X _10940_/X _10744_/A vssd1 vssd1 vccd1 vccd1 _10963_/C
+ sky130_fd_sc_hd__a22oi_4
XFILLER_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08385__A _08385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13675_ _13678_/A _13675_/B vssd1 vssd1 vccd1 vccd1 _13676_/A sky130_fd_sc_hd__and2_1
X_10887_ _13932_/Q _10886_/X _10897_/S vssd1 vssd1 vccd1 vccd1 _10888_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12626_ _12695_/S vssd1 vssd1 vccd1 vccd1 _12642_/S sky130_fd_sc_hd__clkbuf_2
X_12557_ _12557_/A vssd1 vssd1 vccd1 vccd1 _14020_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11508_ _11058_/A _11489_/X _11499_/X _11279_/A _11490_/X vssd1 vssd1 vccd1 vccd1
+ _11508_/X sky130_fd_sc_hd__o221a_1
XFILLER_117_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12488_ _14035_/Q _12485_/X _12487_/X _12473_/X vssd1 vssd1 vccd1 vccd1 _12488_/X
+ sky130_fd_sc_hd__a211o_1
X_14227_ _14244_/CLK _14227_/D _13025_/Y vssd1 vssd1 vccd1 vccd1 _14227_/Q sky130_fd_sc_hd__dfrtp_4
X_11439_ _11297_/A _11076_/A _11446_/S vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__mux2_1
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14158_ _14158_/CLK _14158_/D vssd1 vssd1 vccd1 vccd1 _14158_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13109_ _13115_/A vssd1 vssd1 vccd1 vccd1 _13109_/Y sky130_fd_sc_hd__inv_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__B _09663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06980_ _14280_/Q _06968_/X _06979_/X _14376_/Q vssd1 vssd1 vccd1 vccd1 _06980_/X
+ sky130_fd_sc_hd__o211a_1
X_14089_ _14104_/CLK _14089_/D _12737_/Y vssd1 vssd1 vccd1 vccd1 _14089_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12370__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07464__A _07464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12496__A1 _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12496__B2 _14054_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__B _10621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08650_ _08435_/A _08836_/B _08599_/B _08595_/X vssd1 vssd1 vccd1 vccd1 _08656_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07601_ _07601_/A vssd1 vssd1 vccd1 vccd1 _14083_/D sky130_fd_sc_hd__clkbuf_1
X_08581_ _09493_/B _09361_/D _09092_/D _09443_/A vssd1 vssd1 vccd1 vccd1 _08582_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07532_ _14183_/Q _07530_/X _07531_/Y _07528_/A _07519_/X vssd1 vssd1 vccd1 vccd1
+ _14175_/D sky130_fd_sc_hd__o221a_1
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07463_ _07452_/X _07458_/X _07461_/X _07462_/X _14199_/Q vssd1 vssd1 vccd1 vccd1
+ _14199_/D sky130_fd_sc_hd__a32o_1
XFILLER_23_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09202_ _09202_/A _09202_/B _09202_/C vssd1 vssd1 vccd1 vccd1 _09205_/A sky130_fd_sc_hd__nand3_1
XFILLER_22_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07394_ _14211_/Q _07373_/X _07375_/X _07393_/X vssd1 vssd1 vccd1 vccd1 _14211_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09133_ _09133_/A _09133_/B vssd1 vssd1 vccd1 vccd1 _09135_/A sky130_fd_sc_hd__nor2_1
X_09064_ _09063_/A _09063_/B _09063_/C vssd1 vssd1 vccd1 vccd1 _09065_/C sky130_fd_sc_hd__a21o_1
X_08015_ _08128_/A _08126_/A _09834_/A _08289_/A vssd1 vssd1 vccd1 vccd1 _08078_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_89_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08927__B2 _08891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11595__S _11611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12280__A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _10465_/B _09966_/B _09966_/C vssd1 vssd1 vccd1 vccd1 _09967_/B sky130_fd_sc_hd__nand3_1
XFILLER_58_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08917_ _08683_/X _08941_/B _08895_/A _08892_/B vssd1 vssd1 vccd1 vccd1 _08919_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13684__A0 _12681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__A1 _08128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ _09894_/A _09897_/B vssd1 vssd1 vccd1 vccd1 _09897_/X sky130_fd_sc_hd__and2b_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08848_ _08848_/A _08848_/B vssd1 vssd1 vccd1 vccd1 _08849_/C sky130_fd_sc_hd__xnor2_1
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11064__A_N _11014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _08779_/A _08779_/B vssd1 vssd1 vccd1 vccd1 _08779_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10810_ _10853_/B _10810_/B vssd1 vssd1 vccd1 vccd1 _10858_/A sky130_fd_sc_hd__or2_1
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11790_/A _11790_/B vssd1 vssd1 vccd1 vccd1 _11791_/A sky130_fd_sc_hd__or2_4
XFILLER_41_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _10953_/A vssd1 vssd1 vccd1 vccd1 _11184_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_16_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13460_ input87/X _14385_/Q _13460_/S vssd1 vssd1 vccd1 vccd1 _13461_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10672_ _10944_/S vssd1 vssd1 vccd1 vccd1 _11171_/S sky130_fd_sc_hd__buf_2
X_12411_ _12415_/A vssd1 vssd1 vccd1 vccd1 _12411_/Y sky130_fd_sc_hd__inv_2
X_13391_ _12664_/X _14365_/Q _13391_/S vssd1 vssd1 vccd1 vccd1 _13392_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08652__B _09233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12342_ _12348_/A vssd1 vssd1 vccd1 vccd1 _12347_/A sky130_fd_sc_hd__buf_2
XFILLER_103_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12273_ _12273_/A vssd1 vssd1 vccd1 vccd1 _12273_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14012_ _14304_/CLK _14012_/D vssd1 vssd1 vccd1 vccd1 _14012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11224_ _11228_/B _11229_/A _11228_/A vssd1 vssd1 vccd1 vccd1 _11225_/B sky130_fd_sc_hd__a21oi_1
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11155_ _13916_/Q _13917_/Q _11155_/S vssd1 vssd1 vccd1 vccd1 _11155_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10106_ _10106_/A _10106_/B vssd1 vssd1 vccd1 vccd1 _10121_/B sky130_fd_sc_hd__xor2_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12478__A1 _14033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11086_ _11093_/A _11083_/A _11084_/X _11085_/Y vssd1 vssd1 vccd1 vccd1 _11090_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_23_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10037_ _10037_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _10354_/A sky130_fd_sc_hd__xnor2_4
XFILLER_49_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11988_ _11988_/A _13203_/B vssd1 vssd1 vccd1 vccd1 _12001_/B sky130_fd_sc_hd__nor2_1
XFILLER_91_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13727_ _13727_/A vssd1 vssd1 vccd1 vccd1 _14461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10939_ _10946_/B vssd1 vssd1 vccd1 vccd1 _10960_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13658_ _13661_/A _13658_/B vssd1 vssd1 vccd1 vccd1 _13659_/A sky130_fd_sc_hd__and2_1
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12609_ _12609_/A vssd1 vssd1 vccd1 vccd1 _14035_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07409__A1 _07399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13589_ input75/X _14422_/Q _13593_/S vssd1 vssd1 vccd1 vccd1 _13590_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12365__A _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11700__C _11906_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14183__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09674__A _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13196__A _13265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ _09826_/A vssd1 vssd1 vccd1 vccd1 _10151_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07593__A0 _14086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09751_ _09751_/A _09751_/B _09751_/C vssd1 vssd1 vccd1 vccd1 _09751_/Y sky130_fd_sc_hd__nor3_2
XFILLER_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06963_ _14282_/Q _06929_/X _06962_/X _14378_/Q vssd1 vssd1 vccd1 vccd1 _06963_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12469__A1 _08842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08702_ _08701_/A _08701_/C _08701_/B vssd1 vssd1 vccd1 vccd1 _08708_/B sky130_fd_sc_hd__a21o_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09334__A1 _09319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09682_ _09683_/B _09683_/C _09683_/A vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__a21oi_1
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06894_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06894_/X sky130_fd_sc_hd__buf_4
XFILLER_55_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08633_ _09001_/B _08449_/C _09011_/B _09001_/A vssd1 vssd1 vccd1 vccd1 _08634_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08564_ _08727_/A _08564_/B vssd1 vssd1 vccd1 vccd1 _08566_/A sky130_fd_sc_hd__xnor2_1
XFILLER_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07515_ hold34/X _14180_/Q _07517_/S vssd1 vssd1 vccd1 vccd1 _07516_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08495_ _13862_/Q vssd1 vssd1 vccd1 vccd1 _09865_/A sky130_fd_sc_hd__buf_2
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07446_ _07425_/X _07443_/X _07445_/X _07435_/X _14202_/Q vssd1 vssd1 vccd1 vccd1
+ _14202_/D sky130_fd_sc_hd__a32o_1
XANTENNA__08753__A _14009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07377_ _14097_/Q _07363_/X vssd1 vssd1 vccd1 vccd1 _07377_/X sky130_fd_sc_hd__or2b_1
XANTENNA__12275__A _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ _09032_/X _09040_/Y _09114_/Y _09115_/X vssd1 vssd1 vccd1 vccd1 _10632_/B
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__07369__A _14098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__A1 _13895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ _09048_/A _09048_/B _09048_/C vssd1 vssd1 vccd1 vccd1 _09049_/A sky130_fd_sc_hd__a21oi_4
XFILLER_11_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09584__A _09584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ _10206_/B _10016_/B _10208_/A vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__13657__A0 input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12960_ _12960_/A vssd1 vssd1 vccd1 vccd1 _12960_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11911_ _13759_/Q _11911_/B vssd1 vssd1 vccd1 vccd1 _11911_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07832__A _14025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12936_/A _12896_/B vssd1 vssd1 vccd1 vccd1 _12891_/X sky130_fd_sc_hd__or2_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _14339_/Q _11833_/X _11834_/X _13798_/Q _11841_/X vssd1 vssd1 vccd1 vccd1
+ _11842_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ input61/X vssd1 vssd1 vccd1 vccd1 _11774_/A sky130_fd_sc_hd__clkinv_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _13518_/A _13512_/B vssd1 vssd1 vccd1 vccd1 _13513_/A sky130_fd_sc_hd__and2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _13949_/Q vssd1 vssd1 vccd1 vccd1 _11158_/S sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13443_ input82/X _14380_/Q _13443_/S vssd1 vssd1 vccd1 vccd1 _13444_/B sky130_fd_sc_hd__mux2_1
X_10655_ _10655_/A _10664_/B vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__or2_2
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13374_ _12641_/X _14360_/Q _13374_/S vssd1 vssd1 vccd1 vccd1 _13375_/B sky130_fd_sc_hd__mux2_1
XFILLER_70_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10586_ _10586_/A vssd1 vssd1 vccd1 vccd1 _13960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12325_ _12329_/A vssd1 vssd1 vccd1 vccd1 _12325_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12913__A _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09013__B1 _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12256_ _12259_/A vssd1 vssd1 vccd1 vccd1 _12256_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11207_ _11207_/A _11207_/B vssd1 vssd1 vccd1 vccd1 _11208_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12187_ _12187_/A vssd1 vssd1 vccd1 vccd1 _13832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11138_ _10912_/A _11140_/B _11175_/S vssd1 vssd1 vccd1 vccd1 _11138_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11069_ _11111_/B _11115_/B _11111_/A vssd1 vssd1 vccd1 vccd1 _11112_/B sky130_fd_sc_hd__o21a_1
XFILLER_95_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11123__A1 _11119_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11123__B2 _11056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08827__B1 _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13943_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_07300_ _14225_/Q _07300_/B _14166_/Q vssd1 vssd1 vccd1 vccd1 _07313_/C sky130_fd_sc_hd__or3_1
XFILLER_20_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08280_ _08280_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _09749_/A sky130_fd_sc_hd__xor2_1
X_07231_ _07231_/A vssd1 vssd1 vccd1 vccd1 _14269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11711__B _11882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07162_ _14288_/Q _07161_/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07163_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07093_ _07089_/X _14298_/Q _07093_/S vssd1 vssd1 vccd1 vccd1 _07094_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13351__A2 _13236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09803_ _09803_/A _09803_/B vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__xor2_2
XFILLER_8_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07995_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08024_/C sky130_fd_sc_hd__nand2_1
XFILLER_68_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09734_ _08406_/A _08404_/Y _08402_/X _08403_/X vssd1 vssd1 vccd1 vccd1 _09735_/B
+ sky130_fd_sc_hd__o211a_1
X_06946_ _14460_/Q _14284_/Q vssd1 vssd1 vccd1 vccd1 _06946_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08748__A _08789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_io_wbs_clk clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14054_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09665_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _10576_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06877_ _06970_/A vssd1 vssd1 vccd1 vccd1 _06877_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08616_ _08617_/A _08616_/B _08616_/C vssd1 vssd1 vccd1 vccd1 _08738_/A sky130_fd_sc_hd__nand3_1
XFILLER_15_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _08547_/A _09152_/A _08824_/C _08547_/D vssd1 vssd1 vccd1 vccd1 _08584_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__12614__A1 _14037_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10625__B1 _10528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07097__A2 _07085_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _09378_/A vssd1 vssd1 vccd1 vccd1 _09493_/A sky130_fd_sc_hd__buf_4
XFILLER_11_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07429_ _07425_/X _07427_/X _07428_/X _07408_/X _14205_/Q vssd1 vssd1 vccd1 vccd1
+ _14205_/D sky130_fd_sc_hd__a32o_1
XFILLER_11_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _10440_/A _10425_/B vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__or2b_1
XFILLER_109_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10371_ _10572_/A _10583_/A vssd1 vssd1 vccd1 vccd1 _10376_/A sky130_fd_sc_hd__or2_1
XFILLER_108_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _13810_/Q _12095_/X _12109_/X _11931_/X vssd1 vssd1 vccd1 vccd1 _13810_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07827__A _14028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ _13090_/A vssd1 vssd1 vccd1 vccd1 _14248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12041_ _12044_/A _12041_/B vssd1 vssd1 vccd1 vccd1 _12042_/A sky130_fd_sc_hd__and2_1
XFILLER_2_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12550__A0 _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13992_ _14441_/CLK _13992_/D vssd1 vssd1 vccd1 vccd1 _13992_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08658__A _08980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12943_ hold37/A _12928_/A _12942_/X _12934_/X vssd1 vssd1 vccd1 vccd1 _14164_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12853__A1 _14132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12874_ _12917_/A _12883_/B vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__or2_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11825_ _14332_/Q _11808_/X _11823_/X _13791_/Q _11824_/X vssd1 vssd1 vccd1 vccd1
+ _11825_/X sky130_fd_sc_hd__a221o_2
XFILLER_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10616__B1 _07924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11756_ _11756_/A _11756_/B vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__nor2_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08824__C _08824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ _13942_/Q _10708_/B vssd1 vssd1 vccd1 vccd1 _10828_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11687_ _11682_/B _11661_/X _11686_/A vssd1 vssd1 vccd1 vccd1 _11687_/Y sky130_fd_sc_hd__a21oi_1
X_13426_ _13426_/A _13426_/B vssd1 vssd1 vccd1 vccd1 _13427_/A sky130_fd_sc_hd__and2_1
XANTENNA__09001__B _09001_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10638_ _10638_/A _10638_/B vssd1 vssd1 vccd1 vccd1 _10639_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13357_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13375_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10569_ _10598_/A _10598_/B vssd1 vssd1 vccd1 vccd1 _10587_/A sky130_fd_sc_hd__and2_1
X_12308_ _12310_/A vssd1 vssd1 vccd1 vccd1 _12308_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07737__A _14157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13288_ _14338_/Q _13265_/X _13287_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _14338_/D
+ sky130_fd_sc_hd__o211a_1
X_12239_ _12239_/A vssd1 vssd1 vccd1 vccd1 _12239_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07548__A0 _14106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12541__A0 _12924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11895__A2 _11872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07780_ _07780_/A vssd1 vssd1 vccd1 vccd1 _13988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 dout1[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__11706__B _11882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09450_ _09450_/A _09450_/B vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__14371__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08401_ _09729_/A _08399_/Y _08337_/A _08400_/Y vssd1 vssd1 vccd1 vccd1 _08406_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09381_ _14015_/Q _09796_/A vssd1 vssd1 vccd1 vccd1 _09382_/C sky130_fd_sc_hd__nand2_1
XFILLER_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08332_ _08391_/A _08330_/Y _08122_/X _08331_/Y vssd1 vssd1 vccd1 vccd1 _08336_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08263_ _08263_/A _08263_/B vssd1 vssd1 vccd1 vccd1 _08264_/B sky130_fd_sc_hd__nand2_1
X_07214_ _07214_/A vssd1 vssd1 vccd1 vccd1 _14274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08194_ _08194_/A _08194_/B _08194_/C vssd1 vssd1 vccd1 vccd1 _08194_/X sky130_fd_sc_hd__or3_2
XFILLER_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07145_ _13838_/Q vssd1 vssd1 vccd1 vccd1 _07146_/B sky130_fd_sc_hd__inv_2
X_07076_ _07073_/X _14300_/Q _07076_/S vssd1 vssd1 vccd1 vccd1 _07077_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07978_ _08547_/A _09241_/D _09445_/B _08573_/A vssd1 vssd1 vccd1 vccd1 _07985_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__07382__A _14096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09717_ _09710_/X _09720_/A _09706_/Y _09707_/X vssd1 vssd1 vccd1 vccd1 _09717_/X
+ sky130_fd_sc_hd__a211o_1
X_06929_ _06968_/A vssd1 vssd1 vccd1 vccd1 _06929_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08197__B _08198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _09638_/B _09640_/X _09647_/X _09651_/A vssd1 vssd1 vccd1 vccd1 _09650_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_71_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09576_/X _09577_/X _09575_/X _09578_/Y vssd1 vssd1 vccd1 vccd1 _09622_/A
+ sky130_fd_sc_hd__a211oi_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__A _13010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11610_/Y sky130_fd_sc_hd__xnor2_4
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12590_ _12919_/A _14030_/Q _12600_/S vssd1 vssd1 vccd1 vccd1 _12591_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11541_ _14052_/Q _13964_/Q vssd1 vssd1 vccd1 vccd1 _11541_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14260_ _14281_/CLK _14260_/D _13117_/Y vssd1 vssd1 vccd1 vccd1 _14260_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11472_ _11474_/A vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__clkbuf_2
X_13211_ _14356_/Q _13208_/X _13210_/X vssd1 vssd1 vccd1 vccd1 _13211_/X sky130_fd_sc_hd__a21o_1
X_10423_ _10423_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _10423_/X sky130_fd_sc_hd__or2b_1
X_14191_ _14244_/CLK _14191_/D _12981_/Y vssd1 vssd1 vccd1 vccd1 _14191_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13142_ _13146_/A vssd1 vssd1 vccd1 vccd1 _13142_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10354_ _10354_/A _10354_/B vssd1 vssd1 vccd1 vccd1 _10354_/X sky130_fd_sc_hd__and2_1
XANTENNA_input63_A io_wbs_adr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__A _11079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ _12515_/X _14244_/Q _13076_/S vssd1 vssd1 vccd1 vccd1 _13074_/B sky130_fd_sc_hd__mux2_1
X_10285_ _10159_/A _10285_/B vssd1 vssd1 vccd1 vccd1 _10285_/X sky130_fd_sc_hd__and2b_1
X_12024_ _12024_/A vssd1 vssd1 vccd1 vccd1 _13789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13294__A _13315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09491__B _09792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14394__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10711__A _11244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12826__A1 _12209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13975_ _13982_/CLK _13975_/D _12401_/Y vssd1 vssd1 vccd1 vccd1 _13975_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ _12926_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _12926_/X sky130_fd_sc_hd__or2_1
XFILLER_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10301__A2 _10279_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _12885_/A vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _11855_/A vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__clkbuf_4
X_12788_ _14137_/Q _12776_/X _12760_/X vssd1 vssd1 vccd1 vccd1 _12788_/X sky130_fd_sc_hd__a21o_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13251__B2 _14395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09012__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11739_ _13764_/Q _11740_/B vssd1 vssd1 vccd1 vccd1 _11739_/X sky130_fd_sc_hd__and2_1
XFILLER_31_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14458_ _14467_/CLK _14458_/D vssd1 vssd1 vccd1 vccd1 _14458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13409_ _13409_/A _13409_/B vssd1 vssd1 vccd1 vccd1 _13410_/A sky130_fd_sc_hd__and2_1
X_14389_ _14450_/CLK _14389_/D vssd1 vssd1 vccd1 vccd1 _14389_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12373__A _12379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08950_ _08950_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08950_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_29_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07901_ _07901_/A _07901_/B vssd1 vssd1 vccd1 vccd1 _07901_/Y sky130_fd_sc_hd__nor2_1
X_08881_ _08904_/A _08904_/B vssd1 vssd1 vccd1 vccd1 _08883_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11717__A _13830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07832_ _14025_/Q _13971_/Q vssd1 vssd1 vccd1 vccd1 _07834_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08298__A _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10621__A _10621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07763_ _07763_/A vssd1 vssd1 vccd1 vccd1 _07763_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09502_ _09540_/A _09540_/C _09540_/B vssd1 vssd1 vccd1 vccd1 _09502_/Y sky130_fd_sc_hd__a21oi_1
X_07694_ _14140_/Q _07740_/A _07744_/A _14139_/Q _07693_/X vssd1 vssd1 vccd1 vccd1
+ _07694_/X sky130_fd_sc_hd__a221o_1
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07930__A _10547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ _09431_/X _09433_/B vssd1 vssd1 vccd1 vccd1 _09435_/A sky130_fd_sc_hd__and2b_1
XFILLER_80_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09364_ _09364_/A _09364_/B _09364_/C vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__nand3_1
XFILLER_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08315_ _08315_/A _08315_/B vssd1 vssd1 vccd1 vccd1 _08316_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09295_ _09295_/A _09223_/A vssd1 vssd1 vccd1 vccd1 _09305_/A sky130_fd_sc_hd__or2b_1
X_08246_ _08246_/A _08214_/A vssd1 vssd1 vccd1 vccd1 _08257_/B sky130_fd_sc_hd__or2b_1
XANTENNA__09857__A _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _09786_/A vssd1 vssd1 vccd1 vccd1 _10302_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ _06973_/A _07127_/X _14385_/Q vssd1 vssd1 vccd1 vccd1 _07129_/S sky130_fd_sc_hd__o21a_1
XANTENNA__07377__A _14097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07059_ _14414_/Q _07059_/B _14446_/Q vssd1 vssd1 vccd1 vccd1 _07059_/X sky130_fd_sc_hd__and3b_1
XFILLER_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput160 _14315_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[23] sky130_fd_sc_hd__buf_2
XANTENNA__06983__A1 _14312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput171 _14296_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[4] sky130_fd_sc_hd__buf_2
XFILLER_0_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__xnor2_1
XFILLER_43_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08185__B1 _08091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08001__A _08291_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13760_ _14354_/CLK _13760_/D _11951_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10972_ _11181_/A _10957_/X _10959_/X _10975_/A vssd1 vssd1 vccd1 vccd1 _10972_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12711_ _12715_/A vssd1 vssd1 vccd1 vccd1 _12711_/Y sky130_fd_sc_hd__inv_2
X_13691_ _12688_/X _14451_/Q _13704_/S vssd1 vssd1 vccd1 vccd1 _13692_/B sky130_fd_sc_hd__mux2_1
XFILLER_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12458__A _12817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12642_ _12641_/X _14044_/Q _12642_/S vssd1 vssd1 vccd1 vccd1 _12643_/B sky130_fd_sc_hd__mux2_1
XFILLER_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13233__A1 _14359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12573_ _12576_/A _12573_/B vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__and2_1
XFILLER_12_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11524_ _08941_/B _11510_/X _11522_/X _11523_/X vssd1 vssd1 vccd1 vccd1 _13862_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14312_ _14453_/CLK _14312_/D _13181_/Y vssd1 vssd1 vccd1 vccd1 _14312_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_12_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13289__A _13332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14243_ _14256_/CLK _14243_/D vssd1 vssd1 vccd1 vccd1 _14243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_109_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11455_ _11510_/A vssd1 vssd1 vccd1 vccd1 _11455_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__06903__B _07085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _10478_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _10459_/B sky130_fd_sc_hd__xnor2_1
X_14174_ _14179_/CLK _14174_/D _12959_/Y vssd1 vssd1 vccd1 vccd1 _14174_/Q sky130_fd_sc_hd__dfrtp_1
X_11386_ hold9/X _11390_/B vssd1 vssd1 vccd1 vccd1 _11386_/X sky130_fd_sc_hd__or2_1
XFILLER_113_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13125_ _13128_/A vssd1 vssd1 vccd1 vccd1 _13125_/Y sky130_fd_sc_hd__inv_2
X_10337_ _10337_/A _10350_/B vssd1 vssd1 vccd1 vccd1 _10347_/A sky130_fd_sc_hd__xnor2_1
XFILLER_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _14238_/Q _13041_/A _13055_/X _13053_/X vssd1 vssd1 vccd1 vccd1 _14238_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10268_ _10268_/A _10268_/B vssd1 vssd1 vccd1 vccd1 _10297_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ _13785_/Q _12000_/X _12003_/X _13825_/Q vssd1 vssd1 vccd1 vccd1 _12008_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11537__A _14056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10199_ _10199_/A _10199_/B vssd1 vssd1 vccd1 vccd1 _10200_/B sky130_fd_sc_hd__and2_1
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08479__A1 _09493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13958_ _13963_/CLK _13958_/D _12380_/Y vssd1 vssd1 vccd1 vccd1 _13958_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12909_ _12909_/A _12913_/B vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__or2_1
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13889_ _13892_/CLK _13889_/D _12295_/Y vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfrtp_1
XFILLER_59_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12368__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12087__B input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08100_ _08750_/A vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__buf_2
X_09080_ _09079_/A _09079_/C _09079_/B vssd1 vssd1 vccd1 vccd1 _09081_/C sky130_fd_sc_hd__a21o_1
X_08031_ _13875_/Q vssd1 vssd1 vccd1 vccd1 _08097_/B sky130_fd_sc_hd__clkbuf_2
Xinput40 io_wbs_adr[16] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__13199__A _13306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput51 io_wbs_adr[26] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_1
Xinput62 io_wbs_adr[7] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_4
Xinput73 io_wbs_datwr[16] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_4
Xinput84 io_wbs_datwr[26] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_2
Xinput95 io_wbs_datwr[7] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__buf_4
XFILLER_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09982_ _09880_/A _09880_/B _09981_/X vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__o21ai_1
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08933_ _08896_/A _10156_/A _08948_/D vssd1 vssd1 vccd1 vccd1 _08934_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07925__A _14023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12499__C1 _12498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08864_ _08864_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__nor2_1
XFILLER_29_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07815_ _14037_/Q _13983_/Q vssd1 vssd1 vccd1 vccd1 _07868_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08795_ _08828_/B _09807_/A _09092_/C _08828_/A vssd1 vssd1 vccd1 vccd1 _08797_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_42_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07746_ _14066_/Q _07745_/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__mux2_1
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10277__A1 _10486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ _14135_/Q vssd1 vssd1 vccd1 vccd1 _07687_/A sky130_fd_sc_hd__inv_2
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12278__A _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _09340_/X _09341_/X _09342_/Y _09343_/X vssd1 vssd1 vccd1 vccd1 _09416_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08890__B2 _08891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ _09305_/A _09303_/X _09304_/A vssd1 vssd1 vccd1 vccd1 _09626_/B sky130_fd_sc_hd__a21o_1
XFILLER_32_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ _09361_/A _09361_/B _09807_/B _09866_/A vssd1 vssd1 vccd1 vccd1 _09281_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_32_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08491__A _09297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ _08265_/B _08227_/Y _08170_/A _08170_/Y vssd1 vssd1 vccd1 vccd1 _08234_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_107_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11240_ _11240_/A _11240_/B vssd1 vssd1 vccd1 vccd1 _11241_/B sky130_fd_sc_hd__nor2_1
XFILLER_5_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11171_ _13921_/Q _13922_/Q _11171_/S vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06956__A1 _14283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10122_ _10122_/A vssd1 vssd1 vccd1 vccd1 _10122_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11357__A _14057_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _10053_/A _10053_/B vssd1 vssd1 vccd1 vccd1 _10064_/A sky130_fd_sc_hd__xnor2_1
XFILLER_48_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input26_A dout1[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13812_ _14400_/CLK _13812_/D vssd1 vssd1 vccd1 vccd1 _13812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10955_ _13895_/Q _10674_/A _10771_/Y _10954_/X vssd1 vssd1 vccd1 vccd1 _10955_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13743_ _13743_/A vssd1 vssd1 vccd1 vccd1 _14466_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07133__A1 _14279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11092__A _11092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13674_ _12668_/X _14446_/Q _13687_/S vssd1 vssd1 vccd1 vccd1 _13675_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10886_ _10836_/S _10879_/C _10884_/Y _10885_/X vssd1 vssd1 vccd1 vccd1 _10886_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06892__B1 _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12625_ _12669_/A vssd1 vssd1 vccd1 vccd1 _12695_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_19_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08633__A1 _09001_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ _12576_/A _12556_/B vssd1 vssd1 vccd1 vccd1 _12557_/A sky130_fd_sc_hd__and2_1
XFILLER_12_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11507_ _11502_/A _11506_/X _10686_/X vssd1 vssd1 vccd1 vccd1 _11507_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12487_ _08128_/B _12486_/X _12476_/X _14051_/Q vssd1 vssd1 vccd1 vccd1 _12487_/X
+ sky130_fd_sc_hd__a22o_1
X_11438_ _11482_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11478_/A sky130_fd_sc_hd__nand2_1
X_14226_ _14244_/CLK _14226_/D _13024_/Y vssd1 vssd1 vccd1 vccd1 _14226_/Q sky130_fd_sc_hd__dfrtp_1
X_14157_ _14158_/CLK _14157_/D vssd1 vssd1 vccd1 vccd1 _14157_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10870__S _10875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ _13892_/Q _11363_/X _11367_/X _11396_/A vssd1 vssd1 vccd1 vccd1 _13892_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _13115_/A vssd1 vssd1 vccd1 vccd1 _13108_/Y sky130_fd_sc_hd__inv_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _14104_/CLK _14088_/D _12736_/Y vssd1 vssd1 vccd1 vccd1 _14088_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_112_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13039_ _13254_/A vssd1 vssd1 vccd1 vccd1 _13039_/X sky130_fd_sc_hd__clkbuf_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10171__A _10171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07600_ _14083_/Q input30/X _07604_/S vssd1 vssd1 vccd1 vccd1 _07601_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08580_ _08580_/A _08580_/B _09092_/C _09870_/A vssd1 vssd1 vccd1 vccd1 _08637_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_82_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07531_ _14175_/Q _07534_/A vssd1 vssd1 vccd1 vccd1 _07531_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12098__A _12147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_33_io_wbs_clk_A clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07462_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07462_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09201_ _09424_/B _09866_/A _09199_/D _09424_/A vssd1 vssd1 vccd1 vccd1 _09202_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07393_ _07376_/X _07390_/X _07392_/X _07379_/X vssd1 vssd1 vccd1 vccd1 _07393_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11730__A _13827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09132_ _09132_/A _09132_/B _09792_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09133_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__08624__A1 _08623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08624__B2 _08623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09200__A _14021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ _09063_/A _09063_/B _09063_/C vssd1 vssd1 vccd1 vccd1 _09065_/B sky130_fd_sc_hd__nand3_2
XFILLER_8_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08014_ _09545_/D vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__buf_4
XFILLER_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08927__A2 _09943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12561__A input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14305__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ _09966_/B _09966_/C _10465_/B vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__a21o_1
X_08916_ _08916_/A _08916_/B vssd1 vssd1 vccd1 vccd1 _08924_/A sky130_fd_sc_hd__and2_1
XANTENNA__10081__A _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09896_ _09896_/A _09896_/B vssd1 vssd1 vccd1 vccd1 _09902_/B sky130_fd_sc_hd__and2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09870__A _09870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _08850_/A _08850_/C _08879_/A vssd1 vssd1 vccd1 vccd1 _08849_/B sky130_fd_sc_hd__a21o_1
XFILLER_18_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08778_ _08776_/A _08777_/A _08776_/B _08781_/A _08781_/B vssd1 vssd1 vccd1 vccd1
+ _08778_/X sky130_fd_sc_hd__o32a_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08486__A _13860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07390__A _14094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _07727_/Y _14159_/Q _07757_/S vssd1 vssd1 vccd1 vccd1 _07729_/X sky130_fd_sc_hd__mux2_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07115__A1 _14295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10740_ _10923_/S vssd1 vssd1 vccd1 vccd1 _10953_/A sky130_fd_sc_hd__buf_2
XFILLER_53_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _13947_/Q vssd1 vssd1 vccd1 vccd1 _10944_/S sky130_fd_sc_hd__clkbuf_2
X_12410_ _12410_/A vssd1 vssd1 vccd1 vccd1 _12415_/A sky130_fd_sc_hd__buf_2
XFILLER_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13390_ _13390_/A vssd1 vssd1 vccd1 vccd1 _14364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08652__C _09074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ _12341_/A vssd1 vssd1 vccd1 vccd1 _12341_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12272_ _12273_/A vssd1 vssd1 vccd1 vccd1 _12272_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14011_ _14304_/CLK _14011_/D vssd1 vssd1 vccd1 vccd1 _14011_/Q sky130_fd_sc_hd__dfxtp_2
X_11223_ _13904_/Q vssd1 vssd1 vccd1 vccd1 _11291_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ _11032_/A _13915_/Q _11155_/S vssd1 vssd1 vccd1 vccd1 _11154_/X sky130_fd_sc_hd__mux2_1
X_10105_ _10106_/A _10106_/B vssd1 vssd1 vccd1 vccd1 _10120_/A sky130_fd_sc_hd__or2_1
XANTENNA__11087__A _11142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11085_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10036_ _10045_/A _10036_/B vssd1 vssd1 vccd1 vccd1 _10037_/B sky130_fd_sc_hd__xor2_2
XFILLER_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13822__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11987_ input33/X input44/X _12429_/A vssd1 vssd1 vccd1 vccd1 _13203_/B sky130_fd_sc_hd__or3_2
Xclkbuf_leaf_12_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14041_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13726_ _13729_/A _13726_/B vssd1 vssd1 vccd1 vccd1 _13727_/A sky130_fd_sc_hd__and2_1
X_10938_ _13903_/Q _13904_/Q _13905_/Q _13906_/Q _10944_/S _10954_/A vssd1 vssd1 vccd1
+ vccd1 _10938_/X sky130_fd_sc_hd__mux4_1
XFILLER_31_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13657_ input93/X _14441_/Q _13670_/S vssd1 vssd1 vccd1 vccd1 _13658_/B sky130_fd_sc_hd__mux2_1
X_10869_ _10869_/A _10869_/B vssd1 vssd1 vccd1 vccd1 _10869_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12608_ _12615_/A _12608_/B vssd1 vssd1 vccd1 vccd1 _12609_/A sky130_fd_sc_hd__and2_1
XFILLER_118_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13588_ _13588_/A vssd1 vssd1 vccd1 vccd1 _14421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12539_ _12539_/A vssd1 vssd1 vccd1 vccd1 _14015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14209_ _14217_/CLK _14209_/D _13002_/Y vssd1 vssd1 vccd1 vccd1 _14209_/Q sky130_fd_sc_hd__dfrtp_1
X_14471__183 vssd1 vssd1 vccd1 vccd1 _14471__183/HI io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_99_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10613__B _10613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08790__B1 _13859_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06962_ _14426_/Q _06961_/Y _06931_/X vssd1 vssd1 vccd1 vccd1 _06962_/X sky130_fd_sc_hd__a21o_1
X_09750_ _09781_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09750_/Y sky130_fd_sc_hd__nand2_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08701_ _08701_/A _08701_/B _08701_/C vssd1 vssd1 vccd1 vccd1 _08709_/A sky130_fd_sc_hd__nand3_1
XFILLER_100_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_51_io_wbs_clk clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14400_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09690__A _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ _09681_/A _09598_/B vssd1 vssd1 vccd1 vccd1 _09683_/C sky130_fd_sc_hd__or2b_1
X_06893_ _07090_/A vssd1 vssd1 vccd1 vccd1 _06973_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08632_ _08632_/A _09001_/B _08918_/B _08899_/A vssd1 vssd1 vccd1 vccd1 _08998_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08563_ _08727_/A _08564_/B vssd1 vssd1 vccd1 vccd1 _08567_/A sky130_fd_sc_hd__or2b_1
XFILLER_81_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07514_ _07514_/A vssd1 vssd1 vccd1 vccd1 _14181_/D sky130_fd_sc_hd__clkbuf_1
X_08494_ _08560_/A _08490_/Y _09000_/A _08494_/D vssd1 vssd1 vccd1 vccd1 _08560_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07445_ _14085_/Q _07432_/X _07433_/X _13885_/Q _07444_/X vssd1 vssd1 vccd1 vccd1
+ _07445_/X sky130_fd_sc_hd__a221o_1
XFILLER_11_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12556__A _12576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08753__B _09000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07376_ _07376_/A vssd1 vssd1 vccd1 vccd1 _07376_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09115_ _09114_/B _09114_/C _09114_/A vssd1 vssd1 vccd1 vccd1 _09115_/X sky130_fd_sc_hd__o21a_1
XFILLER_109_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09046_ _08979_/A _08981_/B _08979_/B vssd1 vssd1 vccd1 vccd1 _09048_/C sky130_fd_sc_hd__o21ba_2
XFILLER_85_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13354__B1 _13201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09948_ _09948_/A _09946_/B vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__or2b_1
XFILLER_86_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09879_ _10174_/A _10173_/A vssd1 vssd1 vccd1 vccd1 _09880_/B sky130_fd_sc_hd__xor2_1
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11910_ _13818_/Q _11872_/A _11908_/X _11909_/Y hold38/X vssd1 vssd1 vccd1 vccd1
+ _13758_/D sky130_fd_sc_hd__o221a_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ _14144_/Q _12885_/X _12889_/X _12879_/X vssd1 vssd1 vccd1 vccd1 _14144_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _14004_/Q _11797_/A _11830_/X _14123_/Q vssd1 vssd1 vccd1 vccd1 _11841_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _12951_/A vssd1 vssd1 vccd1 vccd1 _12193_/A sky130_fd_sc_hd__buf_2
XFILLER_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10643__A1 _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13511_ _12610_/X _14400_/Q _13511_/S vssd1 vssd1 vccd1 vccd1 _13512_/B sky130_fd_sc_hd__mux2_1
XFILLER_41_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _11207_/A _10746_/A _10748_/A vssd1 vssd1 vccd1 vccd1 _10818_/B sky130_fd_sc_hd__mux2_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input93_A io_wbs_datwr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13442_ _13442_/A vssd1 vssd1 vccd1 vccd1 _14379_/D sky130_fd_sc_hd__clkbuf_1
X_10654_ _10836_/S vssd1 vssd1 vccd1 vccd1 _10826_/A sky130_fd_sc_hd__buf_2
XANTENNA__13593__A0 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13373_ _13373_/A vssd1 vssd1 vccd1 vccd1 _14359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10585_ _13960_/Q _10584_/X _10585_/S vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12324_ _12348_/A vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__buf_2
XFILLER_103_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12255_ _12255_/A vssd1 vssd1 vccd1 vccd1 _13858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09013__A1 _08573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09013__B2 _08012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06911__B _06942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ _13908_/Q vssd1 vssd1 vccd1 vccd1 _11302_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12186_ _13832_/Q _13059_/B _13111_/B vssd1 vssd1 vccd1 vccd1 _12187_/A sky130_fd_sc_hd__and3b_1
XFILLER_69_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11137_ _13909_/Q vssd1 vssd1 vccd1 vccd1 _11457_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11068_ _11107_/B _11068_/B vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08524__B1 _09000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _10059_/A _10080_/A vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__and2b_1
XFILLER_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12084__B1 _12021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08827__A1 _09132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13709_ _13712_/A _13709_/B vssd1 vssd1 vccd1 vccd1 _13710_/A sky130_fd_sc_hd__and2_1
XANTENNA__08573__B _08573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07230_ _14269_/Q _07229_/X _07236_/S vssd1 vssd1 vccd1 vccd1 _07231_/A sky130_fd_sc_hd__mux2_1
X_07161_ _14104_/Q _07140_/X _07143_/X vssd1 vssd1 vccd1 vccd1 _07161_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07092_ _07090_/X _07091_/X _14362_/Q vssd1 vssd1 vccd1 vccd1 _07093_/S sky130_fd_sc_hd__o21a_1
XANTENNA__12823__B _12952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09802_ _10048_/A _10352_/A vssd1 vssd1 vccd1 vccd1 _10435_/B sky130_fd_sc_hd__xnor2_4
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07994_ _07994_/A _07994_/B vssd1 vssd1 vccd1 vccd1 _08320_/B sky130_fd_sc_hd__xnor2_2
XFILLER_45_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07933__A _14022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06945_ _06945_/A vssd1 vssd1 vccd1 vccd1 _14317_/D sky130_fd_sc_hd__clkbuf_1
X_09733_ _09731_/Y _09697_/A _09739_/B _09732_/X vssd1 vssd1 vccd1 vccd1 _09739_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11455__A _11510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ _07087_/A vssd1 vssd1 vccd1 vccd1 _06970_/A sky130_fd_sc_hd__buf_2
X_09664_ _09649_/Y _09663_/Y _09650_/A vssd1 vssd1 vccd1 vccd1 _09664_/X sky130_fd_sc_hd__a21o_1
XFILLER_28_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08615_ _08615_/A _08615_/B vssd1 vssd1 vccd1 vccd1 _08616_/C sky130_fd_sc_hd__xnor2_1
XFILLER_83_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09595_ _08370_/X _09595_/B vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__and2b_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08546_ _09905_/B vssd1 vssd1 vccd1 vccd1 _08824_/C sky130_fd_sc_hd__clkbuf_2
X_08477_ _13859_/Q vssd1 vssd1 vccd1 vccd1 _09941_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12286__A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07428_ _14088_/Q _07404_/X _07406_/X hold35/X _07417_/X vssd1 vssd1 vccd1 vccd1
+ _07428_/X sky130_fd_sc_hd__a221o_1
XANTENNA__10518__B _10562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ _14100_/Q _07336_/X vssd1 vssd1 vccd1 vccd1 _07359_/X sky130_fd_sc_hd__or2b_1
XFILLER_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ _10377_/B _10370_/B vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__or2_1
XFILLER_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09029_ _09029_/A _09029_/B _09029_/C vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__nand3_2
XFILLER_105_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12040_ _13794_/Q _12038_/X _12039_/X _13810_/Q vssd1 vssd1 vccd1 vccd1 _12041_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12550__A1 _08128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07843__A _14030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13991_ _14441_/CLK _13991_/D vssd1 vssd1 vccd1 vccd1 _13991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08658__B _08658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12942_ _12942_/A _12942_/B vssd1 vssd1 vccd1 vccd1 _12942_/X sky130_fd_sc_hd__or2_1
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _12898_/B vssd1 vssd1 vccd1 vccd1 _12883_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _13997_/Q _11845_/B _12254_/B _14116_/Q vssd1 vssd1 vccd1 vccd1 _11824_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10616__A1 _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12196__A input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ input37/X input36/X input39/X input38/X vssd1 vssd1 vccd1 vccd1 _11756_/B
+ sky130_fd_sc_hd__or4_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08824__D _09084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ _13943_/Q _10708_/B vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11686_ _11686_/A _11686_/B _11686_/C vssd1 vssd1 vccd1 vccd1 _13776_/D sky130_fd_sc_hd__nor3_1
XANTENNA__13566__A0 _12673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13425_ input76/X _14375_/Q _13425_/S vssd1 vssd1 vccd1 vccd1 _13426_/B sky130_fd_sc_hd__mux2_1
X_10637_ _10637_/A vssd1 vssd1 vccd1 vccd1 _10638_/A sky130_fd_sc_hd__inv_2
XANTENNA__12924__A _12924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13356_ _14355_/Q _13265_/A _13355_/X _13343_/X vssd1 vssd1 vccd1 vccd1 _14355_/D
+ sky130_fd_sc_hd__o211a_1
X_10568_ _13962_/Q _10550_/X _10565_/X _10567_/X vssd1 vssd1 vccd1 vccd1 _13962_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_6_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ _12310_/A vssd1 vssd1 vccd1 vccd1 _12307_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13287_ _14418_/Q _13284_/X _13285_/X _13286_/X vssd1 vssd1 vccd1 vccd1 _13287_/X
+ sky130_fd_sc_hd__a211o_1
X_10499_ _10498_/B _10498_/C _10498_/A vssd1 vssd1 vccd1 vccd1 _10507_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12238_ _12239_/A vssd1 vssd1 vccd1 vccd1 _12238_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07548__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12541__A1 _08716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12169_ input94/X vssd1 vssd1 vccd1 vccd1 _12919_/A sky130_fd_sc_hd__buf_6
XFILLER_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_2_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14284_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_65_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput5 dout1[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10855__A1 _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ _08336_/A _08336_/B _08336_/C vssd1 vssd1 vccd1 vccd1 _08400_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_80_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09380_ _08579_/A _09817_/A _09803_/A _09165_/A vssd1 vssd1 vccd1 vccd1 _09382_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_80_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08331_ _08122_/A _08122_/B _08122_/C vssd1 vssd1 vccd1 vccd1 _08331_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07484__B1 _07460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ _08262_/A _08262_/B vssd1 vssd1 vccd1 vccd1 _08263_/B sky130_fd_sc_hd__nand2_1
X_07213_ _14274_/Q _07212_/X _07219_/S vssd1 vssd1 vccd1 vccd1 _07214_/A sky130_fd_sc_hd__mux2_1
X_08193_ _08193_/A _08193_/B vssd1 vssd1 vccd1 vccd1 _08194_/C sky130_fd_sc_hd__nand2_1
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07236__A0 _14267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ _14107_/Q _07140_/X _07143_/X vssd1 vssd1 vccd1 vccd1 _07144_/X sky130_fd_sc_hd__a21o_4
XANTENNA__07928__A _08249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08750__C _09865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07075_ _07051_/X _07074_/X _14364_/Q vssd1 vssd1 vccd1 vccd1 _07076_/S sky130_fd_sc_hd__o21a_1
XFILLER_10_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07977_ _09153_/A vssd1 vssd1 vccd1 vccd1 _08573_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09716_ _09706_/Y _09707_/X _09710_/X _09720_/A vssd1 vssd1 vccd1 vccd1 _09718_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06928_ _06928_/A vssd1 vssd1 vccd1 vccd1 _14319_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09647_ _09651_/A _09652_/A _09647_/C vssd1 vssd1 vccd1 vccd1 _09647_/X sky130_fd_sc_hd__and3b_1
X_06859_ _14400_/Q _06858_/Y _06855_/Y _14403_/Q vssd1 vssd1 vccd1 vccd1 _06875_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_28_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11913__A hold5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09578_ _09573_/Y _09574_/X _09521_/Y _09527_/X vssd1 vssd1 vccd1 vccd1 _09578_/Y
+ sky130_fd_sc_hd__a211oi_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08925__C _08925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08529_/A _08529_/B vssd1 vssd1 vccd1 vccd1 _08530_/B sky130_fd_sc_hd__nor2_1
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11540_ _14053_/Q _13965_/Q vssd1 vssd1 vccd1 vccd1 _11601_/A sky130_fd_sc_hd__or2_1
XFILLER_51_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11471_ _11471_/A _11471_/B vssd1 vssd1 vccd1 vccd1 _11471_/X sky130_fd_sc_hd__or2_1
XFILLER_51_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08941__B _08941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07227__A0 _14270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13210_ _13341_/A vssd1 vssd1 vccd1 vccd1 _13210_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12220__A0 _12218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ _10438_/C _10422_/B vssd1 vssd1 vccd1 vccd1 _10440_/A sky130_fd_sc_hd__or2_1
XFILLER_104_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14190_ _14284_/CLK _14190_/D _12978_/Y vssd1 vssd1 vccd1 vccd1 _14190_/Q sky130_fd_sc_hd__dfrtp_1
X_13141_ _13147_/A vssd1 vssd1 vccd1 vccd1 _13146_/A sky130_fd_sc_hd__clkbuf_4
X_10353_ _10353_/A _10353_/B vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__xnor2_2
XFILLER_87_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13072_ _13072_/A vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input56_A io_wbs_adr[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _10284_/A _10284_/B vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__xnor2_2
XFILLER_105_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12023_ _12026_/A _12023_/B vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__and2_1
XANTENNA__13575__A _13592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13974_ _13982_/CLK _13974_/D _12400_/Y vssd1 vssd1 vccd1 vccd1 _13974_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12925_ _14157_/Q _12915_/X _12924_/X _12920_/X vssd1 vssd1 vccd1 vccd1 _14157_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12919__A _12919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07702__A1 _14147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07702__B2 _14148_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12856_ _13042_/B _12900_/B vssd1 vssd1 vccd1 vccd1 _12885_/A sky130_fd_sc_hd__nor2_2
XFILLER_34_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _13786_/Q _11793_/X _11806_/X vssd1 vssd1 vccd1 vccd1 _11807_/X sky130_fd_sc_hd__a21o_2
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12787_ _14153_/Q _12783_/X _12774_/X _14129_/Q vssd1 vssd1 vccd1 vccd1 _12787_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_38_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09012__B _09153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _13765_/Q _11714_/X _11716_/A _11737_/X vssd1 vssd1 vccd1 vccd1 _13765_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11969__S _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14457_ _14457_/CLK _14457_/D vssd1 vssd1 vccd1 vccd1 _14457_/Q sky130_fd_sc_hd__dfxtp_1
X_11669_ _11669_/A _11682_/C vssd1 vssd1 vccd1 vccd1 _11669_/X sky130_fd_sc_hd__and2_1
XANTENNA__12654__A input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07748__A _14154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13408_ _12561_/X _14370_/Q _13408_/S vssd1 vssd1 vccd1 vccd1 _13409_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14388_ _14440_/CLK _14388_/D vssd1 vssd1 vccd1 vccd1 _14388_/Q sky130_fd_sc_hd__dfxtp_1
X_13339_ _14350_/Q _13332_/X _13338_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _14350_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09963__A _10000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13711__A0 input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13485__A _13485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07900_ _07900_/A _07900_/B vssd1 vssd1 vccd1 vccd1 _07901_/A sky130_fd_sc_hd__or2_1
X_08880_ _08880_/A _08880_/B vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__xor2_1
XFILLER_97_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07831_ _14024_/Q _13970_/Q vssd1 vssd1 vccd1 vccd1 _07918_/A sky130_fd_sc_hd__nand2_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07762_ _07762_/A vssd1 vssd1 vccd1 vccd1 _14061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09501_ _09540_/A _09540_/B _09540_/C vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__and3_1
XFILLER_112_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_0_0_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_io_wbs_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_07693_ _14139_/Q _07744_/A _07673_/X _07692_/X vssd1 vssd1 vccd1 vccd1 _07693_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09432_ _09479_/B _09479_/D _09473_/B _09479_/A vssd1 vssd1 vccd1 vccd1 _09433_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09363_ _09145_/B _09806_/A _09200_/B _09145_/A vssd1 vssd1 vccd1 vccd1 _09364_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13242__A2 _13236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08314_ _08315_/A _08315_/B _08316_/B vssd1 vssd1 vccd1 vccd1 _08322_/B sky130_fd_sc_hd__or3_2
X_09294_ _09294_/A _09294_/B _09294_/C vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__nand3_4
XFILLER_36_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08245_ _08245_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _09771_/A sky130_fd_sc_hd__xnor2_2
X_08176_ _08941_/A vssd1 vssd1 vccd1 vccd1 _08944_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__11556__A2 _13955_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07127_ _14433_/Q _07134_/B _14465_/Q vssd1 vssd1 vccd1 vccd1 _07127_/X sky130_fd_sc_hd__and3b_1
XFILLER_107_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09873__A _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ _14270_/Q _07046_/X _07057_/X _14366_/Q vssd1 vssd1 vccd1 vccd1 _07058_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput150 _14306_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[14] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_40_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput161 _14316_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[24] sky130_fd_sc_hd__buf_2
XFILLER_115_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12505__A1 _14057_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput172 _14297_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[5] sky130_fd_sc_hd__buf_2
XANTENNA__13395__A _13467_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08185__A1 _08937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10971_ _10971_/A vssd1 vssd1 vccd1 vccd1 _10975_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12710_ _12722_/A vssd1 vssd1 vccd1 vccd1 _12715_/A sky130_fd_sc_hd__buf_2
XFILLER_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11492__A1 _08767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13690_ _13724_/A vssd1 vssd1 vccd1 vccd1 _13704_/S sky130_fd_sc_hd__buf_2
XFILLER_71_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12641_ input92/X vssd1 vssd1 vccd1 vccd1 _12641_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13233__A2 _13215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12177__C _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12572_ _12515_/X _14025_/Q _12583_/S vssd1 vssd1 vccd1 vccd1 _12573_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14311_ _14452_/CLK _14311_/D _13180_/Y vssd1 vssd1 vccd1 vccd1 _14311_/Q sky130_fd_sc_hd__dfrtp_4
X_11523_ _11032_/A _11513_/X _11499_/A _11271_/A _11514_/X vssd1 vssd1 vccd1 vccd1
+ _11523_/X sky130_fd_sc_hd__o221a_1
XFILLER_54_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14242_ _14250_/CLK _14242_/D vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
X_11454_ _11454_/A vssd1 vssd1 vccd1 vccd1 _13875_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ _10455_/B _10405_/B vssd1 vssd1 vccd1 vccd1 _10451_/B sky130_fd_sc_hd__and2_1
X_14173_ _14179_/CLK _14173_/D _12958_/Y vssd1 vssd1 vccd1 vccd1 _14173_/Q sky130_fd_sc_hd__dfrtp_1
X_11385_ _13886_/Q _11379_/X _11383_/X _11384_/X vssd1 vssd1 vccd1 vccd1 _13886_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124_ _13128_/A vssd1 vssd1 vccd1 vccd1 _13124_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09783__A _10597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10336_ _09969_/A _10186_/A _09968_/B vssd1 vssd1 vccd1 vccd1 _10350_/B sky130_fd_sc_hd__a21bo_1
XANTENNA_output162_A _14317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ hold29/A _13051_/X _13032_/X vssd1 vssd1 vccd1 vccd1 _13055_/X sky130_fd_sc_hd__a21o_1
X_10267_ _09996_/A _09996_/B _10266_/X vssd1 vssd1 vccd1 vccd1 _10598_/B sky130_fd_sc_hd__o21a_1
XFILLER_61_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12006_ _12006_/A vssd1 vssd1 vccd1 vccd1 _13784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_79_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10198_ _10208_/A _10208_/C _10208_/B vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__a21oi_2
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13957_ _14020_/CLK _13957_/D _12378_/Y vssd1 vssd1 vccd1 vccd1 _13957_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12908_ _14150_/Q _12901_/X _12906_/X _12907_/X vssd1 vssd1 vccd1 vccd1 _14150_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_62_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13888_ _13892_/CLK _13888_/D _12294_/Y vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfrtp_1
X_12839_ _12839_/A vssd1 vssd1 vccd1 vccd1 _14127_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08284__D _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12432__B1 _12485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08030_ _09378_/B vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput30 dout1[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
Xinput41 io_wbs_adr[17] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
Xinput52 io_wbs_adr[27] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_1
Xinput63 io_wbs_adr[8] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput74 io_wbs_datwr[17] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_6
Xinput85 io_wbs_datwr[27] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_2
Xinput96 io_wbs_datwr[8] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07611__A0 _14078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09981_ _10174_/A _10173_/A vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__or2b_1
XFILLER_118_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08932_ _08932_/A _08932_/B vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10632__A _10632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08863_ _09132_/A _09241_/B _09906_/A _08863_/D vssd1 vssd1 vccd1 vccd1 _08864_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07814_ _07878_/A vssd1 vssd1 vccd1 vccd1 _07919_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_85_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08794_ _14009_/Q _08794_/B vssd1 vssd1 vccd1 vccd1 _08798_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07745_ _07744_/Y _14155_/Q _07757_/S vssd1 vssd1 vccd1 vccd1 _07745_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12559__A _12576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07676_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07676_/X sky130_fd_sc_hd__xor2_2
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09415_ _09191_/Y _09192_/Y _09263_/X _09261_/Y vssd1 vssd1 vccd1 vccd1 _09415_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__08890__A2 _10081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _09346_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09360_/A sky130_fd_sc_hd__nand2_2
XFILLER_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09277_ _09277_/A _09277_/B _09277_/C vssd1 vssd1 vccd1 vccd1 _09277_/Y sky130_fd_sc_hd__nand3_1
XFILLER_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08228_ _08170_/A _08170_/Y _08265_/B _08227_/Y vssd1 vssd1 vccd1 vccd1 _08274_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ _08160_/B _08160_/C _08160_/A vssd1 vssd1 vccd1 vccd1 _08170_/A sky130_fd_sc_hd__o21a_1
XFILLER_49_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07602__A0 _14082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11170_ _13923_/Q _13924_/Q _11171_/S vssd1 vssd1 vccd1 vccd1 _11170_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10121_ _10280_/B _10121_/B vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__xnor2_1
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10052_ _10351_/B _10052_/B vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08012__A _08012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13811_ _14335_/CLK _13811_/D vssd1 vssd1 vccd1 vccd1 _13811_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07851__A _14034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input19_A dout1[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13742_ _13745_/A _13742_/B vssd1 vssd1 vccd1 vccd1 _13743_/A sky130_fd_sc_hd__and2_1
X_10954_ _10954_/A _13896_/Q _10679_/A vssd1 vssd1 vccd1 vccd1 _10954_/X sky130_fd_sc_hd__or3b_1
XFILLER_17_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12188__B input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13673_ _13744_/S vssd1 vssd1 vccd1 vccd1 _13687_/S sky130_fd_sc_hd__clkbuf_2
X_10885_ _13974_/Q _10900_/B vssd1 vssd1 vccd1 vccd1 _10885_/X sky130_fd_sc_hd__and2_1
XFILLER_19_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12624_ _12624_/A _12828_/B _12828_/C _12441_/A vssd1 vssd1 vccd1 vccd1 _12669_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_106_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12555_ _12936_/A _08150_/A _12555_/S vssd1 vssd1 vccd1 vccd1 _12556_/B sky130_fd_sc_hd__mux2_1
XFILLER_106_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11506_ _11506_/A _11506_/B vssd1 vssd1 vccd1 vccd1 _11506_/X sky130_fd_sc_hd__and2_1
X_12486_ _12486_/A vssd1 vssd1 vccd1 vccd1 _12486_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10436__B _10436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14225_ _14283_/CLK _14225_/D _13022_/Y vssd1 vssd1 vccd1 vccd1 _14225_/Q sky130_fd_sc_hd__dfrtp_1
X_11437_ _11437_/A vssd1 vssd1 vccd1 vccd1 _11482_/B sky130_fd_sc_hd__inv_2
XANTENNA__12932__A _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14156_ _14158_/CLK _14156_/D vssd1 vssd1 vccd1 vccd1 _14156_/Q sky130_fd_sc_hd__dfxtp_1
X_11368_ _13857_/Q _11536_/A _07904_/A vssd1 vssd1 vccd1 vccd1 _11396_/A sky130_fd_sc_hd__o21a_2
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ _13107_/A vssd1 vssd1 vccd1 vccd1 _14253_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _10393_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10320_/B sky130_fd_sc_hd__or2_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14211_/CLK _14087_/D _12734_/Y vssd1 vssd1 vccd1 vccd1 _14087_/Q sky130_fd_sc_hd__dfrtp_2
X_11299_ _11320_/A _11325_/A _11321_/A vssd1 vssd1 vccd1 vccd1 _11317_/C sky130_fd_sc_hd__o21ba_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13038_ _14232_/Q _13041_/A vssd1 vssd1 vccd1 vccd1 _13038_/X sky130_fd_sc_hd__or2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_41_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14467_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__10248__B1_N _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12379__A _12379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07530_ _14178_/Q _14177_/Q _14176_/Q _14175_/Q _07521_/B vssd1 vssd1 vccd1 vccd1
+ _07530_/X sky130_fd_sc_hd__o41a_1
XFILLER_23_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07461_ _14082_/Q _07459_/X _07460_/X _13882_/Q _07444_/X vssd1 vssd1 vccd1 vccd1
+ _07461_/X sky130_fd_sc_hd__a221o_1
XFILLER_35_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09200_ _14021_/Q _09200_/B vssd1 vssd1 vccd1 vccd1 _09202_/B sky130_fd_sc_hd__and2_1
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07392_ _14210_/Q _14212_/Q _07415_/S vssd1 vssd1 vccd1 vccd1 _07392_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09131_ _09241_/B _09241_/D _09445_/B _09241_/A vssd1 vssd1 vccd1 vccd1 _09133_/A
+ sky130_fd_sc_hd__a22oi_4
X_09062_ _08986_/A _08986_/C _08986_/B vssd1 vssd1 vccd1 vccd1 _09063_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__09200__B _09200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08013_ _08126_/A _08208_/C _08289_/A _08128_/A vssd1 vssd1 vccd1 vccd1 _08020_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09964_ _08980_/B _10487_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10465_/B sky130_fd_sc_hd__o21ba_2
X_08915_ _08915_/A _08915_/B vssd1 vssd1 vccd1 vccd1 _08916_/B sky130_fd_sc_hd__or2_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09895_ _09895_/A _09895_/B vssd1 vssd1 vccd1 vccd1 _09896_/B sky130_fd_sc_hd__nand2_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13673__A _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08846_ _08850_/A _08879_/A _08850_/C vssd1 vssd1 vccd1 vccd1 _08849_/A sky130_fd_sc_hd__nand3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08767__A _08905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__B _11906_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08777_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08781_/B sky130_fd_sc_hd__xnor2_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _07764_/S vssd1 vssd1 vccd1 vccd1 _07757_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07659_ _14070_/Q _07663_/A vssd1 vssd1 vccd1 vccd1 _07660_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10670_ _10777_/B _10670_/B vssd1 vssd1 vccd1 vccd1 _10670_/Y sky130_fd_sc_hd__nand2_2
XFILLER_9_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09329_ _09329_/A _09399_/B _09329_/C _09329_/D vssd1 vssd1 vccd1 vccd1 _09329_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_90_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09812__A1 _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08652__D _09206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _12341_/A vssd1 vssd1 vccd1 vccd1 _12340_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08007__A _08623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ _12273_/A vssd1 vssd1 vccd1 vccd1 _12271_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11907__C1 hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14010_ _14304_/CLK _14010_/D vssd1 vssd1 vccd1 vccd1 _14010_/Q sky130_fd_sc_hd__dfxtp_1
X_11222_ _11294_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__and2_1
XFILLER_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _13918_/Q _13919_/Q _13920_/Q _13921_/Q _11155_/S _11186_/S vssd1 vssd1 vccd1
+ vccd1 _11153_/X sky130_fd_sc_hd__mux4_2
XFILLER_1_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10104_ _10100_/A _10100_/B _10103_/X vssd1 vssd1 vccd1 vccd1 _10106_/B sky130_fd_sc_hd__a21oi_4
X_11084_ _11097_/B _11097_/C _11083_/X vssd1 vssd1 vccd1 vccd1 _11084_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__11087__B _11087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ _09922_/Y _10033_/Y _10034_/Y vssd1 vssd1 vccd1 vccd1 _10354_/B sky130_fd_sc_hd__a21o_1
XFILLER_48_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output125_A _11851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11986_ input55/X vssd1 vssd1 vccd1 vccd1 _12429_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13725_ input83/X _14461_/Q _13738_/S vssd1 vssd1 vccd1 vccd1 _13726_/B sky130_fd_sc_hd__mux2_1
X_10937_ _10971_/A _10932_/X _10934_/X _10765_/A _10936_/X vssd1 vssd1 vccd1 vccd1
+ _11029_/A sky130_fd_sc_hd__o221a_2
XFILLER_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13656_ _13744_/S vssd1 vssd1 vccd1 vccd1 _13670_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10868_ _10868_/A _10868_/B _10874_/A vssd1 vssd1 vccd1 vccd1 _10869_/B sky130_fd_sc_hd__nor3_1
XFILLER_32_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12607_ _12932_/A _14035_/Q _12621_/S vssd1 vssd1 vccd1 vccd1 _12608_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11550__B _13953_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13060__B1 _14240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13587_ _13590_/A _13587_/B vssd1 vssd1 vccd1 vccd1 _13588_/A sky130_fd_sc_hd__and2_1
X_10799_ _10879_/B _10879_/C _10798_/Y vssd1 vssd1 vccd1 vccd1 _10873_/C sky130_fd_sc_hd__a21boi_2
XFILLER_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12538_ _12551_/A _12538_/B vssd1 vssd1 vccd1 vccd1 _12539_/A sky130_fd_sc_hd__and2_1
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12469_ _08842_/A _12465_/X _12454_/X _14047_/Q vssd1 vssd1 vccd1 vccd1 _12469_/X
+ sky130_fd_sc_hd__a22o_1
X_14208_ _14211_/CLK _14208_/D _13001_/Y vssd1 vssd1 vccd1 vccd1 _14208_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10177__B2 _10173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14139_ _14158_/CLK _14139_/D vssd1 vssd1 vccd1 vccd1 _14139_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_99_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08790__A1 _09457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10613__C _10613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06961_ _14458_/Q _14282_/Q vssd1 vssd1 vccd1 vccd1 _06961_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08700_ _08693_/A _08693_/C _08693_/B vssd1 vssd1 vccd1 vccd1 _08701_/C sky130_fd_sc_hd__o21ai_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09680_ _09680_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__or2b_1
X_06892_ _06883_/X _06885_/X _06891_/X _07087_/A vssd1 vssd1 vccd1 vccd1 _07090_/A
+ sky130_fd_sc_hd__o31a_2
X_08631_ _09361_/C vssd1 vssd1 vccd1 vccd1 _08918_/B sky130_fd_sc_hd__buf_6
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08562_ _08568_/A _08562_/B vssd1 vssd1 vccd1 vccd1 _08564_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07513_ hold26/X _14181_/Q _07517_/S vssd1 vssd1 vccd1 vccd1 _07514_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13797__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08493_ _08748_/B vssd1 vssd1 vccd1 vccd1 _08494_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07444_ _07471_/A vssd1 vssd1 vccd1 vccd1 _07444_/X sky130_fd_sc_hd__clkbuf_2
X_07375_ _07399_/A vssd1 vssd1 vccd1 vccd1 _07375_/X sky130_fd_sc_hd__clkbuf_2
X_09114_ _09114_/A _09114_/B _09114_/C vssd1 vssd1 vccd1 vccd1 _09114_/Y sky130_fd_sc_hd__nor3_2
X_09045_ _09045_/A vssd1 vssd1 vccd1 vccd1 _09048_/A sky130_fd_sc_hd__inv_2
XFILLER_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09865__B _09865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11904__A2 _11872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10092__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09947_ _10195_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _10016_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11916__A hold5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09878_ _10039_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _10173_/A sky130_fd_sc_hd__xnor2_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08497__A _09870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08829_ _08829_/A _08829_/B vssd1 vssd1 vccd1 vccd1 _08830_/B sky130_fd_sc_hd__nor2_1
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _14003_/Q _11797_/X _11834_/X _13797_/Q _11839_/X vssd1 vssd1 vccd1 vccd1
+ _11840_/X sky130_fd_sc_hd__a221o_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _13989_/Q _11809_/A _11770_/X _14232_/Q vssd1 vssd1 vccd1 vccd1 _11785_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13510_ _13510_/A vssd1 vssd1 vccd1 vccd1 _14399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _10757_/B _10722_/B vssd1 vssd1 vccd1 vccd1 _10748_/A sky130_fd_sc_hd__nand2_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__B2 _13797_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13441_ _13444_/A _13441_/B vssd1 vssd1 vccd1 vccd1 _13442_/A sky130_fd_sc_hd__and2_1
X_10653_ _10875_/S vssd1 vssd1 vccd1 vccd1 _10836_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_103_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input86_A io_wbs_datwr[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13372_ _13375_/A _13372_/B vssd1 vssd1 vccd1 vccd1 _13373_/A sky130_fd_sc_hd__and2_1
X_10584_ _10576_/C _10582_/Y _10583_/X _10547_/A vssd1 vssd1 vccd1 vccd1 _10584_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ _12385_/A vssd1 vssd1 vccd1 vccd1 _12348_/A sky130_fd_sc_hd__clkbuf_4
X_12254_ _13858_/Q _12254_/B _13037_/C _13111_/B vssd1 vssd1 vccd1 vccd1 _12255_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_119_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09013__A2 _08494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11205_ _11457_/A _11305_/B vssd1 vssd1 vccd1 vccd1 _11311_/B sky130_fd_sc_hd__nand2_1
X_12185_ _12185_/A vssd1 vssd1 vccd1 vccd1 _13111_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11136_ _11134_/A _11110_/X _11135_/X _10826_/X vssd1 vssd1 vccd1 vccd1 _13911_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11067_ _11010_/B _11067_/B vssd1 vssd1 vccd1 vccd1 _11068_/B sky130_fd_sc_hd__and2b_1
XFILLER_27_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08524__A1 _08978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__B2 _08978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10018_ _10092_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _10080_/A sky130_fd_sc_hd__and2_1
XFILLER_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_5_0_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_io_wbs_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_63_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08827__A2 _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ _13772_/Q _13774_/Q _12223_/A vssd1 vssd1 vccd1 vccd1 _11970_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12084__B2 _13822_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13708_ input78/X _14456_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13709_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08573__C _08824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13639_ _13744_/S vssd1 vssd1 vccd1 vccd1 _13653_/S sky130_fd_sc_hd__buf_2
X_07160_ _07160_/A vssd1 vssd1 vccd1 vccd1 _14289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14445__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07091_ _14410_/Q _07098_/B _14442_/Q vssd1 vssd1 vccd1 vccd1 _07091_/X sky130_fd_sc_hd__and3b_1
XANTENNA__12392__A _12410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07015__A1 _14308_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09801_ _09801_/A _09801_/B vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__and2_2
XFILLER_114_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_45_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07993_ _08571_/A _09999_/B vssd1 vssd1 vccd1 vccd1 _07994_/B sky130_fd_sc_hd__nand2_1
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09732_ _09729_/X _09728_/Y _09727_/Y _09727_/B vssd1 vssd1 vccd1 vccd1 _09732_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06944_ _06941_/X _14317_/Q _06944_/S vssd1 vssd1 vccd1 vccd1 _06945_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09206__A _09553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _09663_/A _09663_/B vssd1 vssd1 vccd1 vccd1 _09663_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06875_ _06875_/A _06875_/B _06875_/C vssd1 vssd1 vccd1 vccd1 _07087_/A sky130_fd_sc_hd__or3_4
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08110__A _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08614_ _08905_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _08615_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09594_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09680_/A sky130_fd_sc_hd__nor2_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08545_ _14018_/Q vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _13860_/Q vssd1 vssd1 vccd1 vccd1 _09905_/B sky130_fd_sc_hd__buf_2
XFILLER_39_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08483__C _09491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07427_ _07431_/A _07427_/B vssd1 vssd1 vccd1 vccd1 _07427_/X sky130_fd_sc_hd__or2_1
XANTENNA__10087__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07358_ _14218_/Q _07347_/X _07348_/X _07357_/X vssd1 vssd1 vccd1 vccd1 _14218_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07289_ hold21/X _14229_/Q _07519_/A vssd1 vssd1 vccd1 vccd1 _07290_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11410__S _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09028_ _09025_/Y _09026_/X _08675_/B _08675_/Y vssd1 vssd1 vccd1 vccd1 _09029_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_105_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08754__B2 _08828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13962__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ _14441_/CLK _13990_/D vssd1 vssd1 vccd1 vccd1 _13990_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10550__A _10629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12941_ hold3/A _12928_/X _12940_/X _12934_/X vssd1 vssd1 vccd1 vccd1 _14163_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _12885_/A vssd1 vssd1 vccd1 vccd1 _12872_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _11823_/A vssd1 vssd1 vccd1 vccd1 _11823_/X sky130_fd_sc_hd__buf_2
XFILLER_27_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11754_ input41/X input40/X input43/X input42/X vssd1 vssd1 vccd1 vccd1 _11756_/A
+ sky130_fd_sc_hd__or4_2
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12196__B input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _11216_/A _10705_/B vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__and2_1
X_11685_ _11682_/B _11661_/X _13776_/Q vssd1 vssd1 vccd1 vccd1 _11686_/C sky130_fd_sc_hd__a21oi_1
X_13424_ _13424_/A vssd1 vssd1 vccd1 vccd1 _14374_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09786__A _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10636_ _10636_/A _10636_/B vssd1 vssd1 vccd1 vccd1 _10639_/A sky130_fd_sc_hd__and2_1
XANTENNA__09001__D _09091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355_ _14435_/Q _13216_/X _13354_/X _13341_/X vssd1 vssd1 vccd1 vccd1 _13355_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10567_ _10614_/A _10558_/X _10566_/Y _09788_/A vssd1 vssd1 vccd1 vccd1 _10567_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__06922__B _14287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12306_ _12310_/A vssd1 vssd1 vccd1 vccd1 _12306_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13286_ _14370_/Q _13236_/X _13299_/A vssd1 vssd1 vccd1 vccd1 _13286_/X sky130_fd_sc_hd__a21o_1
X_10498_ _10498_/A _10498_/B _10498_/C vssd1 vssd1 vccd1 vccd1 _10508_/A sky130_fd_sc_hd__and3_1
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ _12239_/A vssd1 vssd1 vccd1 vccd1 _12237_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12940__A _12940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ _13828_/Q _12095_/A _12167_/X _12161_/X vssd1 vssd1 vccd1 vccd1 _13828_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10552__B2 _10551_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12829__A0 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11119_ _11119_/A vssd1 vssd1 vccd1 vccd1 _11119_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_96_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12099_ _12173_/B vssd1 vssd1 vccd1 vccd1 _12112_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 dout1[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09170__A1 _09216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08865__A _08980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08330_ _08391_/A _08391_/B _08391_/C vssd1 vssd1 vccd1 vccd1 _08330_/Y sky130_fd_sc_hd__nor3_1
XFILLER_33_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07484__A1 _14077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ _08262_/A _08262_/B vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__or2_1
XFILLER_119_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07212_ _14090_/Q _13890_/Q _07218_/S vssd1 vssd1 vccd1 vccd1 _07212_/X sky130_fd_sc_hd__mux2_2
XANTENNA__09696__A _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08192_ _08403_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08193_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07236__A1 _07235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07143_ _07186_/A vssd1 vssd1 vccd1 vccd1 _07143_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09630__C1 _09396_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13011__A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__D _13860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _14412_/Q _07098_/B _14444_/Q vssd1 vssd1 vccd1 vccd1 _07074_/X sky130_fd_sc_hd__and3b_1
XFILLER_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08105__A _09234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07976_ _14020_/Q vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _09715_/A _09715_/B _09715_/C vssd1 vssd1 vccd1 vccd1 _09720_/A sky130_fd_sc_hd__or3_1
X_06927_ _06924_/X _14319_/Q _06927_/S vssd1 vssd1 vccd1 vccd1 _06928_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09646_ _09631_/Y _09642_/X _09641_/Y _09404_/X vssd1 vssd1 vccd1 vccd1 _09647_/C
+ sky130_fd_sc_hd__a211o_1
X_06858_ _13779_/Q vssd1 vssd1 vccd1 vccd1 _06858_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _09690_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09577_/X sky130_fd_sc_hd__or2_1
XFILLER_71_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _09241_/A _09241_/B _09074_/B _09206_/B vssd1 vssd1 vccd1 vccd1 _08529_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08459_ _09296_/D vssd1 vssd1 vccd1 vccd1 _09875_/A sky130_fd_sc_hd__buf_4
XFILLER_51_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11470_ _09998_/A _11455_/X _11468_/X _11469_/X vssd1 vssd1 vccd1 vccd1 _13873_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07227__A1 _07226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _10421_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10422_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12220__A1 _07323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10545__A _10562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13140_ _13140_/A vssd1 vssd1 vccd1 vccd1 _13140_/Y sky130_fd_sc_hd__inv_2
X_10352_ _10352_/A _10420_/B vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__xnor2_2
XFILLER_87_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13071_ _13071_/A vssd1 vssd1 vccd1 vccd1 _14243_/D sky130_fd_sc_hd__clkbuf_1
X_10283_ _10283_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10284_/B sky130_fd_sc_hd__xnor2_2
XFILLER_3_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12022_ _13789_/Q _12020_/X _12021_/X _13829_/Q vssd1 vssd1 vccd1 vccd1 _12023_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input49_A io_wbs_adr[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13484__A0 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13973_ _13982_/CLK _13973_/D _12399_/Y vssd1 vssd1 vccd1 vccd1 _13973_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12924_ _12924_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _12924_/X sky130_fd_sc_hd__or2_1
XFILLER_73_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12855_ _12855_/A vssd1 vssd1 vccd1 vccd1 _14132_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _14327_/Q _11833_/A _11770_/X _14235_/Q _11805_/X vssd1 vssd1 vccd1 vccd1
+ _11806_/X sky130_fd_sc_hd__a221o_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _14111_/Q _12782_/X _12784_/X _12785_/X _12207_/X vssd1 vssd1 vccd1 vccd1
+ _14111_/D sky130_fd_sc_hd__o221a_1
XANTENNA__12000__A _12000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11732_/B _11736_/Y _11730_/B _13825_/Q vssd1 vssd1 vccd1 vccd1 _11737_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _14457_/CLK _14456_/D vssd1 vssd1 vccd1 vccd1 _14456_/Q sky130_fd_sc_hd__dfxtp_1
X_11668_ _06855_/Y _11664_/Y _11667_/X vssd1 vssd1 vccd1 vccd1 _13782_/D sky130_fd_sc_hd__o21a_1
X_13407_ _13407_/A vssd1 vssd1 vccd1 vccd1 _14369_/D sky130_fd_sc_hd__clkbuf_1
X_10619_ _10619_/A _10619_/B vssd1 vssd1 vccd1 vccd1 _10619_/Y sky130_fd_sc_hd__xnor2_1
X_14387_ _14467_/CLK _14387_/D vssd1 vssd1 vccd1 vccd1 _14387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11599_ _13854_/Q _11598_/Y _11611_/S vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__mux2_1
X_13338_ _14430_/Q _13327_/X _13337_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13338_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13269_ _14334_/Q _13265_/X _13268_/X _13254_/X vssd1 vssd1 vccd1 vccd1 _14334_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09963__B _09963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07830_ _14026_/Q _13972_/Q vssd1 vssd1 vccd1 vccd1 _07914_/A sky130_fd_sc_hd__nor2_1
XFILLER_97_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13475__A0 _13084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07761_ _14061_/Q _07760_/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07762_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09500_ _09488_/A _09488_/B _09488_/C vssd1 vssd1 vccd1 vccd1 _09540_/C sky130_fd_sc_hd__a21o_1
X_07692_ _14138_/Q _07673_/B _07674_/Y _14137_/Q _07691_/X vssd1 vssd1 vccd1 vccd1
+ _07692_/X sky130_fd_sc_hd__o221a_1
XANTENNA__08595__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09431_ _09479_/A _09479_/B _09479_/D _09473_/B vssd1 vssd1 vccd1 vccd1 _09431_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06901__B1 _06877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ _09362_/A _09844_/B vssd1 vssd1 vccd1 vccd1 _09364_/B sky130_fd_sc_hd__and2_1
XFILLER_36_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09446__A2 _08291_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08313_ _08313_/A _08353_/A vssd1 vssd1 vccd1 vccd1 _08316_/B sky130_fd_sc_hd__and2_1
X_09293_ _09212_/B _09212_/C _09212_/A vssd1 vssd1 vccd1 vccd1 _09294_/C sky130_fd_sc_hd__a21bo_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08244_ _08244_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _08245_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08175_ _14008_/Q vssd1 vssd1 vccd1 vccd1 _08941_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07126_ _14289_/Q _06968_/A _07125_/X _14385_/Q vssd1 vssd1 vccd1 vccd1 _07126_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07057_ _14414_/Q _07056_/Y _07048_/X vssd1 vssd1 vccd1 vccd1 _07057_/X sky130_fd_sc_hd__a21o_1
Xoutput140 _11816_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[5] sky130_fd_sc_hd__buf_2
XFILLER_82_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput151 _14307_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[15] sky130_fd_sc_hd__buf_2
Xoutput162 _14317_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[25] sky130_fd_sc_hd__buf_2
Xoutput173 _14298_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[6] sky130_fd_sc_hd__buf_2
XFILLER_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11067__A_N _11010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07959_ _08132_/A _08251_/A _09848_/A _09842_/A vssd1 vssd1 vccd1 vccd1 _07966_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_101_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13615__S _13628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10970_ _11029_/A _11026_/A _10970_/C _11035_/A vssd1 vssd1 vccd1 vccd1 _11020_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_46_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09629_ _09629_/A _09635_/B vssd1 vssd1 vccd1 vccd1 _09631_/B sky130_fd_sc_hd__xor2_1
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12640_ _12640_/A vssd1 vssd1 vccd1 vccd1 _14043_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ _12571_/A vssd1 vssd1 vccd1 vccd1 _14024_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14310_ _14453_/CLK _14310_/D _13179_/Y vssd1 vssd1 vccd1 vccd1 _14310_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _11517_/A _11521_/Y _11464_/X vssd1 vssd1 vccd1 vccd1 _11522_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07849__A _14033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _14256_/CLK _14241_/D vssd1 vssd1 vccd1 vccd1 _14241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11453_ _10503_/S _11451_/X _11534_/S vssd1 vssd1 vccd1 vccd1 _11454_/A sky130_fd_sc_hd__mux2_1
X_10404_ _10404_/A _10404_/B _10404_/C vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__nand3_1
XFILLER_109_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14172_ _14179_/CLK _14172_/D _12957_/Y vssd1 vssd1 vccd1 vccd1 _14172_/Q sky130_fd_sc_hd__dfrtp_1
X_11384_ _13850_/Q _11390_/B vssd1 vssd1 vccd1 vccd1 _11384_/X sky130_fd_sc_hd__or2_1
X_13123_ _13147_/A vssd1 vssd1 vccd1 vccd1 _13128_/A sky130_fd_sc_hd__buf_2
X_10335_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10337_/A sky130_fd_sc_hd__xnor2_1
XFILLER_65_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _14237_/Q _13041_/X _13052_/X _13053_/X vssd1 vssd1 vccd1 vccd1 _14237_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10266_ _09996_/A _09996_/B _10032_/A _10032_/B vssd1 vssd1 vccd1 vccd1 _10266_/X
+ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_31_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13867_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_output155_A _14292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10722__B _10722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ _12008_/A _12005_/B vssd1 vssd1 vccd1 vccd1 _12006_/A sky130_fd_sc_hd__and2_1
XFILLER_87_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10197_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10208_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13457__A0 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11834__A _11848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13956_ _13963_/CLK _13956_/D _12377_/Y vssd1 vssd1 vccd1 vccd1 _13956_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12907_ _12920_/A vssd1 vssd1 vccd1 vccd1 _12907_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13887_ _14198_/CLK _13887_/D _12291_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12838_ _12847_/A _12838_/B vssd1 vssd1 vccd1 vccd1 _12839_/A sky130_fd_sc_hd__and2_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12432__A1 _08966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12769_ _14108_/Q _12800_/A vssd1 vssd1 vccd1 vccd1 _12769_/X sky130_fd_sc_hd__or2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12432__B2 _14024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput20 dout1[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_2
X_14439_ _14442_/CLK _14439_/D vssd1 vssd1 vccd1 vccd1 _14439_/Q sky130_fd_sc_hd__dfxtp_2
Xinput31 dout1[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__14186__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14164_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput42 io_wbs_adr[18] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput53 io_wbs_adr[28] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_1
Xinput64 io_wbs_adr[9] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
Xinput75 io_wbs_datwr[18] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_4
XFILLER_116_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput86 io_wbs_datwr[28] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput97 io_wbs_datwr[9] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09980_ _09980_/A _09980_/B vssd1 vssd1 vccd1 vccd1 _10290_/A sky130_fd_sc_hd__xor2_2
XFILLER_103_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08931_ _14008_/Q _10061_/A _08928_/A _08940_/A vssd1 vssd1 vccd1 vccd1 _08932_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_69_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10632__B _10632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08862_ _08978_/B _08494_/D _09942_/A _08978_/A vssd1 vssd1 vccd1 vccd1 _08864_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07813_ _07904_/A _07921_/C vssd1 vssd1 vccd1 vccd1 _07878_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13448__A0 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08793_ _08799_/A _08799_/C _08799_/B vssd1 vssd1 vccd1 vccd1 _08820_/B sky130_fd_sc_hd__a21o_1
XFILLER_84_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07744_ _07744_/A vssd1 vssd1 vccd1 vccd1 _07744_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_26_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07675_ _07675_/A _07675_/B vssd1 vssd1 vccd1 vccd1 _07676_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09414_ _09414_/A _09660_/A vssd1 vssd1 vccd1 vccd1 _09421_/C sky130_fd_sc_hd__nor2_2
XFILLER_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09345_ _09345_/A _09345_/B _09345_/C vssd1 vssd1 vccd1 vccd1 _09345_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__09868__B _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09276_ _09276_/A _09276_/B _09276_/C vssd1 vssd1 vccd1 vccd1 _09276_/X sky130_fd_sc_hd__or3_1
X_08227_ _08226_/A _08226_/B _08226_/C vssd1 vssd1 vccd1 vccd1 _08227_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10095__A _10333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ _08195_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08160_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09052__B1 _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07109_ _07109_/A vssd1 vssd1 vccd1 vccd1 _14296_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11919__A hold5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08089_ _14010_/Q vssd1 vssd1 vccd1 vccd1 _08828_/B sky130_fd_sc_hd__buf_2
XFILLER_84_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10120_ _10120_/A _10120_/B _10120_/C vssd1 vssd1 vccd1 vccd1 _10638_/B sky130_fd_sc_hd__and3_1
XANTENNA__13687__A0 _12561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10051_ _10214_/A _10056_/B _10050_/X vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__o21a_1
XFILLER_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13810_ _14335_/CLK _13810_/D vssd1 vssd1 vccd1 vccd1 _13810_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07118__B1 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09658__A2 _09273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13741_ input89/X _14466_/Q _13744_/S vssd1 vssd1 vccd1 vccd1 _13742_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09124__A _13871_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10953_ _10953_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _10953_/X sky130_fd_sc_hd__or2_1
XFILLER_113_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13672_ _13672_/A vssd1 vssd1 vccd1 vccd1 _14445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10884_ _10884_/A _10884_/B _10884_/C vssd1 vssd1 vccd1 vccd1 _10884_/Y sky130_fd_sc_hd__nand3_1
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12623_ _12623_/A vssd1 vssd1 vccd1 vccd1 _14039_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13611__A0 input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12485__A _12485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12554_ _12637_/A vssd1 vssd1 vccd1 vccd1 _12576_/A sky130_fd_sc_hd__buf_2
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11505_ _10215_/A _11486_/X _11503_/X _11504_/X vssd1 vssd1 vccd1 vccd1 _13866_/D
+ sky130_fd_sc_hd__a22o_1
X_12485_ _12485_/A vssd1 vssd1 vccd1 vccd1 _12485_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12178__B1 _11920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14224_ _14224_/CLK _14224_/D _13021_/Y vssd1 vssd1 vccd1 vccd1 _14224_/Q sky130_fd_sc_hd__dfrtp_1
X_11436_ _11294_/A _11002_/B _11436_/S vssd1 vssd1 vccd1 vccd1 _11437_/A sky130_fd_sc_hd__mux2_1
X_14155_ _14158_/CLK _14155_/D vssd1 vssd1 vccd1 vccd1 _14155_/Q sky130_fd_sc_hd__dfxtp_1
X_11367_ _13856_/Q _11377_/B vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__or2_1
XFILLER_99_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06930__B _14286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13106_ _13106_/A _13106_/B vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__and2_1
XFILLER_112_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _10393_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10369_/C sky130_fd_sc_hd__nand2_1
XFILLER_98_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14086_ _14104_/CLK _14086_/D _12733_/Y vssd1 vssd1 vccd1 vccd1 _14086_/Q sky130_fd_sc_hd__dfrtp_2
X_11298_ _11317_/B _11298_/B vssd1 vssd1 vccd1 vccd1 _11321_/A sky130_fd_sc_hd__or2_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _13037_/A _13037_/B _13037_/C vssd1 vssd1 vccd1 vccd1 _13041_/A sky130_fd_sc_hd__and3_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ _10423_/A vssd1 vssd1 vccd1 vccd1 _10395_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13939_ _13947_/CLK _13939_/D _12357_/Y vssd1 vssd1 vccd1 vccd1 _13939_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07460_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07460_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09969__A _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06883__A2 _13778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07391_ _14227_/Q vssd1 vssd1 vccd1 vccd1 _07415_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09130_ _09130_/A _09130_/B _09130_/C vssd1 vssd1 vccd1 vccd1 _09137_/A sky130_fd_sc_hd__nand3_2
XFILLER_31_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09061_ _08435_/A _08684_/A _09060_/A _09060_/C vssd1 vssd1 vccd1 vccd1 _09063_/B
+ sky130_fd_sc_hd__a22o_1
X_08012_ _08012_/A vssd1 vssd1 vccd1 vccd1 _08128_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__07596__A0 _14085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09963_ _10000_/B _09963_/B vssd1 vssd1 vccd1 vccd1 _10276_/B sky130_fd_sc_hd__and2_2
XANTENNA__08113__A _08113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ _08960_/A _08960_/B _08887_/Y _08913_/Y vssd1 vssd1 vccd1 vccd1 _08914_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_44_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09894_ _09894_/A _09897_/B vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__xnor2_4
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08803_/A _08803_/B _08814_/B _08803_/D vssd1 vssd1 vccd1 vccd1 _08850_/C
+ sky130_fd_sc_hd__o22ai_2
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08767__B _08767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08776_ _08776_/A _08776_/B vssd1 vssd1 vccd1 vccd1 _08777_/B sky130_fd_sc_hd__or2_1
XFILLER_38_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ _07727_/A vssd1 vssd1 vccd1 vccd1 _07727_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_66_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07658_ _14145_/Q _07716_/A _07716_/B _14144_/Q _07657_/Y vssd1 vssd1 vccd1 vccd1
+ _07658_/X sky130_fd_sc_hd__o32a_1
XANTENNA__08783__A _08783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07589_ _14088_/Q input4/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07590_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11413__S _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_52_io_wbs_clk_A clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09328_ _09307_/X _09308_/Y _09277_/A _09277_/Y vssd1 vssd1 vccd1 vccd1 _09329_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ _09274_/B _09274_/C _09274_/A vssd1 vssd1 vccd1 vccd1 _09259_/Y sky130_fd_sc_hd__a21oi_2
X_12270_ _12273_/A vssd1 vssd1 vccd1 vccd1 _12270_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11221_ _11221_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11294_/B sky130_fd_sc_hd__xnor2_2
XFILLER_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12580__A0 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _11139_/X _11151_/X _11152_/S vssd1 vssd1 vccd1 vccd1 _11152_/X sky130_fd_sc_hd__mux2_2
XANTENNA__09328__A1 _09307_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ _10143_/B _10143_/A vssd1 vssd1 vccd1 vccd1 _10103_/X sky130_fd_sc_hd__and2b_1
XFILLER_110_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11083_ _11083_/A _11083_/B vssd1 vssd1 vccd1 vccd1 _11083_/X sky130_fd_sc_hd__and2_1
XFILLER_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A dout1[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10034_ _10090_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _10034_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11985_ _13202_/A vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10646__B1 _09788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10936_ _10936_/A _10936_/B vssd1 vssd1 vccd1 vccd1 _10936_/X sky130_fd_sc_hd__or2_1
XFILLER_95_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13724_ _13724_/A vssd1 vssd1 vccd1 vccd1 _13738_/S sky130_fd_sc_hd__buf_2
XANTENNA__07511__A0 hold32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13655_ _13655_/A vssd1 vssd1 vccd1 vccd1 _14440_/D sky130_fd_sc_hd__clkbuf_1
X_10867_ _10867_/A vssd1 vssd1 vccd1 vccd1 _13936_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__06925__B _06942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12606_ _12606_/A vssd1 vssd1 vccd1 vccd1 _14034_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13060__A1 _11990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13586_ input74/X _14421_/Q _13593_/S vssd1 vssd1 vccd1 vccd1 _13587_/B sky130_fd_sc_hd__mux2_1
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10798_ _10873_/B _10798_/B vssd1 vssd1 vccd1 vccd1 _10798_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12537_ _12922_/A _08842_/A _12537_/S vssd1 vssd1 vccd1 vccd1 _12538_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12468_ _13995_/Q _12460_/X _12467_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _13995_/D
+ sky130_fd_sc_hd__o211a_1
X_11419_ _11517_/A _11517_/B vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__or2_1
X_14207_ _14211_/CLK _14207_/D _13000_/Y vssd1 vssd1 vccd1 vccd1 _14207_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12399_ _12403_/A vssd1 vssd1 vccd1 vccd1 _12399_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07578__A0 _14093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14138_ _14158_/CLK _14138_/D vssd1 vssd1 vccd1 vccd1 _14138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14069_ _14075_/CLK _14069_/D _12712_/Y vssd1 vssd1 vccd1 vccd1 _14069_/Q sky130_fd_sc_hd__dfrtp_2
X_06960_ _06960_/A vssd1 vssd1 vccd1 vccd1 _14315_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11126__A1 _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06891_ _06891_/A _06891_/B _06890_/X vssd1 vssd1 vccd1 vccd1 _06891_/X sky130_fd_sc_hd__or3b_1
XFILLER_67_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08630_ _09000_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _08630_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08561_ _08561_/A _08591_/A vssd1 vssd1 vccd1 vccd1 _08562_/B sky130_fd_sc_hd__xnor2_1
XFILLER_78_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07512_ _07512_/A vssd1 vssd1 vccd1 vccd1 _14182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08492_ _13862_/Q vssd1 vssd1 vccd1 vccd1 _08748_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__07502__A0 hold18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07443_ _07458_/A _07443_/B vssd1 vssd1 vccd1 vccd1 _07443_/X sky130_fd_sc_hd__or2_1
XFILLER_74_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13051__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ _07374_/A vssd1 vssd1 vccd1 vccd1 _07399_/A sky130_fd_sc_hd__clkbuf_2
X_09113_ _09110_/X _09111_/Y _09029_/B _09030_/A vssd1 vssd1 vccd1 vccd1 _09114_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07012__A _07090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09044_ _09044_/A _09188_/B vssd1 vssd1 vccd1 vccd1 _09050_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07947__A _13871_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13354__A2 _13236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07569__A0 _14097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12562__A0 _12561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10092__B _10092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10573__C1 _10632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09946_ _09948_/A _09946_/B vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__xnor2_4
XFILLER_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09877_ _09928_/A _10067_/A vssd1 vssd1 vccd1 vccd1 _09947_/B sky130_fd_sc_hd__xnor2_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08828_ _08828_/A _08828_/B _09361_/D _09092_/D vssd1 vssd1 vccd1 vccd1 _08829_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08759_ _08785_/B _08785_/C _08785_/A vssd1 vssd1 vccd1 vccd1 _08760_/C sky130_fd_sc_hd__a21bo_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11932__A input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10628__B1 _10528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11770_ _13035_/A vssd1 vssd1 vccd1 vccd1 _11770_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08944__C _08944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10721_ _10758_/A _10950_/S _10721_/C vssd1 vssd1 vccd1 vccd1 _10722_/B sky130_fd_sc_hd__nor3_4
XANTENNA__09402__A _09402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ input81/X _14379_/Q _13443_/S vssd1 vssd1 vccd1 vccd1 _13441_/B sky130_fd_sc_hd__mux2_1
X_10652_ _10652_/A vssd1 vssd1 vccd1 vccd1 _10652_/X sky130_fd_sc_hd__buf_2
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09797__A1 _08291_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13371_ input91/X _14359_/Q _13374_/S vssd1 vssd1 vccd1 vccd1 _13372_/B sky130_fd_sc_hd__mux2_1
X_10583_ _10583_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _10583_/X sky130_fd_sc_hd__xor2_2
XFILLER_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12322_ _12322_/A vssd1 vssd1 vccd1 vccd1 _12322_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input79_A io_wbs_datwr[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _12259_/A vssd1 vssd1 vccd1 vccd1 _12253_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11356__B2 _10669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11204_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11305_/B sky130_fd_sc_hd__xnor2_2
X_12184_ input65/X _13609_/A vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__and2_1
XFILLER_79_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11135_ _11135_/A _11135_/B vssd1 vssd1 vccd1 vccd1 _11135_/X sky130_fd_sc_hd__or2_1
XFILLER_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14397__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11066_ _11114_/B _11114_/C _11065_/Y vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__a21boi_1
XFILLER_1_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10730__B _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10017_ _10205_/A _10017_/B vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08524__A2 _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12003__A _12021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12938__A _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12084__A2 _12000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ _11968_/A vssd1 vssd1 vccd1 vccd1 _13773_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13707_ _13724_/A vssd1 vssd1 vccd1 vccd1 _13721_/S sky130_fd_sc_hd__clkbuf_2
X_10919_ _11142_/A _11087_/B vssd1 vssd1 vccd1 vccd1 _10920_/A sky130_fd_sc_hd__or2_2
XFILLER_32_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11899_ _13754_/Q _11897_/B _13755_/Q vssd1 vssd1 vccd1 vccd1 _11899_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08573__D _09084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13638_ _13724_/A vssd1 vssd1 vccd1 vccd1 _13744_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13569_ _12610_/X _14416_/Q _13576_/S vssd1 vssd1 vccd1 vccd1 _13570_/B sky130_fd_sc_hd__mux2_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11595__A1 _11592_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07090_ _07090_/A vssd1 vssd1 vccd1 vccd1 _07090_/X sky130_fd_sc_hd__buf_4
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12544__A0 _12926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09800_ _09800_/A _10280_/B vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07992_ _09800_/A vssd1 vssd1 vccd1 vccd1 _09999_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06943_ _06934_/X _06942_/X _14381_/Q vssd1 vssd1 vccd1 vccd1 _06944_/S sky130_fd_sc_hd__o21a_1
X_09731_ _09777_/B _09731_/B vssd1 vssd1 vccd1 vccd1 _09731_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13764__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09662_ _09662_/A _10596_/C vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__or2_1
X_06874_ _14445_/Q _14269_/Q vssd1 vssd1 vccd1 vccd1 _06874_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09206__B _09206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08613_ _08613_/A _08613_/B vssd1 vssd1 vccd1 vccd1 _08616_/B sky130_fd_sc_hd__or2_1
XFILLER_27_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07007__A _07085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09593_ _09593_/A _09593_/B vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08544_ _08726_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _08727_/A sky130_fd_sc_hd__or2_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08279__A1 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08475_ _09378_/B vssd1 vssd1 vccd1 vccd1 _09493_/B sky130_fd_sc_hd__buf_2
X_07426_ _14204_/Q _14206_/Q _07442_/S vssd1 vssd1 vccd1 vccd1 _07427_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07357_ _07349_/X _07355_/X _07356_/X _07352_/X vssd1 vssd1 vccd1 vccd1 _07357_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08451__A1 _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07288_ _07288_/A vssd1 vssd1 vccd1 vccd1 _14230_/D sky130_fd_sc_hd__clkbuf_1
X_09027_ _08675_/B _08675_/Y _09025_/Y _09026_/X vssd1 vssd1 vccd1 vccd1 _09029_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_117_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09892__A _09892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09400__B1 _09319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13618__S _13628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10831__A _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _08893_/A _09807_/X _09806_/X vssd1 vssd1 vccd1 vccd1 _09930_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__08301__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11138__S _11175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12940_ _12940_/A _12940_/B vssd1 vssd1 vccd1 vccd1 _12940_/X sky130_fd_sc_hd__or2_1
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _14137_/Q _12857_/X _12870_/X _12866_/X vssd1 vssd1 vccd1 vccd1 _14137_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11662__A hold6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _13790_/Q _11793_/X _11821_/X vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__a21o_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13263__A1 _14365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _11753_/A vssd1 vssd1 vccd1 vccd1 _11753_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11813__A2 _11808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _11244_/A vssd1 vssd1 vccd1 vccd1 _11216_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11684_ _13777_/Q _11686_/B _11683_/Y vssd1 vssd1 vccd1 vccd1 _13777_/D sky130_fd_sc_hd__o21a_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13423_ _13426_/A _13423_/B vssd1 vssd1 vccd1 vccd1 _13424_/A sky130_fd_sc_hd__and2_1
X_10635_ _10645_/A _10645_/B vssd1 vssd1 vccd1 vccd1 _10636_/B sky130_fd_sc_hd__or2_1
X_13354_ _14387_/Q _13236_/A _13201_/X _14467_/Q vssd1 vssd1 vccd1 vccd1 _13354_/X
+ sky130_fd_sc_hd__a22o_1
X_10566_ _10566_/A _10566_/B vssd1 vssd1 vccd1 vccd1 _10566_/Y sky130_fd_sc_hd__nand2_1
X_12305_ _12317_/A vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__buf_2
XFILLER_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13285_ _14450_/Q _13315_/A _13218_/X _14402_/Q vssd1 vssd1 vccd1 vccd1 _13285_/X
+ sky130_fd_sc_hd__a22o_1
X_10497_ _10503_/S _10497_/B vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__xnor2_1
XFILLER_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11329__B2 _10669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12236_ _12239_/A vssd1 vssd1 vccd1 vccd1 _12236_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12167_ _12917_/A _12173_/B vssd1 vssd1 vccd1 vccd1 _12167_/X sky130_fd_sc_hd__or2_1
XFILLER_110_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11118_ _10831_/X _11114_/C _11117_/Y _11100_/X _11061_/A vssd1 vssd1 vccd1 vccd1
+ _13918_/D sky130_fd_sc_hd__a32o_1
XFILLER_110_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12829__A1 _14125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ _12147_/A vssd1 vssd1 vccd1 vccd1 _12173_/B sky130_fd_sc_hd__clkbuf_1
X_11049_ _11135_/A _11131_/B _11131_/A vssd1 vssd1 vccd1 vccd1 _11129_/A sky130_fd_sc_hd__o21ba_1
XFILLER_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11501__A1 _08836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 dout1[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09170__A2 _09168_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09458__B1 _09792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11291__B _11291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14412__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08260_ _09771_/B _08219_/B _08218_/A vssd1 vssd1 vccd1 vccd1 _08262_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07484__A2 _11746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07211_ _07211_/A vssd1 vssd1 vccd1 vccd1 _14275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08191_ _09635_/A vssd1 vssd1 vccd1 vccd1 _08403_/A sky130_fd_sc_hd__buf_2
XFILLER_118_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07142_ _13893_/Q _07203_/A vssd1 vssd1 vccd1 vccd1 _07186_/A sky130_fd_sc_hd__and2_1
XFILLER_69_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10635__B _10645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07073_ _14268_/Q _07046_/X _07072_/X _14364_/Q vssd1 vssd1 vccd1 vccd1 _07073_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06995__A1 _14278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08138__A2_N _10000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09217__A _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ _09792_/B vssd1 vssd1 vccd1 vccd1 _09445_/B sky130_fd_sc_hd__buf_2
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06926_ _06894_/X _06925_/X _14383_/Q vssd1 vssd1 vccd1 vccd1 _06927_/S sky130_fd_sc_hd__o21a_1
X_09714_ _09692_/Y _09709_/X _09708_/B _09708_/Y vssd1 vssd1 vccd1 vccd1 _09715_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06857_ _14403_/Q _06855_/Y _06856_/Y _14402_/Q vssd1 vssd1 vccd1 vccd1 _06875_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09645_ _09401_/A _09401_/B _09644_/Y vssd1 vssd1 vccd1 vccd1 _09652_/A sky130_fd_sc_hd__o21bai_4
XFILLER_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09576_ _09634_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09576_/X sky130_fd_sc_hd__or2_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07171__S _07183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _09165_/C vssd1 vssd1 vccd1 vccd1 _09074_/B sky130_fd_sc_hd__buf_2
XFILLER_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09887__A _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ _09132_/B vssd1 vssd1 vccd1 vccd1 _08468_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08791__A _08791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07409_ _07399_/X _07402_/X _07407_/X _07408_/X _14209_/Q vssd1 vssd1 vccd1 vccd1
+ _14209_/D sky130_fd_sc_hd__a32o_1
XFILLER_13_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08389_ _08389_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _09698_/C sky130_fd_sc_hd__xnor2_1
XFILLER_104_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10826__A _10826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10420_ _10421_/A _10420_/B vssd1 vssd1 vccd1 vccd1 _10438_/C sky130_fd_sc_hd__and2_1
XFILLER_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10351_ _10384_/A _10351_/B vssd1 vssd1 vccd1 vccd1 _10353_/A sky130_fd_sc_hd__xor2_2
XFILLER_100_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12508__B1 _14007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13070_ _13070_/A _13070_/B vssd1 vssd1 vccd1 vccd1 _13071_/A sky130_fd_sc_hd__and2_1
X_10282_ _10282_/A _10282_/B vssd1 vssd1 vccd1 vccd1 _10284_/A sky130_fd_sc_hd__nor2_2
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12021_ _12021_/A vssd1 vssd1 vccd1 vccd1 _12021_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_21_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14102_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__11657__A _13778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09127__A _09127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08031__A _13875_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13484__A1 _14392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13972_ _13988_/CLK _13972_/D _12397_/Y vssd1 vssd1 vccd1 vccd1 _13972_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__08966__A _08966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12923_ _14156_/Q _12915_/X _12922_/X _12920_/X vssd1 vssd1 vccd1 vccd1 _14156_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _13070_/A _12854_/B vssd1 vssd1 vccd1 vccd1 _12855_/A sky130_fd_sc_hd__and2_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _13992_/Q _11809_/A _11800_/X _14111_/Q vssd1 vssd1 vccd1 vccd1 _11805_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12785_ _14136_/Q _12776_/X _12760_/X vssd1 vssd1 vccd1 vccd1 _12785_/X sky130_fd_sc_hd__a21o_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11736_ _13764_/Q _11740_/B _13765_/Q vssd1 vssd1 vccd1 vccd1 _11736_/Y sky130_fd_sc_hd__o21ai_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ _14457_/CLK _14455_/D vssd1 vssd1 vccd1 vccd1 _14455_/Q sky130_fd_sc_hd__dfxtp_1
X_11667_ _13781_/Q _11669_/A _11661_/X _11680_/D _13782_/Q vssd1 vssd1 vccd1 vccd1
+ _11667_/X sky130_fd_sc_hd__a41o_1
XFILLER_30_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13406_ _13409_/A _13406_/B vssd1 vssd1 vccd1 vccd1 _13407_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_60_io_wbs_clk clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14367_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10618_ _10626_/A _10626_/B _10260_/A vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__o21ai_1
X_14386_ _14467_/CLK _14386_/D vssd1 vssd1 vccd1 vccd1 _14386_/Q sky130_fd_sc_hd__dfxtp_1
X_11598_ _11598_/A _11598_/B vssd1 vssd1 vccd1 vccd1 _11598_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__08206__A _08621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07110__A _14439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13337_ _14382_/Q _13328_/X _13336_/X _14462_/Q vssd1 vssd1 vccd1 vccd1 _13337_/X
+ sky130_fd_sc_hd__a22o_1
X_10549_ _09725_/X _09741_/A _09745_/B _10622_/A vssd1 vssd1 vccd1 vccd1 _10549_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13268_ _14414_/Q _13199_/X _13266_/X _13267_/X vssd1 vssd1 vccd1 vccd1 _13268_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_2_1_0_io_wbs_clk_A clkbuf_2_1_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12219_ _13062_/A _12226_/B vssd1 vssd1 vccd1 vccd1 _12220_/S sky130_fd_sc_hd__or2_1
X_13199_ _13306_/A vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11722__A1 _13829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__A2 _10524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07760_ _07688_/B _14150_/Q _07764_/S vssd1 vssd1 vccd1 vccd1 _07760_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07691_ _14137_/Q _07674_/Y _07676_/X _14136_/Q _07690_/X vssd1 vssd1 vccd1 vccd1
+ _07691_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12398__A _12410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08595__B _08791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09430_ _09430_/A _09430_/B _09430_/C vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__nand3_1
XFILLER_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13227__A1 _14358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09361_ _09361_/A _09361_/B _09361_/C _09361_/D vssd1 vssd1 vccd1 vccd1 _09364_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_21_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08312_ _08312_/A _08982_/B _08313_/A _08312_/D vssd1 vssd1 vccd1 vccd1 _08353_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_75_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09292_ _09291_/A _09291_/C _09291_/B vssd1 vssd1 vccd1 vccd1 _09294_/B sky130_fd_sc_hd__a21o_1
X_08243_ _08243_/A _08243_/B _08243_/C vssd1 vssd1 vccd1 vccd1 _08244_/B sky130_fd_sc_hd__and3_1
XANTENNA__13952__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_57_io_wbs_clk_A clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13022__A _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08174_ _08170_/Y _08171_/X _08084_/Y _08122_/X vssd1 vssd1 vccd1 vccd1 _08194_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07125_ _14433_/Q _07124_/Y _06970_/A vssd1 vssd1 vccd1 vccd1 _07125_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07056_ _14446_/Q _14270_/Q vssd1 vssd1 vccd1 vccd1 _07056_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07955__A _13869_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput130 _11859_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[25] sky130_fd_sc_hd__buf_2
XFILLER_115_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput141 _11819_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[6] sky130_fd_sc_hd__buf_2
Xoutput152 _14308_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[16] sky130_fd_sc_hd__buf_2
XFILLER_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput163 _14318_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[26] sky130_fd_sc_hd__buf_2
Xoutput174 _14299_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[7] sky130_fd_sc_hd__buf_2
XFILLER_0_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11995__C_N input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07958_ _09803_/B vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__buf_4
X_06909_ _14262_/Q _06873_/X _06908_/X _14358_/Q vssd1 vssd1 vccd1 vccd1 _06909_/X
+ sky130_fd_sc_hd__o211a_1
X_07889_ _07847_/A _07847_/B _07847_/C vssd1 vssd1 vccd1 vccd1 _07890_/B sky130_fd_sc_hd__o21a_1
XFILLER_71_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09628_ _09694_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09635_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09559_ _09558_/A _09558_/B _09558_/C vssd1 vssd1 vccd1 vccd1 _09560_/C sky130_fd_sc_hd__a21o_1
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13631__S _13634_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12570_ _12576_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _12571_/A sky130_fd_sc_hd__and2_1
XFILLER_54_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11521_ _11521_/A _11521_/B vssd1 vssd1 vccd1 vccd1 _11521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14240_ _14441_/CLK _14240_/D vssd1 vssd1 vccd1 vccd1 _14240_/Q sky130_fd_sc_hd__dfxtp_1
X_11452_ _11452_/A _11452_/B _07806_/B vssd1 vssd1 vccd1 vccd1 _11534_/S sky130_fd_sc_hd__nor3b_4
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08026__A _09297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ _10404_/B _10404_/C _10404_/A vssd1 vssd1 vccd1 vccd1 _10455_/B sky130_fd_sc_hd__a21o_1
X_14171_ _14179_/CLK _14171_/D _12956_/Y vssd1 vssd1 vccd1 vccd1 _14171_/Q sky130_fd_sc_hd__dfrtp_1
X_11383_ _11396_/A vssd1 vssd1 vccd1 vccd1 _11383_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__06959__A1 _14315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input61_A io_wbs_adr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13122_ _13153_/A vssd1 vssd1 vccd1 vccd1 _13147_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10334_ _10306_/A _10306_/B _10333_/X vssd1 vssd1 vccd1 vccd1 _10349_/B sky130_fd_sc_hd__a21oi_1
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13053_ _13254_/A vssd1 vssd1 vccd1 vccd1 _13053_/X sky130_fd_sc_hd__buf_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _10610_/A _10615_/A _10626_/A _10261_/X _10264_/X vssd1 vssd1 vccd1 vccd1
+ _10598_/A sky130_fd_sc_hd__o41a_1
XFILLER_105_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12004_ _13784_/Q _12000_/X _12003_/X _13824_/Q vssd1 vssd1 vccd1 vccd1 _12005_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10196_ _10206_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10208_/C sky130_fd_sc_hd__nand2_1
XFILLER_61_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output148_A _14304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13825__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13955_ _13963_/CLK _13955_/D _12376_/Y vssd1 vssd1 vccd1 vccd1 _13955_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07136__A1 _14292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12906_ _12906_/A _12913_/B vssd1 vssd1 vccd1 vccd1 _12906_/X sky130_fd_sc_hd__or2_1
XFILLER_59_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13886_ _14198_/CLK _13886_/D _12290_/Y vssd1 vssd1 vccd1 vccd1 _13886_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12633_/X _14127_/Q _12846_/S vssd1 vssd1 vccd1 vccd1 _12838_/B sky130_fd_sc_hd__mux2_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12768_/A _13037_/B _13037_/C vssd1 vssd1 vccd1 vccd1 _12800_/A sky130_fd_sc_hd__and3_2
XANTENNA__12432__A2 _12486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11719_ _13770_/Q _11719_/B vssd1 vssd1 vccd1 vccd1 _11719_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12699_ _14059_/Q _13111_/B _12699_/C vssd1 vssd1 vccd1 vccd1 _12700_/A sky130_fd_sc_hd__and3b_1
X_14438_ _14440_/CLK _14438_/D vssd1 vssd1 vccd1 vccd1 _14438_/Q sky130_fd_sc_hd__dfxtp_1
Xinput10 dout1[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
Xinput21 dout1[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput32 dout1[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput43 io_wbs_adr[19] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
Xinput54 io_wbs_adr[29] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_1
Xinput65 io_wbs_cyc vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_4
X_14369_ _14417_/CLK _14369_/D vssd1 vssd1 vccd1 vccd1 _14369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09061__A1 _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput76 io_wbs_datwr[19] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09061__B2 _09060_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput87 io_wbs_datwr[29] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput98 io_wbs_rst vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__buf_4
XANTENNA__07072__B1 _07048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _08928_/A _08940_/A _14008_/Q _10061_/A vssd1 vssd1 vccd1 vccd1 _08932_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08861_ _08861_/A _08861_/B _08861_/C vssd1 vssd1 vccd1 vccd1 _08872_/A sky130_fd_sc_hd__nand3_1
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07812_ _11362_/A vssd1 vssd1 vccd1 vccd1 _07904_/A sky130_fd_sc_hd__inv_2
X_08792_ _08821_/B _08821_/C _08821_/A vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__a21bo_1
XFILLER_42_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07743_ _07743_/A vssd1 vssd1 vccd1 vccd1 _14067_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13017__A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07674_ _07674_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _07674_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_52_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _09411_/X _09410_/Y _09344_/X _09339_/X vssd1 vssd1 vccd1 vccd1 _09660_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_80_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09344_ _09340_/X _09341_/X _09342_/Y _09343_/X vssd1 vssd1 vccd1 vccd1 _09344_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09275_ _09198_/A _09198_/Y _09229_/X _09230_/Y vssd1 vssd1 vccd1 vccd1 _09275_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08226_ _08226_/A _08226_/B _08226_/C vssd1 vssd1 vccd1 vccd1 _08265_/B sky130_fd_sc_hd__or3_1
XFILLER_20_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08157_ _08223_/C _08157_/B vssd1 vssd1 vccd1 vccd1 _08195_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09884__B _13860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09052__B2 _08925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ _07104_/X _14296_/Q _07108_/S vssd1 vssd1 vccd1 vccd1 _07109_/A sky130_fd_sc_hd__mux2_1
X_08088_ _14011_/Q vssd1 vssd1 vccd1 vccd1 _08796_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07039_ _14448_/Q _14272_/Q vssd1 vssd1 vccd1 vccd1 _07039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10050_ _10124_/B _10050_/B vssd1 vssd1 vccd1 vccd1 _10050_/X sky130_fd_sc_hd__or2_1
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11935__A _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11654__B _13952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13740_ _13740_/A vssd1 vssd1 vccd1 vccd1 _14465_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10952_ _13897_/Q _13898_/Q _11169_/S vssd1 vssd1 vccd1 vccd1 _10953_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13671_ _13678_/A _13671_/B vssd1 vssd1 vccd1 vccd1 _13672_/A sky130_fd_sc_hd__and2_1
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10883_ _10883_/A vssd1 vssd1 vccd1 vccd1 _13933_/D sky130_fd_sc_hd__clkbuf_1
X_12622_ _12635_/A _12622_/B vssd1 vssd1 vccd1 vccd1 _12623_/A sky130_fd_sc_hd__and2_1
XFILLER_40_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12553_ _13428_/A vssd1 vssd1 vccd1 vccd1 _12637_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11504_ _11061_/A _11489_/X _11499_/X _11282_/A _11490_/X vssd1 vssd1 vccd1 vccd1
+ _11504_/X sky130_fd_sc_hd__o221a_1
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ _13999_/Q _12481_/X _12483_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _13999_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12178__A1 _11990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14223_ _14281_/CLK _14223_/D _13020_/Y vssd1 vssd1 vccd1 vccd1 _14223_/Q sky130_fd_sc_hd__dfrtp_1
X_11435_ _11487_/A _11487_/B vssd1 vssd1 vccd1 vccd1 _11482_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14154_ _14158_/CLK _14154_/D vssd1 vssd1 vccd1 vccd1 _14154_/Q sky130_fd_sc_hd__dfxtp_1
X_11366_ _11407_/B vssd1 vssd1 vccd1 vccd1 _11377_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13105_ _12654_/X hold18/A _13105_/S vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__mux2_1
X_10317_ _10366_/A _10317_/B vssd1 vssd1 vccd1 vccd1 _10319_/B sky130_fd_sc_hd__xnor2_1
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11297_ _11297_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__nor2_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _14211_/CLK _14085_/D _12732_/Y vssd1 vssd1 vccd1 vccd1 _14085_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13036_ _13034_/X _14241_/Q _13036_/S vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__mux2_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _08980_/B _10276_/B _10487_/A vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__o21bai_2
XFILLER_26_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10179_ _10188_/A _10188_/B vssd1 vssd1 vccd1 vccd1 _10180_/A sky130_fd_sc_hd__or2_1
XFILLER_93_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13938_ _13943_/CLK _13938_/D _12356_/Y vssd1 vssd1 vccd1 vccd1 _13938_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13869_ _13946_/CLK _13869_/D _12270_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11580__A _14055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07390_ _14094_/Q _07363_/A vssd1 vssd1 vccd1 vccd1 _07390_/X sky130_fd_sc_hd__or2b_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09282__A1 _09425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__A _10206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09060_ _09060_/A _09060_/B _09060_/C vssd1 vssd1 vccd1 vccd1 _09063_/A sky130_fd_sc_hd__nand3_1
X_08011_ _09792_/A vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09962_ _10000_/B _09962_/B vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__nor2_4
XFILLER_83_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08913_ _08957_/A _08957_/B _08912_/A vssd1 vssd1 vccd1 vccd1 _08913_/Y sky130_fd_sc_hd__a21oi_1
X_09893_ _09893_/A _10017_/B vssd1 vssd1 vccd1 vccd1 _09897_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08844_ _08844_/A _08844_/B _08844_/C vssd1 vssd1 vccd1 vccd1 _08879_/A sky130_fd_sc_hd__nor3_2
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11474__B _11533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08775_ _09188_/A _08767_/B _08770_/B _08774_/X vssd1 vssd1 vccd1 vccd1 _08781_/A
+ sky130_fd_sc_hd__a31oi_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _14071_/Q _07720_/X hold2/X _07725_/Y vssd1 vssd1 vccd1 vccd1 _14071_/D sky130_fd_sc_hd__o22a_1
XFILLER_84_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07657_ _14071_/Q _07660_/A vssd1 vssd1 vccd1 vccd1 _07657_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__12586__A _12611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__A _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13054__C1 _13053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07588_ _07588_/A vssd1 vssd1 vccd1 vccd1 _14089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09327_ _09399_/A _09325_/Y _09245_/A _09248_/A vssd1 vssd1 vccd1 vccd1 _09329_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09895__A _09895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ _09258_/A vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__clkbuf_2
X_08209_ _08251_/A vssd1 vssd1 vccd1 vccd1 _09762_/A sky130_fd_sc_hd__clkbuf_4
X_09189_ _09184_/Y _09185_/X _09118_/Y _09110_/X vssd1 vssd1 vccd1 vccd1 _09189_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11220_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13210__A _13341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__A _14023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12580__A1 _14027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _13922_/Q _13923_/Q _13924_/Q _13925_/Q _10967_/S _10777_/B vssd1 vssd1 vccd1
+ vccd1 _11151_/X sky130_fd_sc_hd__mux4_1
X_10102_ _10333_/A _10095_/B _10101_/X vssd1 vssd1 vccd1 vccd1 _10143_/A sky130_fd_sc_hd__a21bo_1
XFILLER_108_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09328__A2 _09308_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11082_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11083_/B sky130_fd_sc_hd__or2_1
X_10033_ _10090_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _10033_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11665__A hold6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input24_A dout1[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11984_ input58/X vssd1 vssd1 vccd1 vccd1 _13202_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13723_ _13723_/A vssd1 vssd1 vccd1 vccd1 _14460_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10646__A1 _10565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10935_ _13902_/Q _13903_/Q _13904_/Q _13905_/Q _10931_/A _13948_/Q vssd1 vssd1 vccd1
+ vccd1 _10936_/B sky130_fd_sc_hd__mux4_1
XFILLER_56_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13654_ _13661_/A _13654_/B vssd1 vssd1 vccd1 vccd1 _13655_/A sky130_fd_sc_hd__and2_1
XFILLER_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10866_ _13936_/Q _10865_/X _10871_/S vssd1 vssd1 vccd1 vccd1 _10867_/A sky130_fd_sc_hd__mux2_1
X_12605_ _12615_/A _12605_/B vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__and2_1
XFILLER_13_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13585_ _13585_/A vssd1 vssd1 vccd1 vccd1 _14420_/D sky130_fd_sc_hd__clkbuf_1
X_10797_ _13933_/Q _10797_/B vssd1 vssd1 vccd1 vccd1 _10798_/B sky130_fd_sc_hd__nor2_1
XFILLER_9_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07102__B _14264_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12551_/A sky130_fd_sc_hd__clkbuf_1
X_12467_ _14030_/Q _12464_/X _12466_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _12467_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_69_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14206_ _14211_/CLK _14206_/D _12999_/Y vssd1 vssd1 vccd1 vccd1 _14206_/Q sky130_fd_sc_hd__dfrtp_1
X_11418_ _11273_/A _11054_/A _11425_/S vssd1 vssd1 vccd1 vccd1 _11517_/B sky130_fd_sc_hd__mux2_1
X_12398_ _12410_/A vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__buf_2
XANTENNA__08214__A _08214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14137_ _14152_/CLK _14137_/D vssd1 vssd1 vccd1 vccd1 _14137_/Q sky130_fd_sc_hd__dfxtp_1
X_11349_ _11271_/A _10845_/X _11348_/X _10669_/X vssd1 vssd1 vccd1 vccd1 _13897_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10582__B1 _10547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14068_ _14075_/CLK _14068_/D _12711_/Y vssd1 vssd1 vccd1 vccd1 _14068_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11126__A2 _11110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13019_ _13022_/A vssd1 vssd1 vccd1 vccd1 _13019_/Y sky130_fd_sc_hd__inv_2
X_06890_ _14393_/Q _11659_/A _06864_/Y _14390_/Q _06889_/Y vssd1 vssd1 vccd1 vccd1
+ _06890_/X sky130_fd_sc_hd__o221a_1
XFILLER_79_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11294__B _11294_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08560_ _08560_/A _08560_/B vssd1 vssd1 vccd1 vccd1 _08591_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07511_ hold32/X _14182_/Q _07517_/S vssd1 vssd1 vccd1 vccd1 _07512_/A sky130_fd_sc_hd__mux2_1
X_08491_ _09297_/A vssd1 vssd1 vccd1 vccd1 _09000_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07442_ _14201_/Q _14203_/Q _07442_/S vssd1 vssd1 vccd1 vccd1 _07443_/B sky130_fd_sc_hd__mux2_1
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07373_ _07373_/A vssd1 vssd1 vccd1 vccd1 _07373_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13051__A2 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09112_ _09029_/B _09030_/A _09110_/X _09111_/Y vssd1 vssd1 vccd1 vccd1 _09114_/B
+ sky130_fd_sc_hd__a211oi_2
X_09043_ _09999_/B vssd1 vssd1 vccd1 vccd1 _09188_/B sky130_fd_sc_hd__buf_6
XFILLER_11_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13030__A _13115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12562__A1 _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09945_ _10039_/A _10171_/B vssd1 vssd1 vccd1 vccd1 _09946_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13511__A0 _12610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ _08494_/D _09807_/X _09806_/X vssd1 vssd1 vccd1 vccd1 _10067_/A sky130_fd_sc_hd__o21a_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07174__S _07183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08827_ _09132_/B _09887_/A _09906_/A _09132_/A vssd1 vssd1 vccd1 vccd1 _08829_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07741__A1 _14156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _08758_/A _08758_/B _08758_/C vssd1 vssd1 vccd1 vccd1 _08785_/A sky130_fd_sc_hd__nand3_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08794__A _14009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__B1 _11823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07709_ _07706_/Y hold3/X _07723_/A vssd1 vssd1 vccd1 vccd1 _07709_/X sky130_fd_sc_hd__mux2_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08689_/A _08966_/C vssd1 vssd1 vccd1 vccd1 _08690_/B sky130_fd_sc_hd__xnor2_2
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13290__A2 _13315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08944__D _08944_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10720_ _10946_/A vssd1 vssd1 vccd1 vccd1 _10721_/C sky130_fd_sc_hd__clkbuf_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10548__B _10565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _10651_/A vssd1 vssd1 vccd1 vccd1 _10652_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13370_ _13370_/A vssd1 vssd1 vccd1 vccd1 _14358_/D sky130_fd_sc_hd__clkbuf_1
X_10582_ _09655_/B _09664_/X _10574_/X _10547_/A vssd1 vssd1 vccd1 vccd1 _10582_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_107_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12763__B _12900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12321_ _12322_/A vssd1 vssd1 vccd1 vccd1 _12321_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12252_ _12252_/A vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__buf_4
XFILLER_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11356__A2 _10845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ _11207_/B _11208_/A _10700_/X vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__a21o_1
X_12183_ _13042_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _13059_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08969__A _09044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ _11134_/A _11134_/B vssd1 vssd1 vccd1 vccd1 _11135_/B sky130_fd_sc_hd__and2_1
XFILLER_62_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11065_ _11111_/B _11065_/B vssd1 vssd1 vccd1 vccd1 _11065_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10016_ _10206_/B _10016_/B vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__xor2_2
XFILLER_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11967_ _13771_/Q _13773_/Q _13184_/A vssd1 vssd1 vccd1 vccd1 _11968_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13281__A2 _13306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13115__A _13115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ _13706_/A vssd1 vssd1 vccd1 vccd1 _14455_/D sky130_fd_sc_hd__clkbuf_1
X_10918_ _10918_/A vssd1 vssd1 vccd1 vccd1 _11142_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11898_ hold31/X _11882_/X _11896_/X _11897_/Y _11885_/X vssd1 vssd1 vccd1 vccd1
+ _13754_/D sky130_fd_sc_hd__o221a_1
XANTENNA__13569__A0 _12610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08209__A _08251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13637_ _13637_/A _13637_/B vssd1 vssd1 vccd1 vccd1 _13724_/A sky130_fd_sc_hd__nand2_2
XFILLER_38_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09237__A1 _08867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10849_ _11322_/A _10840_/B _10846_/X _10848_/Y vssd1 vssd1 vccd1 vccd1 _10849_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13568_ _13568_/A vssd1 vssd1 vccd1 vccd1 _14415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12519_ _12536_/A vssd1 vssd1 vccd1 vccd1 _12534_/A sky130_fd_sc_hd__clkbuf_1
X_13499_ _13502_/A _13499_/B vssd1 vssd1 vccd1 vccd1 _13500_/A sky130_fd_sc_hd__and2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13741__A0 input89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12544__A1 _08632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10555__B1 _10644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07991_ _08070_/C vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__buf_2
XFILLER_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09730_ _09727_/B _09727_/Y _09728_/Y _09729_/X vssd1 vssd1 vccd1 vccd1 _09739_/B
+ sky130_fd_sc_hd__o211ai_4
X_06942_ _14429_/Q _06942_/B _14461_/Q vssd1 vssd1 vccd1 vccd1 _06942_/X sky130_fd_sc_hd__and3b_1
XFILLER_80_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09661_ _10613_/B _09421_/C _10613_/C _09414_/A _09660_/Y vssd1 vssd1 vccd1 vccd1
+ _10596_/C sky130_fd_sc_hd__a311oi_4
X_06873_ _06968_/A vssd1 vssd1 vccd1 vccd1 _06873_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_83_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08612_ _08613_/A _08613_/B vssd1 vssd1 vccd1 vccd1 _08617_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ _09592_/A _09592_/B _09592_/C vssd1 vssd1 vccd1 vccd1 _09592_/Y sky130_fd_sc_hd__nand3_1
X_08543_ _08543_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _08726_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07487__B1 _07528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08474_ _09165_/A _09217_/B _09145_/D _13859_/Q vssd1 vssd1 vccd1 vccd1 _08484_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_39_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08119__A _09590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07425_ _07452_/A vssd1 vssd1 vccd1 vccd1 _07425_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12864__A _12909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07239__A0 _14082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07958__A _09803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ _14217_/Q _14219_/Q _07360_/S vssd1 vssd1 vccd1 vccd1 _07356_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07287_ hold23/X _14230_/Q _07519_/A vssd1 vssd1 vccd1 vccd1 _07288_/A sky130_fd_sc_hd__mux2_1
XANTENNA__08451__A2 _10215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09026_ _09048_/B _09025_/B _09025_/C _09025_/D vssd1 vssd1 vccd1 vccd1 _09026_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13732__A0 input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14028_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09892__B _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08789__A _08789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09928_ _09928_/A vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__buf_2
XFILLER_86_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10849__A1 _11322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09859_ _10091_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__xor2_1
XFILLER_59_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_64_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_46_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11943__A _11947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13634__S _13634_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12870_ _12913_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _12870_/X sky130_fd_sc_hd__or2_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _14331_/Q _11833_/A _11797_/X _13996_/Q _11820_/X vssd1 vssd1 vccd1 vccd1
+ _11821_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _14059_/Q _14258_/Q _11752_/C vssd1 vssd1 vccd1 vccd1 _11753_/A sky130_fd_sc_hd__or3_4
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09132__B _09132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08029__A _14016_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10782_/A vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__buf_2
XFILLER_109_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09219__A1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ _13777_/Q _11686_/B _11686_/A vssd1 vssd1 vccd1 vccd1 _11683_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input91_A io_wbs_datwr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ input75/X _14374_/Q _13425_/S vssd1 vssd1 vccd1 vccd1 _13423_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_50_io_wbs_clk clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14451_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10634_ _10634_/A _10634_/B vssd1 vssd1 vccd1 vccd1 _10634_/Y sky130_fd_sc_hd__nor2_1
X_13353_ _14354_/Q _13265_/A _13352_/X _13343_/X vssd1 vssd1 vccd1 vccd1 _14354_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10565_ _10564_/X _10565_/B _10565_/C vssd1 vssd1 vccd1 vccd1 _10565_/X sky130_fd_sc_hd__and3b_1
XANTENNA__14364__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12304_ _12304_/A vssd1 vssd1 vccd1 vccd1 _12304_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13284_ _13306_/A vssd1 vssd1 vccd1 vccd1 _13284_/X sky130_fd_sc_hd__clkbuf_2
X_10496_ _10496_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__nor2_1
XANTENNA_output178_A _14167_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11329__A2 _10845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12235_ _12239_/A vssd1 vssd1 vccd1 vccd1 _12235_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12166_ input93/X vssd1 vssd1 vccd1 vccd1 _12917_/A sky130_fd_sc_hd__buf_6
XFILLER_69_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11117_ _11062_/X _11117_/B _11117_/C vssd1 vssd1 vccd1 vccd1 _11117_/Y sky130_fd_sc_hd__nand3b_1
X_12097_ _13113_/B _13470_/A _12828_/C vssd1 vssd1 vccd1 vccd1 _12147_/A sky130_fd_sc_hd__or3_4
XFILLER_7_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11048_ _11048_/A _11048_/B _11048_/C vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__and3_1
XFILLER_64_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 dout1[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09458__A1 _08823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12999_ _13003_/A vssd1 vssd1 vccd1 vccd1 _12999_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09458__B2 _08445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07210_ _14275_/Q _07209_/X _07219_/S vssd1 vssd1 vccd1 vccd1 _07211_/A sky130_fd_sc_hd__mux2_1
X_08190_ _09635_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08193_/A sky130_fd_sc_hd__or2_1
XANTENNA__07778__A _10629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10916__B _11087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12765__A1 _14125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07141_ _13839_/Q _13838_/Q vssd1 vssd1 vccd1 vccd1 _07203_/A sky130_fd_sc_hd__nor2_2
XFILLER_119_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07072_ _14412_/Q _07071_/Y _07048_/X vssd1 vssd1 vccd1 vccd1 _07072_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08402__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__A1 _08251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ _13872_/Q vssd1 vssd1 vccd1 vccd1 _09792_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_45_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09713_ _08403_/A _09585_/B _09712_/X vssd1 vssd1 vccd1 vccd1 _09715_/B sky130_fd_sc_hd__o21a_1
XFILLER_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06925_ _14431_/Q _06942_/B _14463_/Q vssd1 vssd1 vccd1 vccd1 _06925_/X sky130_fd_sc_hd__and3b_1
XFILLER_68_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09644_ _09696_/A _09644_/B vssd1 vssd1 vccd1 vccd1 _09644_/Y sky130_fd_sc_hd__nor2_1
X_06856_ _13781_/Q vssd1 vssd1 vccd1 vccd1 _06856_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09575_ _09521_/Y _09527_/X _09573_/Y _09574_/X vssd1 vssd1 vccd1 vccd1 _09575_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08494__D _08494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08526_ _08796_/B vssd1 vssd1 vccd1 vccd1 _09241_/B sky130_fd_sc_hd__buf_2
XFILLER_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08457_ _08796_/B vssd1 vssd1 vccd1 vccd1 _09132_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08791__B _08791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07408_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07408_/X sky130_fd_sc_hd__clkbuf_2
X_08388_ _08388_/A _08388_/B vssd1 vssd1 vccd1 vccd1 _08389_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07339_ _07482_/S vssd1 vssd1 vccd1 vccd1 _07360_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10350_ _10337_/A _10350_/B vssd1 vssd1 vccd1 vccd1 _10360_/B sky130_fd_sc_hd__and2b_1
XFILLER_118_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12508__A1 _11990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ _09009_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08015__C _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10281_ _10280_/B _10281_/B vssd1 vssd1 vccd1 vccd1 _10282_/B sky130_fd_sc_hd__and2b_1
X_12020_ _12059_/A vssd1 vssd1 vccd1 vccd1 _12020_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09408__A _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09127__B _09127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13971_ _13986_/CLK _13971_/D _12396_/Y vssd1 vssd1 vccd1 vccd1 _13971_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08966__B _10486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__A1 _11010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _12922_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__or2_1
XFILLER_4_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12692__A0 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12853_ _12654_/X _14132_/Q _12853_/S vssd1 vssd1 vccd1 vccd1 _12854_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _13194_/A vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08982__A _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12784_ _14152_/Q _12783_/X _12774_/X _14128_/Q vssd1 vssd1 vccd1 vccd1 _12784_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _13763_/Q vssd1 vssd1 vccd1 vccd1 _11740_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14454_ _14457_/CLK _14454_/D vssd1 vssd1 vccd1 vccd1 _14454_/Q sky130_fd_sc_hd__dfxtp_1
X_11666_ hold5/X _14259_/D vssd1 vssd1 vccd1 vccd1 _11680_/D sky130_fd_sc_hd__nor2_1
XANTENNA__13754__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13405_ _12681_/X _14369_/Q _13408_/S vssd1 vssd1 vccd1 vccd1 _13406_/B sky130_fd_sc_hd__mux2_1
X_10617_ _10614_/Y _10616_/Y _13956_/Q _10545_/X vssd1 vssd1 vccd1 vccd1 _13956_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_70_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14385_ _14464_/CLK _14385_/D vssd1 vssd1 vccd1 vccd1 _14385_/Q sky130_fd_sc_hd__dfxtp_1
X_11597_ _11539_/Y _11597_/B vssd1 vssd1 vccd1 vccd1 _11598_/B sky130_fd_sc_hd__and2b_1
X_13336_ _13336_/A vssd1 vssd1 vccd1 vccd1 _13336_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07110__B _14263_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ _10546_/X _10565_/B _10548_/C vssd1 vssd1 vccd1 vccd1 _10548_/X sky130_fd_sc_hd__and3b_1
XFILLER_6_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11848__A _11848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ _14366_/Q _13236_/X _13210_/X vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__a21o_1
X_10479_ _10503_/S _10447_/B _10446_/A vssd1 vssd1 vccd1 vccd1 _10480_/C sky130_fd_sc_hd__a21o_1
X_12218_ input66/X vssd1 vssd1 vccd1 vccd1 _12218_/X sky130_fd_sc_hd__buf_6
XFILLER_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13198_ _13526_/A vssd1 vssd1 vccd1 vccd1 _13306_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12149_ _13822_/Q _12146_/X _12148_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _13822_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09128__B1 _09127_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07690_ _14136_/Q _07676_/X _07680_/Y _07689_/X vssd1 vssd1 vccd1 vccd1 _07690_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08595__C _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13227__A2 _13215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _09360_/A _09360_/B vssd1 vssd1 vccd1 vccd1 _09360_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08103__A1 _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ _09145_/B _09296_/D _09217_/D _09145_/A vssd1 vssd1 vccd1 vccd1 _08312_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09291_ _09291_/A _09291_/B _09291_/C vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__nand3_2
X_08242_ _08243_/B _08243_/C _08243_/A vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__a21oi_1
XFILLER_21_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08173_ _08194_/A vssd1 vssd1 vccd1 vccd1 _08173_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07124_ _14465_/Q _14289_/Q vssd1 vssd1 vccd1 vccd1 _07124_/Y sky130_fd_sc_hd__nand2_1
XFILLER_119_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07055_ _07055_/A vssd1 vssd1 vccd1 vccd1 _14303_/D sky130_fd_sc_hd__clkbuf_1
Xoutput120 _11844_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[16] sky130_fd_sc_hd__buf_2
Xoutput131 _11861_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[26] sky130_fd_sc_hd__buf_2
XFILLER_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput142 _11822_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[7] sky130_fd_sc_hd__buf_2
Xoutput153 _14309_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[17] sky130_fd_sc_hd__buf_2
Xoutput164 _14319_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[27] sky130_fd_sc_hd__buf_2
XANTENNA__11174__A0 _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput175 _14300_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[8] sky130_fd_sc_hd__buf_2
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07971__A _09153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07957_ _13868_/Q vssd1 vssd1 vccd1 vccd1 _09803_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_29_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11477__A1 _10486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ _14406_/Q _06907_/Y _06877_/X vssd1 vssd1 vccd1 vccd1 _06908_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12674__A0 _12673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ _07886_/Y _07887_/X _07890_/A _13979_/Q vssd1 vssd1 vccd1 vccd1 _13979_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09627_ _09360_/A _09360_/B _09626_/X vssd1 vssd1 vccd1 vccd1 _09634_/B sky130_fd_sc_hd__a21oi_2
XFILLER_55_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09558_ _09558_/A _09558_/B _09558_/C vssd1 vssd1 vccd1 vccd1 _09560_/B sky130_fd_sc_hd__nand3_1
X_08509_ _09865_/A vssd1 vssd1 vccd1 vccd1 _09092_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_12_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09489_ _09489_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09499_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ _10061_/A _11510_/X _11518_/X _11519_/X vssd1 vssd1 vccd1 vccd1 _13863_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_1_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14244_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11451_ _11451_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11451_/X sky130_fd_sc_hd__xor2_1
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _10430_/S _10429_/A vssd1 vssd1 vccd1 vccd1 _10404_/A sky130_fd_sc_hd__xor2_1
X_14170_ _14258_/CLK _14170_/D vssd1 vssd1 vccd1 vccd1 _14170_/Q sky130_fd_sc_hd__dfxtp_1
X_11382_ _13887_/Q _11379_/X _11370_/X _11381_/X vssd1 vssd1 vccd1 vccd1 _13887_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13121_ _13121_/A vssd1 vssd1 vccd1 vccd1 _13121_/Y sky130_fd_sc_hd__inv_2
X_10333_ _10333_/A _10333_/B vssd1 vssd1 vccd1 vccd1 _10333_/X sky130_fd_sc_hd__and2_1
XFILLER_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input54_A io_wbs_adr[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ hold25/A _13051_/X _13032_/X vssd1 vssd1 vccd1 vccd1 _13052_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10264_ _10610_/A _10615_/A _10263_/Y vssd1 vssd1 vccd1 vccd1 _10264_/X sky130_fd_sc_hd__or3b_1
XFILLER_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08042__A _09491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ _12021_/A vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10195_ _10195_/A _10195_/B vssd1 vssd1 vccd1 vccd1 _10204_/A sky130_fd_sc_hd__xnor2_1
XFILLER_105_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08581__A1 _09493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08581__B2 _09443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11607__S _11611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12665__A0 _12664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13954_ _13963_/CLK _13954_/D _12375_/Y vssd1 vssd1 vccd1 vccd1 _13954_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12905_ _14149_/Q _12901_/X _12904_/X _12892_/X vssd1 vssd1 vccd1 vccd1 _14149_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13885_ _14198_/CLK _13885_/D _12289_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12836_ _12836_/A vssd1 vssd1 vccd1 vccd1 _14126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12767_ hold12/A _12761_/X _12766_/X vssd1 vssd1 vccd1 vccd1 _12767_/X sky130_fd_sc_hd__o21a_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _11730_/B vssd1 vssd1 vccd1 vccd1 _11718_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12698_ _12703_/A vssd1 vssd1 vccd1 vccd1 _12698_/Y sky130_fd_sc_hd__inv_2
X_14437_ _14451_/CLK _14437_/D vssd1 vssd1 vccd1 vccd1 _14437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11649_ _11649_/A vssd1 vssd1 vccd1 vccd1 _13842_/D sky130_fd_sc_hd__clkbuf_1
Xinput11 dout1[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 dout1[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_2
Xinput33 io_wbs_adr[0] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
Xinput44 io_wbs_adr[1] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_4
Xinput55 io_wbs_adr[2] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_2
X_14368_ _14417_/CLK _14368_/D vssd1 vssd1 vccd1 vccd1 _14368_/Q sky130_fd_sc_hd__dfxtp_1
Xinput66 io_wbs_datwr[0] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_4
XFILLER_7_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput77 io_wbs_datwr[1] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__buf_2
Xinput88 io_wbs_datwr[2] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_8
X_13319_ _14378_/Q _13307_/X _13315_/X _14458_/Q vssd1 vssd1 vccd1 vccd1 _13319_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11578__A _14054_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput99 io_wbs_stb vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__buf_6
X_14299_ _14411_/CLK _14299_/D _13165_/Y vssd1 vssd1 vccd1 vccd1 _14299_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11297__B _11297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ _08944_/C _10215_/A vssd1 vssd1 vccd1 vccd1 _08880_/A sky130_fd_sc_hd__nand2_1
XFILLER_85_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07811_ _07808_/X _07810_/Y _07807_/Y vssd1 vssd1 vccd1 vccd1 _13986_/D sky130_fd_sc_hd__o21ba_1
XFILLER_85_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08791_ _08791_/A _08791_/B _09905_/B _09941_/B vssd1 vssd1 vccd1 vccd1 _08821_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_78_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07742_ _14067_/Q _07741_/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07743_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07673_ _14138_/Q _07673_/B vssd1 vssd1 vccd1 vccd1 _07673_/X sky130_fd_sc_hd__and2_1
XFILLER_25_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09412_ _09339_/X _09344_/X _09410_/Y _09411_/X vssd1 vssd1 vccd1 vccd1 _09414_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13081__A0 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _09338_/X _09337_/Y _09274_/Y _09274_/B vssd1 vssd1 vccd1 vccd1 _09343_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09274_ _09274_/A _09274_/B _09274_/C vssd1 vssd1 vccd1 vccd1 _09274_/Y sky130_fd_sc_hd__nand3_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ _09685_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08226_/C sky130_fd_sc_hd__xnor2_1
XFILLER_119_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08156_ _08201_/A _08156_/B vssd1 vssd1 vccd1 vccd1 _08157_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07107_ _07090_/X _07106_/X _14360_/Q vssd1 vssd1 vccd1 vccd1 _07108_/S sky130_fd_sc_hd__o21a_1
X_08087_ _14011_/Q _08796_/B _08097_/B vssd1 vssd1 vccd1 vccd1 _08091_/A sky130_fd_sc_hd__and3_2
XANTENNA__07177__S _07183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07038_ _07038_/A vssd1 vssd1 vccd1 vccd1 _14305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08989_ _08989_/A _08989_/B _08989_/C vssd1 vssd1 vccd1 vccd1 _08991_/B sky130_fd_sc_hd__nand3_4
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13208__A _13236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12647__A0 _12645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12112__A _12936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10951_ _10951_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _10963_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13670_ _12664_/X _14445_/Q _13670_/S vssd1 vssd1 vccd1 vccd1 _13671_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10882_ _13933_/Q _10881_/Y _10897_/S vssd1 vssd1 vccd1 vccd1 _10883_/A sky130_fd_sc_hd__mux2_1
X_12621_ _12942_/A _14039_/Q _12621_/S vssd1 vssd1 vccd1 vccd1 _12622_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09421__A _10621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ _12552_/A vssd1 vssd1 vccd1 vccd1 _14019_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08037__A _08097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11503_ _11497_/A _11502_/X _11472_/X vssd1 vssd1 vccd1 vccd1 _11503_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12483_ _14034_/Q _12464_/X _12482_/X _12473_/X vssd1 vssd1 vccd1 vccd1 _12483_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_11_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14222_ _14244_/CLK _14222_/D _13019_/Y vssd1 vssd1 vccd1 vccd1 _14222_/Q sky130_fd_sc_hd__dfrtp_1
X_11434_ _11291_/A _11007_/B _11446_/S vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07054__A1 _14303_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14153_ _14158_/CLK _14153_/D vssd1 vssd1 vccd1 vccd1 _14153_/Q sky130_fd_sc_hd__dfxtp_1
X_11365_ _11365_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _11407_/B sky130_fd_sc_hd__nor2_2
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13104_ _13104_/A vssd1 vssd1 vccd1 vccd1 _14252_/D sky130_fd_sc_hd__clkbuf_1
X_10316_ _10293_/A _10293_/B _10315_/X vssd1 vssd1 vccd1 vccd1 _10317_/B sky130_fd_sc_hd__a21o_1
XFILLER_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11138__A0 _10912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14084_ _14211_/CLK _14084_/D _12731_/Y vssd1 vssd1 vccd1 vccd1 _14084_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_output160_A _14315_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11296_ _11324_/B _11324_/C _11324_/A vssd1 vssd1 vccd1 vccd1 _11325_/A sky130_fd_sc_hd__a21oi_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _13035_/A _13203_/B vssd1 vssd1 vccd1 vccd1 _13036_/S sky130_fd_sc_hd__and2_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10247_ _10250_/A _10250_/B vssd1 vssd1 vccd1 vccd1 _10254_/A sky130_fd_sc_hd__or2_1
XFILLER_78_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10178_ _10178_/A vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__inv_2
XFILLER_26_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06939__B _14285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12638__A0 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13937_ _13943_/CLK _13937_/D _12353_/Y vssd1 vssd1 vccd1 vccd1 _13937_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13552__S _13559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06868__B2 _14397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13868_ _13946_/CLK _13868_/D _12269_/Y vssd1 vssd1 vccd1 vccd1 _13868_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12819_ hold3/X _12772_/X _12803_/A _14147_/Q _12809_/X vssd1 vssd1 vccd1 vccd1 _12819_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__13063__A0 _12218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13799_ _14400_/CLK _13799_/D vssd1 vssd1 vccd1 vccd1 _13799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14448__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08010_ _13873_/Q vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _10091_/A _10195_/A vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__or2_1
XFILLER_103_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08912_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _08957_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09892_ _09892_/A _10083_/A vssd1 vssd1 vccd1 vccd1 _10017_/B sky130_fd_sc_hd__xnor2_4
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08843_ _08834_/A _08834_/C _08834_/B vssd1 vssd1 vccd1 vccd1 _08844_/C sky130_fd_sc_hd__a21oi_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08774_ _08769_/B _08774_/B vssd1 vssd1 vccd1 vccd1 _08774_/X sky130_fd_sc_hd__and2b_1
XFILLER_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ _07657_/Y _07723_/X _07724_/X vssd1 vssd1 vccd1 vccd1 _07725_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_69_io_wbs_clk_A clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_38_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07656_ _07656_/A _07656_/B vssd1 vssd1 vccd1 vccd1 _07700_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09241__A _09241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07587_ _14089_/Q input5/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07588_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09326_ _09245_/A _09248_/A _09399_/A _09325_/Y vssd1 vssd1 vccd1 vccd1 _09399_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_16_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09257_ _09274_/A _09258_/A _09274_/C vssd1 vssd1 vccd1 vccd1 _09257_/X sky130_fd_sc_hd__and3_1
X_08208_ _08249_/A _08208_/B _08208_/C _09963_/B vssd1 vssd1 vccd1 vccd1 _08208_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09188_ _09188_/A _09188_/B _09188_/C vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__and3_2
XANTENNA__11907__A2 _11872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ _08213_/B _08203_/B vssd1 vssd1 vccd1 vccd1 _08141_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08784__A1 _08842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__A _11240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08784__B2 _08716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _10971_/A _11145_/X _11147_/X _10765_/A _11149_/X vssd1 vssd1 vccd1 vccd1
+ _11249_/A sky130_fd_sc_hd__o221a_1
XFILLER_108_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10101_ _10101_/A _10333_/B vssd1 vssd1 vccd1 vccd1 _10101_/X sky130_fd_sc_hd__or2b_1
XANTENNA__11946__A _11947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11081_ _11099_/B _11099_/C _11080_/X vssd1 vssd1 vccd1 vccd1 _11097_/C sky130_fd_sc_hd__a21bo_1
XFILLER_1_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10032_ _10032_/A _10032_/B vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__xnor2_2
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input17_A dout1[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ _12762_/C _12951_/A _11766_/B vssd1 vssd1 vccd1 vccd1 _11994_/A sky130_fd_sc_hd__or3b_1
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13722_ _13729_/A _13722_/B vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__and2_1
X_10934_ _10713_/A _10933_/X _10916_/X vssd1 vssd1 vccd1 vccd1 _10934_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13653_ input92/X _14440_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13654_/B sky130_fd_sc_hd__mux2_1
X_10865_ _11119_/A _10858_/C _10863_/X _10864_/X vssd1 vssd1 vccd1 vccd1 _10865_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12604_ _12930_/A _14034_/Q _12621_/S vssd1 vssd1 vccd1 vccd1 _12605_/B sky130_fd_sc_hd__mux2_1
X_13584_ _13590_/A _13584_/B vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__and2_1
X_10796_ _10884_/B _10884_/C _10884_/A vssd1 vssd1 vccd1 vccd1 _10879_/C sky130_fd_sc_hd__a21o_1
XFILLER_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12535_ _12535_/A vssd1 vssd1 vccd1 vccd1 _14014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_71_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12466_ _08983_/A _12465_/X _12454_/X _14046_/Q vssd1 vssd1 vccd1 vccd1 _12466_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14205_ _14211_/CLK _14205_/D _12997_/Y vssd1 vssd1 vccd1 vccd1 _14205_/Q sky130_fd_sc_hd__dfrtp_1
X_11417_ _11521_/A _11521_/B vssd1 vssd1 vccd1 vccd1 _11517_/A sky130_fd_sc_hd__or2_1
X_12397_ _12397_/A vssd1 vssd1 vccd1 vccd1 _12397_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08775__A1 _09188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14136_ _14152_/CLK _14136_/D vssd1 vssd1 vccd1 vccd1 _14136_/Q sky130_fd_sc_hd__dfxtp_1
X_11348_ _11348_/A _11348_/B vssd1 vssd1 vccd1 vccd1 _11348_/X sky130_fd_sc_hd__xor2_1
XFILLER_113_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14067_ _14179_/CLK _14067_/D _12709_/Y vssd1 vssd1 vccd1 vccd1 _14067_/Q sky130_fd_sc_hd__dfrtp_1
X_11279_ _11279_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__or2_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13018_ _13022_/A vssd1 vssd1 vccd1 vccd1 _13018_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08230__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ _07510_/A vssd1 vssd1 vccd1 vccd1 _14183_/D sky130_fd_sc_hd__clkbuf_1
X_08490_ _08555_/B _09085_/B _09084_/C _08580_/A vssd1 vssd1 vccd1 vccd1 _08490_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_74_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10919__B _11087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07441_ _07425_/X _07439_/X _07440_/X _07435_/X _14203_/Q vssd1 vssd1 vccd1 vccd1
+ _14203_/D sky130_fd_sc_hd__a32o_1
XFILLER_90_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07372_ _14215_/Q _07347_/X _07348_/X _07371_/X vssd1 vssd1 vccd1 vccd1 _14215_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10000__A _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09111_ _09118_/A _09110_/C _09110_/A vssd1 vssd1 vccd1 vccd1 _09111_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09042_ _08973_/A _08973_/B _09041_/X vssd1 vssd1 vccd1 vccd1 _09114_/A sky130_fd_sc_hd__o21a_1
XANTENNA__13311__A _13332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12011__B2 _13826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10573__A1 _10644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09944_ _09893_/A _10191_/B _10173_/B vssd1 vssd1 vccd1 vccd1 _09948_/A sky130_fd_sc_hd__a21oi_4
X_09875_ _09875_/A _09875_/B vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__xnor2_4
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A dout1[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _09134_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08830_/A sky130_fd_sc_hd__nand2_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08757_ _08757_/A _08757_/B vssd1 vssd1 vccd1 vccd1 _08785_/C sky130_fd_sc_hd__xnor2_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08794__B _08794_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _07764_/S vssd1 vssd1 vccd1 vccd1 _07723_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _08688_/A _08688_/B vssd1 vssd1 vccd1 vccd1 _08966_/C sky130_fd_sc_hd__nor2_1
XFILLER_54_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ _07671_/B _07672_/B _07671_/A vssd1 vssd1 vccd1 vccd1 _07670_/A sky130_fd_sc_hd__a21boi_2
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10650_ _10650_/A vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__buf_2
XFILLER_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12786__C1 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ _09277_/A _09277_/Y _09307_/X _09308_/Y vssd1 vssd1 vccd1 vccd1 _09329_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_10_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10581_ _10581_/A vssd1 vssd1 vccd1 vccd1 _13961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13221__A _13341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12320_ _12322_/A vssd1 vssd1 vccd1 vccd1 _12320_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12251_ _12251_/A vssd1 vssd1 vccd1 vccd1 _12251_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11202_ _10652_/X _11185_/X _11143_/X vssd1 vssd1 vccd1 vccd1 _11208_/A sky130_fd_sc_hd__o21ai_2
X_12182_ _12952_/B vssd1 vssd1 vccd1 vccd1 _12828_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08969__B _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _11048_/A _11110_/X _11132_/Y _10826_/X vssd1 vssd1 vccd1 vccd1 _13912_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09146__A _09362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11064_ _11014_/B _11064_/B vssd1 vssd1 vccd1 vccd1 _11065_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08050__A _08146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10015_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10111_/A sky130_fd_sc_hd__nand2_1
XFILLER_92_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output123_A _11850_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11966_ _13153_/A vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__buf_6
XFILLER_45_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12300__A _12304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10917_ _10761_/B _10914_/X _10916_/X vssd1 vssd1 vccd1 vccd1 _10917_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13705_ _13712_/A _13705_/B vssd1 vssd1 vccd1 vccd1 _13706_/A sky130_fd_sc_hd__and2_1
X_11897_ _13754_/Q _11897_/B vssd1 vssd1 vccd1 vccd1 _11897_/Y sky130_fd_sc_hd__nor2_1
X_13636_ _13636_/A vssd1 vssd1 vccd1 vccd1 _14435_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07113__B _07134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10848_ _13981_/Q _10906_/A vssd1 vssd1 vccd1 vccd1 _10848_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09237__A2 _09824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13567_ _13573_/A _13567_/B vssd1 vssd1 vccd1 vccd1 _13568_/A sky130_fd_sc_hd__and2_1
X_10779_ _10905_/B _10783_/A _10782_/A vssd1 vssd1 vccd1 vccd1 _10780_/B sky130_fd_sc_hd__o21ai_1
XFILLER_34_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12518_ _12518_/A vssd1 vssd1 vccd1 vccd1 _14009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13498_ _12660_/X _14396_/Q _13511_/S vssd1 vssd1 vccd1 vccd1 _13499_/B sky130_fd_sc_hd__mux2_1
X_12449_ _08891_/A _12439_/X _12442_/X _14043_/Q vssd1 vssd1 vccd1 vccd1 _12449_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14119_ _14163_/CLK _14119_/D vssd1 vssd1 vccd1 vccd1 _14119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07990_ _09821_/B vssd1 vssd1 vccd1 vccd1 _08070_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_113_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06941_ _14285_/Q _06929_/X _06940_/X _14381_/Q vssd1 vssd1 vccd1 vccd1 _06941_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09660_ _09660_/A _10604_/A vssd1 vssd1 vccd1 vccd1 _09660_/Y sky130_fd_sc_hd__nor2_1
X_06872_ _07027_/A vssd1 vssd1 vccd1 vccd1 _06968_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08611_ _08611_/A _08620_/A vssd1 vssd1 vccd1 vccd1 _08613_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09591_ _09591_/A _09670_/B vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__xnor2_1
XFILLER_82_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ _08571_/A _08783_/A vssd1 vssd1 vccd1 vccd1 _08726_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13306__A _13306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12210__A _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09476__A2 _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08473_ _13860_/Q vssd1 vssd1 vccd1 vccd1 _09145_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07424_ _07399_/X _07422_/X _07423_/X _07408_/X _14206_/Q vssd1 vssd1 vccd1 vccd1
+ _14206_/D sky130_fd_sc_hd__a32o_1
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14016__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07355_ _14101_/Q _07336_/X vssd1 vssd1 vccd1 vccd1 _07355_/X sky130_fd_sc_hd__or2b_1
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07286_ _07286_/A vssd1 vssd1 vccd1 vccd1 _14231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09025_ _09048_/B _09025_/B _09025_/C _09025_/D vssd1 vssd1 vccd1 vccd1 _09025_/Y
+ sky130_fd_sc_hd__nand4_4
XANTENNA__07974__A _13872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _10271_/A _10331_/A vssd1 vssd1 vccd1 vccd1 _10394_/B sky130_fd_sc_hd__xor2_4
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09858_ _08703_/B _09843_/X _09844_/X vssd1 vssd1 vccd1 vccd1 _10090_/B sky130_fd_sc_hd__a21oi_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08809_ _08814_/B _08809_/B vssd1 vssd1 vccd1 vccd1 _08815_/C sky130_fd_sc_hd__xnor2_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09789_ _10634_/A _10485_/A _09788_/X vssd1 vssd1 vccd1 vccd1 _09789_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_74_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11820_ _14239_/Q _13037_/A _11800_/X _14115_/Q vssd1 vssd1 vccd1 vccd1 _11820_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13216__A _13526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12120__A _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11751_ _14257_/Q _13858_/Q _13832_/Q _14170_/Q vssd1 vssd1 vccd1 vccd1 _11752_/C
+ sky130_fd_sc_hd__or4_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09132__C _09792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13650__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _13944_/Q vssd1 vssd1 vccd1 vccd1 _10782_/A sky130_fd_sc_hd__inv_2
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _13776_/Q _11682_/B _11682_/C vssd1 vssd1 vccd1 vccd1 _11686_/B sky130_fd_sc_hd__and3_1
XFILLER_109_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09219__A2 _09803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13421_ _13421_/A vssd1 vssd1 vccd1 vccd1 _14373_/D sky130_fd_sc_hd__clkbuf_1
X_10633_ _10633_/A _10633_/B vssd1 vssd1 vccd1 vccd1 _10634_/B sky130_fd_sc_hd__xnor2_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13352_ _14434_/Q _13216_/X _13351_/X _13341_/X vssd1 vssd1 vccd1 vccd1 _13352_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_input84_A io_wbs_datwr[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ _10564_/A _10564_/B _10564_/C vssd1 vssd1 vccd1 vccd1 _10564_/X sky130_fd_sc_hd__and3_1
XANTENNA__08045__A _14018_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _12304_/A vssd1 vssd1 vccd1 vccd1 _12303_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13283_ _14337_/Q _13265_/X _13282_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _14337_/D
+ sky130_fd_sc_hd__o211a_1
X_10495_ _10495_/A _10495_/B vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__and2_1
XFILLER_68_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12234_ _12252_/A vssd1 vssd1 vccd1 vccd1 _12239_/A sky130_fd_sc_hd__buf_2
XFILLER_29_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12931__C1 _12920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12165_ _13827_/Q _12095_/A _12164_/X _12161_/X vssd1 vssd1 vccd1 vccd1 _13827_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11116_ _11014_/B _11110_/X _11114_/Y _11115_/Y vssd1 vssd1 vccd1 vccd1 _13919_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12096_ input96/X vssd1 vssd1 vccd1 vccd1 _12924_/A sky130_fd_sc_hd__buf_4
XFILLER_104_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11047_ _11048_/B _11048_/C _11048_/A vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__a21oi_1
XFILLER_77_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 dout1[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09458__A2 _09821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12998_ _13004_/A vssd1 vssd1 vccd1 vccd1 _13003_/A sky130_fd_sc_hd__buf_2
XFILLER_75_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12462__A1 _14029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _11953_/A vssd1 vssd1 vccd1 vccd1 _11949_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13619_ _13625_/A _13619_/B vssd1 vssd1 vccd1 vccd1 _13620_/A sky130_fd_sc_hd__and2_1
XANTENNA__14189__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12765__A2 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ _07185_/A vssd1 vssd1 vccd1 vccd1 _07140_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ _14444_/Q _14268_/Q vssd1 vssd1 vccd1 vccd1 _07071_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07973_ _09457_/D vssd1 vssd1 vccd1 vccd1 _09241_/D sky130_fd_sc_hd__buf_2
XFILLER_68_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09712_ _09712_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09712_/X sky130_fd_sc_hd__or2_1
XFILLER_68_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06924_ _14287_/Q _06873_/X _06923_/X _14383_/Q vssd1 vssd1 vccd1 vccd1 _06924_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09643_ _09641_/Y _09404_/X _09631_/Y _09642_/X vssd1 vssd1 vccd1 vccd1 _09651_/A
+ sky130_fd_sc_hd__o211a_1
X_06855_ _13782_/Q vssd1 vssd1 vccd1 vccd1 _06855_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _09573_/B _09573_/C _09573_/A vssd1 vssd1 vccd1 vccd1 _09574_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09233__B _09233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08525_ _08796_/A vssd1 vssd1 vccd1 vccd1 _09241_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13650__A0 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08657__B1 _08656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08456_ _08980_/A _08767_/B vssd1 vssd1 vccd1 vccd1 _08470_/A sky130_fd_sc_hd__nand2_1
X_07407_ _14092_/Q _07404_/X _07406_/X _13892_/Q _07521_/B vssd1 vssd1 vccd1 vccd1
+ _07407_/X sky130_fd_sc_hd__a221o_1
XANTENNA__13402__A0 _12610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08387_ _09683_/A _08387_/B _08387_/C vssd1 vssd1 vccd1 vccd1 _08388_/B sky130_fd_sc_hd__and3_1
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07338_ _14227_/Q vssd1 vssd1 vccd1 vccd1 _07482_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_104_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07269_ _14174_/Q _14173_/Q _14172_/Q _14171_/Q vssd1 vssd1 vccd1 vccd1 _07534_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_118_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ _09007_/B _09007_/C _09007_/A vssd1 vssd1 vccd1 vccd1 _09009_/B sky130_fd_sc_hd__a21oi_1
XFILLER_3_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10280_ _10281_/B _10280_/B vssd1 vssd1 vccd1 vccd1 _10282_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10519__A1 _07924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12115__A _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09127__C _09127_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11954__A _11971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13970_ _13988_/CLK _13970_/D _12395_/Y vssd1 vssd1 vccd1 vccd1 _13970_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_76_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12921_ _14155_/Q _12915_/X _12919_/X _12920_/X vssd1 vssd1 vccd1 vccd1 _14155_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12692__A1 _14056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12852_/A vssd1 vssd1 vccd1 vccd1 _14131_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _13785_/Q _11793_/X _11802_/X vssd1 vssd1 vccd1 vccd1 _11803_/X sky130_fd_sc_hd__a21o_2
XFILLER_55_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12801_/A vssd1 vssd1 vccd1 vccd1 _12783_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12444__A1 _14025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _13766_/Q _11714_/X _11716_/X _11733_/X vssd1 vssd1 vccd1 vccd1 _13766_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07320__B1 _07464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11665_ hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__inv_2
XFILLER_30_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14453_ _14453_/CLK _14453_/D vssd1 vssd1 vccd1 vccd1 _14453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_10_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_109_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13404_ _13404_/A vssd1 vssd1 vccd1 vccd1 _14368_/D sky130_fd_sc_hd__clkbuf_1
X_10616_ _10634_/A _10615_/Y _07924_/X vssd1 vssd1 vccd1 vccd1 _10616_/Y sky130_fd_sc_hd__a21oi_1
X_14384_ _14464_/CLK _14384_/D vssd1 vssd1 vccd1 vccd1 _14384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11596_ _11596_/A vssd1 vssd1 vccd1 vccd1 _13855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13335_ _14349_/Q _13332_/X _13334_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _14349_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10547_ _10547_/A vssd1 vssd1 vccd1 vccd1 _10565_/B sky130_fd_sc_hd__buf_2
X_13266_ _14446_/Q _13201_/X _13204_/X _14398_/Q vssd1 vssd1 vccd1 vccd1 _13266_/X
+ sky130_fd_sc_hd__a22o_1
X_10478_ _10478_/A vssd1 vssd1 vccd1 vccd1 _10503_/S sky130_fd_sc_hd__clkbuf_2
X_12217_ _12209_/X _12210_/X _12226_/B _12215_/X _12216_/X vssd1 vssd1 vccd1 vccd1
+ _13835_/D sky130_fd_sc_hd__o311a_1
X_13197_ _13197_/A _13197_/B vssd1 vssd1 vccd1 vccd1 _13526_/A sky130_fd_sc_hd__nor2_8
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12148_ input81/X _12160_/B vssd1 vssd1 vccd1 vccd1 _12148_/X sky130_fd_sc_hd__or2_1
XFILLER_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09128__A1 _09127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13555__S _13559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ _12079_/A vssd1 vssd1 vccd1 vccd1 _13804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08103__A2 _09233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ _09165_/C vssd1 vssd1 vccd1 vccd1 _09217_/D sky130_fd_sc_hd__clkbuf_2
X_09290_ _09284_/A _09284_/B _09284_/C vssd1 vssd1 vccd1 vccd1 _09291_/C sky130_fd_sc_hd__a21o_1
XFILLER_36_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08241_ _08239_/X _08193_/A _09749_/B _08240_/X vssd1 vssd1 vccd1 vccd1 _09749_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_60_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07939__D _09218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ _08084_/Y _08122_/X _08170_/Y _08171_/X vssd1 vssd1 vccd1 vccd1 _08194_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_119_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07123_ _07123_/A vssd1 vssd1 vccd1 vccd1 _14294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07054_ _07050_/X _14303_/Q _07054_/S vssd1 vssd1 vccd1 vccd1 _07055_/A sky130_fd_sc_hd__mux2_1
Xoutput110 _14069_/Q vssd1 vssd1 vccd1 vccd1 addr1[9] sky130_fd_sc_hd__buf_2
XFILLER_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput121 _11846_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[17] sky130_fd_sc_hd__buf_2
Xoutput132 _11863_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[27] sky130_fd_sc_hd__buf_2
Xoutput143 _11825_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[8] sky130_fd_sc_hd__buf_2
Xoutput154 _14310_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[18] sky130_fd_sc_hd__buf_2
Xoutput165 _14320_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[28] sky130_fd_sc_hd__buf_2
XANTENNA__11174__A1 _11032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput176 _14323_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[9] sky130_fd_sc_hd__buf_2
XFILLER_87_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07956_ _09803_/A vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__buf_2
XFILLER_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06907_ _14438_/Q _14262_/Q vssd1 vssd1 vccd1 vccd1 _06907_/Y sky130_fd_sc_hd__nand2_1
X_07887_ _07886_/A _07848_/A _07848_/B _07874_/S vssd1 vssd1 vccd1 vccd1 _07887_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_29_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09626_ _09626_/A _09626_/B _09626_/C vssd1 vssd1 vccd1 vccd1 _09626_/X sky130_fd_sc_hd__and3_1
XFILLER_16_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09557_ _09475_/B _09475_/C _09475_/A vssd1 vssd1 vccd1 vccd1 _09558_/C sky130_fd_sc_hd__a21bo_1
X_08508_ _09869_/B vssd1 vssd1 vccd1 vccd1 _09361_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_52_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09488_ _09488_/A _09488_/B _09488_/C vssd1 vssd1 vccd1 vccd1 _09540_/A sky130_fd_sc_hd__nand3_2
XFILLER_52_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08439_ _09863_/A vssd1 vssd1 vccd1 vccd1 _08794_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_1_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_8_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11450_ _11142_/B _11087_/B _13945_/Q vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__mux2_1
X_10401_ _10388_/A _10388_/B _10400_/X vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__o21a_2
X_11381_ hold13/X _11390_/B vssd1 vssd1 vccd1 vccd1 _11381_/X sky130_fd_sc_hd__or2_1
X_13120_ _13121_/A vssd1 vssd1 vccd1 vccd1 _13120_/Y sky130_fd_sc_hd__inv_2
X_10332_ _10332_/A _10332_/B vssd1 vssd1 vccd1 vccd1 _10349_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_clkbuf_leaf_76_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_106_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ input33/X input44/X _11988_/A _13037_/A vssd1 vssd1 vccd1 vccd1 _13051_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_11_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _10262_/X _10260_/A _10255_/B vssd1 vssd1 vccd1 vccd1 _10263_/Y sky130_fd_sc_hd__a21oi_1
X_12002_ _12060_/A vssd1 vssd1 vccd1 vccd1 _12021_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_3_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10194_ _10194_/A _10200_/A vssd1 vssd1 vccd1 vccd1 _10195_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input47_A io_wbs_adr[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13953_ _14020_/CLK _13953_/D _12374_/Y vssd1 vssd1 vccd1 vccd1 _13953_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_98_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _12904_/A _12913_/B vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__or2_1
XFILLER_98_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13884_ _14198_/CLK _13884_/D _12288_/Y vssd1 vssd1 vccd1 vccd1 _13884_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _12847_/A _12835_/B vssd1 vssd1 vccd1 vccd1 _12836_/A sky130_fd_sc_hd__and2_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _14149_/Q _12801_/A _12776_/A _14133_/Q _12765_/X vssd1 vssd1 vccd1 vccd1
+ _12766_/X sky130_fd_sc_hd__a221o_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07402__A _07528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ _13830_/Q vssd1 vssd1 vccd1 vccd1 _11717_/Y sky130_fd_sc_hd__inv_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _12697_/A vssd1 vssd1 vccd1 vccd1 _14057_/D sky130_fd_sc_hd__clkbuf_1
X_14436_ _14440_/CLK _14436_/D vssd1 vssd1 vccd1 vccd1 _14436_/Q sky130_fd_sc_hd__dfxtp_1
X_11648_ hold22/A _11647_/X _11652_/S vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 dout1[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 dout1[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 io_wbs_adr[10] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 io_wbs_adr[20] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
X_14367_ _14367_/CLK _14367_/D vssd1 vssd1 vccd1 vccd1 _14367_/Q sky130_fd_sc_hd__dfxtp_1
X_11579_ _11539_/Y _11598_/A _11597_/B vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__o21ai_2
Xinput56 io_wbs_adr[30] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
Xinput67 io_wbs_datwr[10] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
XFILLER_115_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput78 io_wbs_datwr[20] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__07548__S _07548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13318_ _14345_/Q _13311_/X _13317_/X _13301_/X vssd1 vssd1 vccd1 vccd1 _14345_/D
+ sky130_fd_sc_hd__o211a_1
Xinput89 io_wbs_datwr[30] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_2
X_14298_ _14410_/CLK _14298_/D _13164_/Y vssd1 vssd1 vccd1 vccd1 _14298_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_66_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08233__A _08403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13249_ _14330_/Q _13240_/X _13248_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _14330_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11156__A1 _10722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__B2 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07810_ _11452_/A _10664_/B _11452_/B vssd1 vssd1 vccd1 vccd1 _07810_/Y sky130_fd_sc_hd__a21oi_1
X_08790_ _09457_/B _09145_/D _13859_/Q _09457_/A vssd1 vssd1 vccd1 vccd1 _08821_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07741_ _07740_/Y _14156_/Q _07757_/S vssd1 vssd1 vccd1 vccd1 _07741_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07672_ _07672_/A _07672_/B vssd1 vssd1 vccd1 vccd1 _07673_/B sky130_fd_sc_hd__xor2_2
XFILLER_38_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09999__A _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09411_ _09411_/A _09411_/B _09411_/C vssd1 vssd1 vccd1 vccd1 _09411_/X sky130_fd_sc_hd__and3_1
XFILLER_80_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11533__S _11533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _09274_/B _09274_/Y _09337_/Y _09338_/X vssd1 vssd1 vccd1 vccd1 _09342_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_34_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13033__B _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ _09273_/A _09273_/B vssd1 vssd1 vccd1 vccd1 _10627_/B sky130_fd_sc_hd__and2_1
X_08224_ _08224_/A _08224_/B vssd1 vssd1 vccd1 vccd1 _08225_/B sky130_fd_sc_hd__nor2_1
XFILLER_14_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08155_ _08201_/A _08156_/B vssd1 vssd1 vccd1 vccd1 _08223_/C sky130_fd_sc_hd__or2_1
XFILLER_88_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07106_ _14408_/Q _07134_/B _14440_/Q vssd1 vssd1 vccd1 vccd1 _07106_/X sky130_fd_sc_hd__and3b_1
X_08086_ _14010_/Q vssd1 vssd1 vccd1 vccd1 _08796_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_106_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07037_ _07034_/X _14305_/Q _07037_/S vssd1 vssd1 vccd1 vccd1 _07038_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12895__A1 _14146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09760__A1 _09777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08988_ _08654_/A _08654_/C _08654_/B vssd1 vssd1 vccd1 vccd1 _08989_/C sky130_fd_sc_hd__o21bai_2
XFILLER_60_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07939_ _09084_/A _09084_/B _09233_/D _09218_/B vssd1 vssd1 vccd1 vccd1 _08004_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_28_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10950_ _10938_/X _10926_/X _10950_/S vssd1 vssd1 vccd1 vccd1 _10951_/B sky130_fd_sc_hd__mux2_2
XFILLER_44_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09609_ _09586_/B _09586_/Y _09675_/A _09608_/Y vssd1 vssd1 vccd1 vccd1 _09612_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_16_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10881_ _10906_/A _10873_/C _10879_/X _10880_/Y vssd1 vssd1 vccd1 vccd1 _10881_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12620_ _12620_/A vssd1 vssd1 vccd1 vccd1 _14038_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12551_ _12551_/A _12551_/B vssd1 vssd1 vccd1 vccd1 _12552_/A sky130_fd_sc_hd__and2_1
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11502_ _11502_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11502_/X sky130_fd_sc_hd__or2_1
XFILLER_32_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10830__B1 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12482_ _08317_/A _12465_/X _12476_/X _14050_/Q vssd1 vssd1 vccd1 vccd1 _12482_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11433_ _11436_/S vssd1 vssd1 vccd1 vccd1 _11446_/S sky130_fd_sc_hd__buf_2
XFILLER_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14221_ _14284_/CLK _14221_/D _13018_/Y vssd1 vssd1 vccd1 vccd1 _14221_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10189__A2 _10191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12583__A0 _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14152_ _14152_/CLK _14152_/D vssd1 vssd1 vccd1 vccd1 _14152_/Q sky130_fd_sc_hd__dfxtp_1
X_11364_ _13857_/Q vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__inv_2
XANTENNA__10594__C1 _09788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13103_ _13106_/A _13103_/B vssd1 vssd1 vccd1 vccd1 _13104_/A sky130_fd_sc_hd__and2_1
X_10315_ _10292_/B _10315_/B vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__and2b_1
X_14083_ _14217_/CLK _14083_/D _12730_/Y vssd1 vssd1 vccd1 vccd1 _14083_/Q sky130_fd_sc_hd__dfrtp_2
X_11295_ _11320_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11324_/A sky130_fd_sc_hd__or2_1
XFILLER_112_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13034_ hold27/A _11988_/A _13035_/A _13033_/Y _14240_/Q vssd1 vssd1 vccd1 vccd1
+ _13034_/X sky130_fd_sc_hd__a32o_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10246_ _10116_/A _10116_/B _10245_/X vssd1 vssd1 vccd1 vccd1 _10250_/B sky130_fd_sc_hd__a21oi_2
XFILLER_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output153_A _14309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10177_ _10174_/A _10174_/B _10173_/A _10173_/B vssd1 vssd1 vccd1 vccd1 _10178_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12303__A _12304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13936_ _14102_/CLK _13936_/D _12352_/Y vssd1 vssd1 vccd1 vccd1 _13936_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11310__A1 _11087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11310__B2 _10826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13867_ _13867_/CLK _13867_/D _12267_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Q sky130_fd_sc_hd__dfrtp_4
X_12818_ _14121_/Q _12771_/X _12816_/X _12817_/X vssd1 vssd1 vccd1 vccd1 _14121_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13063__A1 _14241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ _14335_/CLK _13798_/D vssd1 vssd1 vccd1 vccd1 _13798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12810__A1 _14159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12752_/A vssd1 vssd1 vccd1 vccd1 _12749_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08490__B2 _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14419_ _14452_/CLK _14419_/D vssd1 vssd1 vccd1 vccd1 _14419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09960_ _09854_/A _09854_/B _09959_/Y vssd1 vssd1 vccd1 vccd1 _10269_/A sky130_fd_sc_hd__o21bai_2
XFILLER_98_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08911_ _08911_/A _08916_/A vssd1 vssd1 vccd1 vccd1 _08912_/B sky130_fd_sc_hd__and2_1
XFILLER_48_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09891_ _10092_/B vssd1 vssd1 vccd1 vccd1 _09893_/A sky130_fd_sc_hd__clkinv_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08842_/A _10171_/A vssd1 vssd1 vccd1 vccd1 _08844_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08735_/A _08735_/B _08735_/C vssd1 vssd1 vccd1 vccd1 _08776_/B sky130_fd_sc_hd__a21oi_1
X_07724_ _07765_/S vssd1 vssd1 vccd1 vccd1 _07724_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07655_ _14073_/Q _07716_/A vssd1 vssd1 vccd1 vccd1 _07656_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09241__B _09241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07586_ _07586_/A vssd1 vssd1 vccd1 vccd1 _14090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_30_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13897_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09325_ _09346_/B _09324_/C _09324_/B vssd1 vssd1 vccd1 vccd1 _09325_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_90_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07808__A1 _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12883__A _12926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ _09254_/Y _09253_/X _09180_/Y _09180_/C vssd1 vssd1 vccd1 vccd1 _09274_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__07977__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08207_ _09762_/B _09999_/A vssd1 vssd1 vccd1 vccd1 _08212_/A sky130_fd_sc_hd__nand2_2
X_09187_ _09187_/A vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12565__B1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ _08621_/A _10000_/B _08213_/A _08134_/Y vssd1 vssd1 vccd1 vccd1 _08203_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08784__A2 _08937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08069_ _08128_/A vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__clkbuf_4
X_10100_ _10100_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10143_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10591__A2 _09663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11080_ _11097_/B _11080_/B vssd1 vssd1 vccd1 vccd1 _11080_/X sky130_fd_sc_hd__and2_1
XFILLER_103_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10031_ _10421_/B _10252_/B _10030_/B _10030_/A vssd1 vssd1 vccd1 vccd1 _10032_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12123__A _12940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13653__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13293__A1 _14339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11982_ _12933_/A vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__buf_2
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13721_ input82/X _14460_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13722_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10933_ _13906_/Q _13907_/Q _13908_/Q _13909_/Q _10931_/A _13948_/Q vssd1 vssd1 vccd1
+ vccd1 _10933_/X sky130_fd_sc_hd__mux4_2
XFILLER_83_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13652_ _13652_/A vssd1 vssd1 vccd1 vccd1 _14439_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10864_ _13978_/Q _10895_/B vssd1 vssd1 vccd1 vccd1 _10864_/X sky130_fd_sc_hd__and2_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _12611_/S vssd1 vssd1 vccd1 vccd1 _12621_/S sky130_fd_sc_hd__buf_2
X_13583_ input73/X _14420_/Q _13593_/S vssd1 vssd1 vccd1 vccd1 _13584_/B sky130_fd_sc_hd__mux2_1
X_10795_ _10879_/B _10795_/B vssd1 vssd1 vccd1 vccd1 _10884_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12534_ _12534_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _12535_/A sky130_fd_sc_hd__and2_1
XFILLER_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13348__A2 _13236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12465_ _12486_/A vssd1 vssd1 vccd1 vccd1 _12465_/X sky130_fd_sc_hd__clkbuf_2
X_14204_ _14211_/CLK _14204_/D _12996_/Y vssd1 vssd1 vccd1 vccd1 _14204_/Q sky130_fd_sc_hd__dfrtp_1
X_11416_ _11271_/A _11032_/A _11425_/S vssd1 vssd1 vccd1 vccd1 _11521_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12396_ _12397_/A vssd1 vssd1 vccd1 vccd1 _12396_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11347_ _11347_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11348_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08775__A2 _08767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14135_ _14152_/CLK _14135_/D vssd1 vssd1 vccd1 vccd1 _14135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ _11341_/B _11345_/A _11341_/A vssd1 vssd1 vccd1 vccd1 _11342_/A sky130_fd_sc_hd__a21oi_1
X_14066_ _14179_/CLK _14066_/D _12708_/Y vssd1 vssd1 vccd1 vccd1 _14066_/Q sky130_fd_sc_hd__dfrtp_1
X_10229_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10229_/X sky130_fd_sc_hd__or2_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13017_ _13116_/A vssd1 vssd1 vccd1 vccd1 _13022_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11531__A1 _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11531__B2 _13895_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__buf_2
XFILLER_95_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11872__A _11872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13919_ _13920_/CLK _13919_/D _12332_/Y vssd1 vssd1 vccd1 vccd1 _13919_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__14415__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07440_ _14086_/Q _07432_/X _07433_/X _13886_/Q _07417_/X vssd1 vssd1 vccd1 vccd1
+ _07440_/X sky130_fd_sc_hd__a221o_1
XANTENNA__13036__A1 _14241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11047__B1 _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07371_ _07349_/X _07369_/X _07370_/X _07352_/X vssd1 vssd1 vccd1 vccd1 _07371_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10000__B _10000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09110_ _09110_/A _09118_/A _09110_/C vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__and3_2
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09041_ _09041_/A _08974_/B vssd1 vssd1 vccd1 vccd1 _09041_/X sky130_fd_sc_hd__or2b_1
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12547__A0 _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11112__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ _10081_/A _09943_/B _10057_/A vssd1 vssd1 vccd1 vccd1 _10173_/B sky130_fd_sc_hd__and3_2
XFILLER_86_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13039__A _13254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _09903_/A vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__buf_4
XFILLER_98_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _08831_/A _08831_/C _08869_/A vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__a21o_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12878__A _12922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08756_ _08756_/A _08756_/B vssd1 vssd1 vccd1 vccd1 _08757_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06876__A _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10089__A1 _10127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14095__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _14148_/Q _07651_/X _07702_/X _14256_/Q vssd1 vssd1 vccd1 vccd1 _07764_/S
+ sky130_fd_sc_hd__o211ai_4
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__A2 _11808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ _08687_/A _08687_/B _08687_/C vssd1 vssd1 vccd1 vccd1 _08688_/B sky130_fd_sc_hd__and3_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _14130_/Q _14065_/Q vssd1 vssd1 vccd1 vccd1 _07671_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07569_ _14097_/Q input14/X _07571_/S vssd1 vssd1 vccd1 vccd1 _07570_/A sky130_fd_sc_hd__mux2_1
XFILLER_110_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09308_ _09393_/A _09393_/C _09393_/B vssd1 vssd1 vccd1 vccd1 _09308_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ _13961_/Q _10579_/Y _10585_/S vssd1 vssd1 vccd1 vccd1 _10581_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09239_ _09239_/A _09239_/B _09239_/C vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__nand3_2
XFILLER_103_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_15_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11022__A _11058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12250_ _12251_/A vssd1 vssd1 vccd1 vccd1 _12250_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11201_ _11216_/B _11217_/A _11213_/A vssd1 vssd1 vccd1 vccd1 _11207_/B sky130_fd_sc_hd__nor3_1
XFILLER_119_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12181_ _12181_/A vssd1 vssd1 vccd1 vccd1 _13042_/A sky130_fd_sc_hd__inv_2
XFILLER_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11132_ _11135_/A _11132_/B vssd1 vssd1 vccd1 vccd1 _11132_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11063_ _11117_/B _11117_/C _11062_/X vssd1 vssd1 vccd1 vccd1 _11114_/C sky130_fd_sc_hd__a21bo_1
XFILLER_62_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09146__B _09870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10014_ _10397_/B _10011_/A vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__or2b_1
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14438__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11965_ _11965_/A vssd1 vssd1 vccd1 vccd1 _11965_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output116_A _11836_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13704_ input76/X _14455_/Q _13704_/S vssd1 vssd1 vccd1 vccd1 _13705_/B sky130_fd_sc_hd__mux2_1
X_10916_ _10916_/A _11087_/B vssd1 vssd1 vccd1 vccd1 _10916_/X sky130_fd_sc_hd__or2_1
XFILLER_17_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11896_ _13754_/Q _11897_/B vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__and2_1
X_13635_ _13644_/A _13635_/B vssd1 vssd1 vccd1 vccd1 _13636_/A sky130_fd_sc_hd__and2_1
XFILLER_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07113__C _14439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10847_ _10900_/B vssd1 vssd1 vccd1 vccd1 _10906_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13412__A _13447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13566_ _12673_/X _14415_/Q _13576_/S vssd1 vssd1 vccd1 vccd1 _13567_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08506__A _09349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10778_ _10713_/A _10755_/Y _10777_/X _10770_/A vssd1 vssd1 vccd1 vccd1 _10783_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07410__A _07464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12517_ _12517_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__and2_1
X_13497_ _13497_/A vssd1 vssd1 vccd1 vccd1 _13511_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12028__A _12216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12448_ _13991_/Q _12422_/X _12447_/X _12203_/X vssd1 vssd1 vccd1 vccd1 _13991_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ _12379_/A vssd1 vssd1 vccd1 vccd1 _12384_/A sky130_fd_sc_hd__buf_2
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14118_ _14163_/CLK _14118_/D vssd1 vssd1 vccd1 vccd1 _14118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06940_ _14429_/Q _06939_/Y _06931_/X vssd1 vssd1 vccd1 vccd1 _06940_/X sky130_fd_sc_hd__a21o_1
X_14049_ _14411_/CLK _14049_/D vssd1 vssd1 vccd1 vccd1 _14049_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11504__A1 _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06871_ _07105_/A vssd1 vssd1 vccd1 vccd1 _07027_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12698__A _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ _08682_/A _08610_/B vssd1 vssd1 vccd1 vccd1 _08620_/A sky130_fd_sc_hd__xor2_2
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09590_ _09590_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09670_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08541_ _08547_/D vssd1 vssd1 vccd1 vccd1 _08783_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08472_ _09378_/B vssd1 vssd1 vccd1 vccd1 _09217_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07423_ _14089_/Q _07404_/X _07406_/X hold39/X _07417_/X vssd1 vssd1 vccd1 vccd1
+ _07423_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09800__A _09800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12217__C1 _12216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_io_wbs_clk_A clkbuf_3_7_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__13322__A _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07354_ _14219_/Q _07347_/X _07348_/X _07353_/X vssd1 vssd1 vccd1 vccd1 _14219_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08416__A _09188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_109_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07285_ _14243_/Q _14231_/Q _07519_/A vssd1 vssd1 vccd1 vccd1 _07286_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06998__A1 _14310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ _09023_/B _09023_/C _09023_/A vssd1 vssd1 vccd1 vccd1 _09025_/D sky130_fd_sc_hd__a21o_1
XANTENNA__11991__A1 _13823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11777__A _13206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11743__A1 _13823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09926_ _09926_/A _09926_/B vssd1 vssd1 vccd1 vccd1 _10331_/A sky130_fd_sc_hd__or2_4
XFILLER_113_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07990__A _09821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _09857_/A _09857_/B vssd1 vssd1 vccd1 vccd1 _10091_/A sky130_fd_sc_hd__xnor2_4
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _08757_/A _08756_/A _08756_/B vssd1 vssd1 vccd1 vccd1 _08809_/B sky130_fd_sc_hd__o21ba_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09788_ _09788_/A vssd1 vssd1 vccd1 vccd1 _09788_/X sky130_fd_sc_hd__buf_2
XFILLER_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _08740_/A _08740_/B vssd1 vssd1 vccd1 vccd1 _08779_/B sky130_fd_sc_hd__xnor2_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11749_/Y hold16/A _07548_/S vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__o21bai_1
XFILLER_54_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _11110_/A vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12208__C1 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11681_/A vssd1 vssd1 vccd1 vccd1 _13778_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13420_ _13426_/A _13420_/B vssd1 vssd1 vccd1 vccd1 _13421_/A sky130_fd_sc_hd__and2_1
X_10632_ _10632_/A _10632_/B vssd1 vssd1 vccd1 vccd1 _10633_/B sky130_fd_sc_hd__nor2_1
X_13351_ _14386_/Q _13236_/A _13336_/X _14466_/Q vssd1 vssd1 vccd1 vccd1 _13351_/X
+ sky130_fd_sc_hd__a22o_1
X_10563_ _07924_/X _10556_/Y _10561_/Y _10562_/X vssd1 vssd1 vccd1 vccd1 _13963_/D
+ sky130_fd_sc_hd__o31a_1
X_12302_ _12304_/A vssd1 vssd1 vccd1 vccd1 _12302_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input77_A io_wbs_datwr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13282_ _14369_/Q _13208_/X _13281_/X _13258_/X vssd1 vssd1 vccd1 vccd1 _13282_/X
+ sky130_fd_sc_hd__a211o_1
X_10494_ _10495_/A _10495_/B vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12233_ _12233_/A vssd1 vssd1 vccd1 vccd1 _12233_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ _12913_/A _12173_/B vssd1 vssd1 vccd1 vccd1 _12164_/X sky130_fd_sc_hd__or2_1
XFILLER_29_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11115_ _11125_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11115_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12095_ _12095_/A vssd1 vssd1 vccd1 vccd1 _12095_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13828__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11046_ _13912_/Q vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__buf_2
XANTENNA__11498__B1 _10686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12311__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06913__A1 _14321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12997_ _12997_/A vssd1 vssd1 vccd1 vccd1 _12997_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07124__B _14289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ _11971_/A vssd1 vssd1 vccd1 vccd1 _11953_/A sky130_fd_sc_hd__buf_2
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11879_ _13748_/Q _13747_/Q _13749_/Q vssd1 vssd1 vccd1 vccd1 _11879_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13142__A _13146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13618_ input84/X _14430_/Q _13628_/S vssd1 vssd1 vccd1 vccd1 _13619_/B sky130_fd_sc_hd__mux2_1
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07140__A _07185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13549_ input94/X _14410_/Q _13559_/S vssd1 vssd1 vccd1 vccd1 _13550_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07070_ _07070_/A vssd1 vssd1 vccd1 vccd1 _14301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07972_ _13873_/Q vssd1 vssd1 vccd1 vccd1 _09457_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_09711_ _09708_/B _09708_/Y _09692_/Y _09709_/X vssd1 vssd1 vccd1 vccd1 _09715_/A
+ sky130_fd_sc_hd__a211oi_1
X_06923_ _14431_/Q _06922_/Y _06877_/X vssd1 vssd1 vccd1 vccd1 _06923_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09642_ _09631_/A _09631_/C _09631_/B vssd1 vssd1 vccd1 vccd1 _09642_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12221__A _12517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__A1 _06894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07315__A _07452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09573_ _09573_/A _09573_/B _09573_/C vssd1 vssd1 vccd1 vccd1 _09573_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__09233__C _09233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _08978_/B _10007_/A _09000_/B _08978_/A vssd1 vssd1 vccd1 vccd1 _08529_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13650__A1 _14439_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09530__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10464__A1 _10302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ _09434_/B vssd1 vssd1 vccd1 vccd1 _08767_/B sky130_fd_sc_hd__buf_6
X_07406_ _07460_/A vssd1 vssd1 vccd1 vccd1 _07406_/X sky130_fd_sc_hd__clkbuf_2
X_08386_ _08387_/B _08387_/C _08298_/A vssd1 vssd1 vccd1 vccd1 _08388_/A sky130_fd_sc_hd__a21oi_1
XFILLER_23_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08146__A _08146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07337_ _14104_/Q _07336_/X vssd1 vssd1 vccd1 vccd1 _07337_/X sky130_fd_sc_hd__or2b_1
XFILLER_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12891__A _12936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07268_ _07264_/Y _07266_/Y _07267_/X vssd1 vssd1 vccd1 vccd1 _07280_/A sky130_fd_sc_hd__a21oi_2
XFILLER_87_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09007_ _09007_/A _09007_/B _09007_/C vssd1 vssd1 vccd1 vccd1 _09009_/A sky130_fd_sc_hd__and3_1
XFILLER_118_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07199_ _07199_/A vssd1 vssd1 vccd1 vccd1 _14278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09909_ _09903_/Y _10171_/B _10153_/B vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__a21oi_2
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12920_ _12920_/A vssd1 vssd1 vccd1 vccd1 _12920_/X sky130_fd_sc_hd__buf_2
XFILLER_111_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12131__A _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12851_ _13070_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12852_/A sky130_fd_sc_hd__and2_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _14326_/Q _11870_/B _11797_/X _13991_/Q _11801_/X vssd1 vssd1 vccd1 vccd1
+ _11802_/X sky130_fd_sc_hd__a221o_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12800_/A vssd1 vssd1 vccd1 vccd1 _12782_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11729_/B _11732_/Y _11718_/X _13826_/Q vssd1 vssd1 vccd1 vccd1 _11733_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14452_/CLK _14452_/D vssd1 vssd1 vccd1 vccd1 _14452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _13781_/Q _11669_/A _11661_/X _11686_/A vssd1 vssd1 vccd1 vccd1 _11664_/Y
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__08056__A _13872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13403_ _13409_/A _13403_/B vssd1 vssd1 vccd1 vccd1 _13404_/A sky130_fd_sc_hd__and2_1
X_10615_ _10615_/A _10615_/B vssd1 vssd1 vccd1 vccd1 _10615_/Y sky130_fd_sc_hd__xnor2_1
X_14383_ _14464_/CLK _14383_/D vssd1 vssd1 vccd1 vccd1 _14383_/Q sky130_fd_sc_hd__dfxtp_1
X_11595_ _13855_/Q _11592_/Y _11611_/S vssd1 vssd1 vccd1 vccd1 _11596_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13334_ _14429_/Q _13327_/X _13333_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13334_/X
+ sky130_fd_sc_hd__a211o_1
X_10546_ _10546_/A _10546_/B _10546_/C vssd1 vssd1 vccd1 vccd1 _10546_/X sky130_fd_sc_hd__and3_1
XFILLER_10_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13265_ _13265_/A vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10477_ _10485_/A _10477_/B vssd1 vssd1 vccd1 vccd1 _10480_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12216_ _12216_/A vssd1 vssd1 vccd1 vccd1 _12216_/X sky130_fd_sc_hd__buf_2
X_13196_ _13265_/A vssd1 vssd1 vccd1 vccd1 _13196_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12147_ _12147_/A vssd1 vssd1 vccd1 vccd1 _12160_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09128__A2 _09127_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ _12081_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12079_/A sky130_fd_sc_hd__and2_1
XFILLER_81_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11029_ _11029_/A _11029_/B vssd1 vssd1 vccd1 vccd1 _11054_/B sky130_fd_sc_hd__xnor2_1
XFILLER_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09053__C _09824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08240_ _08274_/B _08235_/X _08173_/Y _08194_/X vssd1 vssd1 vccd1 vccd1 _08240_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13396__A0 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _08170_/A _08170_/B _08170_/C vssd1 vssd1 vccd1 vccd1 _08171_/X sky130_fd_sc_hd__o21a_1
X_07122_ _07119_/X _14294_/Q _07122_/S vssd1 vssd1 vccd1 vccd1 _07123_/A sky130_fd_sc_hd__mux2_1
XANTENNA__07075__B1 _14364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07053_ _07051_/X _07052_/X _14367_/Q vssd1 vssd1 vccd1 vccd1 _07054_/S sky130_fd_sc_hd__o21a_1
XFILLER_118_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12216__A _12216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput111 _11745_/Y vssd1 vssd1 vccd1 vccd1 csb1 sky130_fd_sc_hd__buf_2
Xoutput122 _11849_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[18] sky130_fd_sc_hd__buf_2
Xoutput133 _11865_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[28] sky130_fd_sc_hd__buf_2
XFILLER_47_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput144 _11827_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[9] sky130_fd_sc_hd__buf_2
Xoutput155 _14292_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[19] sky130_fd_sc_hd__buf_2
XFILLER_82_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput166 _14293_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[29] sky130_fd_sc_hd__buf_2
Xoutput177 _14168_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_spi_cs_no sky130_fd_sc_hd__buf_2
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11774__B _11774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _13869_/Q vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__buf_2
X_06906_ _06906_/A vssd1 vssd1 vccd1 vccd1 _14322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07886_ _07886_/A _07886_/B vssd1 vssd1 vccd1 vccd1 _07886_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ _09396_/C _09396_/Y _09470_/X _09624_/X vssd1 vssd1 vccd1 vccd1 _09631_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09556_ _09555_/A _09555_/B _09555_/C vssd1 vssd1 vccd1 vccd1 _09558_/B sky130_fd_sc_hd__a21o_1
XFILLER_52_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08507_ _08750_/B vssd1 vssd1 vccd1 vccd1 _08823_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09487_ _09437_/B _09437_/C _09437_/A vssd1 vssd1 vccd1 vccd1 _09488_/C sky130_fd_sc_hd__a21bo_1
XFILLER_12_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08438_ _09207_/C vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11014__B _11014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ _08579_/A _13874_/Q _09457_/D _09165_/A vssd1 vssd1 vccd1 vccd1 _09595_/B
+ sky130_fd_sc_hd__a22o_1
X_10400_ _10400_/A _10386_/A vssd1 vssd1 vccd1 vccd1 _10400_/X sky130_fd_sc_hd__or2b_1
X_11380_ _11407_/B vssd1 vssd1 vccd1 vccd1 _11390_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ _10331_/A _10423_/A vssd1 vssd1 vccd1 vccd1 _10332_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12126__A _12942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11030__A _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13050_ _14236_/Q _13041_/X _13049_/X _13039_/X vssd1 vssd1 vccd1 vccd1 _14236_/D
+ sky130_fd_sc_hd__o211a_1
X_10262_ _10254_/A _10254_/B _10254_/C vssd1 vssd1 vccd1 vccd1 _10262_/X sky130_fd_sc_hd__a21o_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12001_ _12059_/A _12001_/B vssd1 vssd1 vccd1 vccd1 _12060_/A sky130_fd_sc_hd__nor2_2
X_10193_ _10199_/A _10199_/B vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__nor2_1
XFILLER_94_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13952_ _14020_/CLK _13952_/D _12372_/Y vssd1 vssd1 vccd1 vccd1 _13952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12903_ _12942_/B vssd1 vssd1 vccd1 vccd1 _12913_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13883_ _14198_/CLK _13883_/D _12287_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12834_ _12515_/X _14126_/Q _12846_/S vssd1 vssd1 vccd1 vccd1 _12835_/B sky130_fd_sc_hd__mux2_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _14125_/Q _13200_/B _12761_/X vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__a21bo_1
XFILLER_43_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11716_/A vssd1 vssd1 vccd1 vccd1 _11716_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A _12696_/B vssd1 vssd1 vccd1 vccd1 _12697_/A sky130_fd_sc_hd__and2_1
XFILLER_30_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14435_ _14467_/CLK _14435_/D vssd1 vssd1 vccd1 vccd1 _14435_/Q sky130_fd_sc_hd__dfxtp_1
X_11647_ _11647_/A _11647_/B vssd1 vssd1 vccd1 vccd1 _11647_/X sky130_fd_sc_hd__xor2_1
Xinput13 dout1[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
Xinput24 dout1[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_2
XANTENNA__07057__B1 _07048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput35 io_wbs_adr[11] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
X_14366_ _14417_/CLK _14366_/D vssd1 vssd1 vccd1 vccd1 _14366_/Q sky130_fd_sc_hd__dfxtp_1
Xinput46 io_wbs_adr[21] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
X_11578_ _14054_/Q _13966_/Q vssd1 vssd1 vccd1 vccd1 _11597_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput57 io_wbs_adr[31] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
X_14474__186 vssd1 vssd1 vccd1 vccd1 _14474__186/HI io_oeb[6] sky130_fd_sc_hd__conb_1
Xinput68 io_wbs_datwr[11] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
X_13317_ _14425_/Q _13306_/X _13316_/X _13299_/X vssd1 vssd1 vccd1 vccd1 _13317_/X
+ sky130_fd_sc_hd__a211o_1
Xinput79 io_wbs_datwr[21] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__clkbuf_4
X_10529_ _09725_/X _09741_/X _09745_/X _09741_/B vssd1 vssd1 vccd1 vccd1 _10530_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14297_ _14410_/CLK _14297_/D _13163_/Y vssd1 vssd1 vccd1 vccd1 _14297_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13248_ _14362_/Q _13215_/X _13247_/X _13222_/X vssd1 vssd1 vccd1 vccd1 _13248_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13179_ _13183_/A vssd1 vssd1 vccd1 vccd1 _13179_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07740_ _07740_/A vssd1 vssd1 vccd1 vccd1 _07740_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_96_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07671_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09999__B _09999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07532__B2 _07528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ _09411_/A _09411_/C _09411_/B vssd1 vssd1 vccd1 vccd1 _09410_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_37_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14104_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09341_ _09635_/A _09341_/B vssd1 vssd1 vccd1 vccd1 _09341_/X sky130_fd_sc_hd__or2_1
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11115__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _09271_/A _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09273_/B sky130_fd_sc_hd__o21ai_4
X_08223_ _08298_/A _08223_/B _08223_/C vssd1 vssd1 vccd1 vccd1 _08224_/B sky130_fd_sc_hd__and3_1
XFILLER_20_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08154_ _08223_/B _08154_/B vssd1 vssd1 vccd1 vccd1 _08156_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07105_ _07105_/A vssd1 vssd1 vccd1 vccd1 _07134_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_49_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08085_ _08160_/C _08082_/Y _08325_/A _08052_/Y vssd1 vssd1 vccd1 vccd1 _08122_/B
+ sky130_fd_sc_hd__o211a_1
X_07036_ _07012_/X _07035_/X _14369_/Q vssd1 vssd1 vccd1 vccd1 _07037_/S sky130_fd_sc_hd__o21a_1
XFILLER_115_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08987_ _08986_/B _08986_/C _08986_/A vssd1 vssd1 vccd1 vccd1 _08989_/B sky130_fd_sc_hd__a21o_1
XFILLER_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07938_ _09817_/B vssd1 vssd1 vccd1 vccd1 _09218_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_95_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07869_ _07869_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07869_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_29_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09608_ _09607_/B _09607_/C _09607_/A vssd1 vssd1 vccd1 vccd1 _09608_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10880_ _13975_/Q _10895_/B vssd1 vssd1 vccd1 vccd1 _10880_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09539_ _09582_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__xnor2_1
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12550_ _12932_/A _08128_/B _12555_/S vssd1 vssd1 vccd1 vccd1 _12551_/B sky130_fd_sc_hd__mux2_1
XFILLER_19_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11501_ _08836_/B _11486_/X _11498_/Y _11500_/X vssd1 vssd1 vccd1 vccd1 _13867_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10830__A1 _10669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12481_ _12481_/A vssd1 vssd1 vccd1 vccd1 _12481_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13240__A _13265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14220_ _14284_/CLK _14220_/D _13016_/Y vssd1 vssd1 vccd1 vccd1 _14220_/Q sky130_fd_sc_hd__dfrtp_1
X_11432_ _11493_/A _11493_/B vssd1 vssd1 vccd1 vccd1 _11487_/A sky130_fd_sc_hd__nand2_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08334__A _09336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12583__A1 _14028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ _14158_/CLK _14151_/D vssd1 vssd1 vccd1 vccd1 _14151_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11363_ _11392_/A vssd1 vssd1 vccd1 vccd1 _11363_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13102_ _12650_/X hold29/A _13105_/S vssd1 vssd1 vccd1 vccd1 _13103_/B sky130_fd_sc_hd__mux2_1
X_10314_ _10314_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10366_/A sky130_fd_sc_hd__xnor2_1
X_14082_ _14217_/CLK _14082_/D _12727_/Y vssd1 vssd1 vccd1 vccd1 _14082_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11294_ _11294_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11295_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13532__A0 _13084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13033_ _13035_/A _13359_/A vssd1 vssd1 vccd1 vccd1 _13033_/Y sky130_fd_sc_hd__nand2_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10245_ _10115_/B _10245_/B vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__and2b_1
XFILLER_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10176_ _10176_/A _10176_/B vssd1 vssd1 vccd1 vccd1 _10180_/B sky130_fd_sc_hd__xnor2_2
XFILLER_79_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output146_A _14302_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_2_0_io_wbs_clk_A clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_75_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_22_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__11846__B1 _11848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13935_ _14102_/CLK _13935_/D _12351_/Y vssd1 vssd1 vccd1 vccd1 _13935_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11310__A2 _10845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13866_ _13867_/CLK _13866_/D _12266_/Y vssd1 vssd1 vccd1 vccd1 _13866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12817_ _12817_/A vssd1 vssd1 vccd1 vccd1 _12817_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13797_ _14335_/CLK _13797_/D vssd1 vssd1 vccd1 vccd1 _13797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12752_/A vssd1 vssd1 vccd1 vccd1 _12748_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12679_ _12679_/A vssd1 vssd1 vccd1 vccd1 _14052_/D sky130_fd_sc_hd__clkbuf_1
X_14418_ _14449_/CLK _14418_/D vssd1 vssd1 vccd1 vccd1 _14418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14349_ _14354_/CLK _14349_/D vssd1 vssd1 vccd1 vccd1 _14349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08910_ _08911_/A _08916_/A vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__nor2_1
XFILLER_48_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09890_ _09883_/Y _10157_/A _10129_/B vssd1 vssd1 vccd1 vccd1 _09894_/A sky130_fd_sc_hd__a21oi_4
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08841_ _10156_/A vssd1 vssd1 vccd1 vccd1 _10171_/A sky130_fd_sc_hd__buf_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08772_ _08772_/A _08772_/B vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07723_ _07723_/A vssd1 vssd1 vccd1 vccd1 _07723_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07654_ _14146_/Q vssd1 vssd1 vccd1 vccd1 _07700_/A sky130_fd_sc_hd__inv_2
XANTENNA__08419__A _09206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07323__A _07363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07585_ _14090_/Q input6/X _07593_/S vssd1 vssd1 vccd1 vccd1 _07586_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09324_ _09346_/B _09324_/B _09324_/C vssd1 vssd1 vccd1 vccd1 _09399_/A sky130_fd_sc_hd__and3_2
XFILLER_34_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07808__A2 _10705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09255_ _09180_/C _09180_/Y _09253_/X _09254_/Y vssd1 vssd1 vccd1 vccd1 _09258_/A
+ sky130_fd_sc_hd__a211o_1
X_08206_ _08621_/A vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__clkbuf_4
X_09186_ _09118_/Y _09110_/X _09184_/Y _09185_/X vssd1 vssd1 vccd1 vccd1 _09187_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12565__A1 _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08137_ _08213_/A _08134_/Y _08621_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _08213_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_88_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07993__A _08571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ _08124_/A _08124_/B vssd1 vssd1 vccd1 vccd1 _08125_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13514__A0 _12681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ _14275_/Q _07007_/X _07018_/X _14371_/Q vssd1 vssd1 vccd1 vccd1 _07019_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11915__A1_N _13820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12404__A _12410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10030_ _10030_/A _10030_/B vssd1 vssd1 vccd1 vccd1 _10252_/B sky130_fd_sc_hd__xor2_1
XFILLER_88_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ _12233_/A vssd1 vssd1 vccd1 vccd1 _11981_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13720_ _13720_/A vssd1 vssd1 vccd1 vccd1 _14459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10932_ _13898_/Q _13899_/Q _13900_/Q _13901_/Q _11169_/S _07798_/A vssd1 vssd1 vccd1
+ vccd1 _10932_/X sky130_fd_sc_hd__mux4_2
XFILLER_72_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ _13661_/A _13651_/B vssd1 vssd1 vccd1 vccd1 _13652_/A sky130_fd_sc_hd__and2_1
XFILLER_72_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10863_ _10863_/A _10863_/B _10869_/A vssd1 vssd1 vccd1 vccd1 _10863_/X sky130_fd_sc_hd__or3_1
XFILLER_13_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _12602_/A vssd1 vssd1 vccd1 vccd1 _14033_/D sky130_fd_sc_hd__clkbuf_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A vssd1 vssd1 vccd1 vccd1 _14419_/D sky130_fd_sc_hd__clkbuf_1
X_10794_ _10768_/B _10768_/A _13932_/Q vssd1 vssd1 vccd1 vccd1 _10795_/B sky130_fd_sc_hd__o21bai_1
XFILLER_40_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12533_ _12919_/A _08983_/A _12537_/S vssd1 vssd1 vccd1 vccd1 _12534_/B sky130_fd_sc_hd__mux2_1
XFILLER_40_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12464_ _12485_/A vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14203_ _14215_/CLK _14203_/D _12995_/Y vssd1 vssd1 vccd1 vccd1 _14203_/Q sky130_fd_sc_hd__dfrtp_1
X_11415_ _11415_/A vssd1 vssd1 vccd1 vccd1 _11425_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__10567__B1 _09788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ _12397_/A vssd1 vssd1 vccd1 vccd1 _12395_/Y sky130_fd_sc_hd__inv_2
XFILLER_67_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14134_ _14149_/CLK _14134_/D vssd1 vssd1 vccd1 vccd1 _14134_/Q sky130_fd_sc_hd__dfxtp_1
X_11346_ _11273_/A _10904_/X _11345_/X _07784_/X vssd1 vssd1 vccd1 vccd1 _13898_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13505__A0 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ _14065_/CLK _14065_/D _12707_/Y vssd1 vssd1 vccd1 vccd1 _14065_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10533__S _10585_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _11338_/A _11277_/B vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__or2_1
XFILLER_3_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13016_ _13016_/A vssd1 vssd1 vccd1 vccd1 _13016_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07408__A _07462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ _10232_/A _10232_/B vssd1 vssd1 vccd1 vccd1 _10228_/X sky130_fd_sc_hd__and2_1
XFILLER_95_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07127__B _07134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__xor2_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13145__A _13146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13918_ _13920_/CLK _13918_/D _12331_/Y vssd1 vssd1 vccd1 vccd1 _13918_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__08239__A _09777_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13849_ _13988_/CLK _13849_/D _12243_/Y vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfrtp_1
XFILLER_63_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07370_ _14214_/Q _14216_/Q _07387_/S vssd1 vssd1 vccd1 vccd1 _07370_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09040_ _08688_/A _08966_/X _09032_/X _09033_/Y vssd1 vssd1 vccd1 vccd1 _09040_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_50_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13744__A0 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__A1 _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__A _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11070__A_N _11007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09942_ _09942_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__xor2_4
XANTENNA__07318__A _07471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ _09873_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09903_/A sky130_fd_sc_hd__xnor2_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08824_ _08983_/B _08982_/A _08824_/C _09084_/D vssd1 vssd1 vccd1 vccd1 _08869_/A
+ sky130_fd_sc_hd__and4_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08755_ _08796_/A _08796_/B _09863_/A _09361_/C vssd1 vssd1 vccd1 vccd1 _08756_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13275__A2 _13315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _07706_/A vssd1 vssd1 vccd1 vccd1 _07706_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_54_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08686_ _08687_/A _08687_/B _08687_/C vssd1 vssd1 vccd1 vccd1 _08688_/A sky130_fd_sc_hd__a21oi_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08149__A _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08151__A1 _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _07674_/A _07674_/B _07626_/A vssd1 vssd1 vccd1 vccd1 _07672_/B sky130_fd_sc_hd__o21ai_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12894__A _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07568_ _07568_/A vssd1 vssd1 vccd1 vccd1 _14098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12786__A1 _14111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09307_ _09393_/A _09393_/B _09393_/C vssd1 vssd1 vccd1 vccd1 _09307_/X sky130_fd_sc_hd__and3_2
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07499_ _14188_/Q _07501_/A _07498_/Y _07399_/X vssd1 vssd1 vccd1 vccd1 _14188_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09238_ _09127_/B _09127_/C _09127_/A vssd1 vssd1 vccd1 vccd1 _09239_/C sky130_fd_sc_hd__o21bai_1
XFILLER_10_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13735__A0 input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ _09095_/A _09094_/B _09094_/A vssd1 vssd1 vccd1 vccd1 _09171_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__09403__A1 _09396_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11200_ _10652_/A _11180_/X _11143_/X vssd1 vssd1 vccd1 vccd1 _11213_/A sky130_fd_sc_hd__o21a_1
XFILLER_108_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12180_ _12180_/A vssd1 vssd1 vccd1 vccd1 _13831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _11131_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11132_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12134__A _12147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09167__B1 _09811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11062_ _11114_/B _11062_/B vssd1 vssd1 vccd1 vccd1 _11062_/X sky130_fd_sc_hd__and2_1
XFILLER_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07717__A1 hold14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13664__S _13670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10013_ _10013_/A _10013_/B vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__xor2_2
XFILLER_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input22_A dout1[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09443__A _09443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13266__A2 _13201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ _11965_/A vssd1 vssd1 vccd1 vccd1 _11964_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08059__A _13871_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13703_ _13703_/A vssd1 vssd1 vccd1 vccd1 _14454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10915_ _13910_/Q vssd1 vssd1 vccd1 vccd1 _11087_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11895_ _13813_/Q _11872_/X _11894_/Y _11874_/X vssd1 vssd1 vccd1 vccd1 _13753_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_output109_A _14068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13634_ input90/X _14435_/Q _13634_/S vssd1 vssd1 vccd1 vccd1 _13635_/B sky130_fd_sc_hd__mux2_1
X_10846_ _10846_/A _10846_/B _10846_/C vssd1 vssd1 vccd1 vccd1 _10846_/X sky130_fd_sc_hd__and3_1
X_13565_ _13565_/A vssd1 vssd1 vccd1 vccd1 _14414_/D sky130_fd_sc_hd__clkbuf_1
X_10777_ _10670_/B _10777_/B vssd1 vssd1 vccd1 vccd1 _10777_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08506__B _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12516_ _12515_/X _08683_/X _12520_/S vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07653__B1 _14145_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13496_ _13496_/A vssd1 vssd1 vccd1 vccd1 _14395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12447_ _14026_/Q _12438_/X _12446_/X _12435_/X vssd1 vssd1 vccd1 vccd1 _12447_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08522__A _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12378_ _12378_/A vssd1 vssd1 vccd1 vccd1 _12378_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _14163_/CLK _14117_/D vssd1 vssd1 vccd1 vccd1 _14117_/Q sky130_fd_sc_hd__dfxtp_1
X_11329_ _11291_/A _10845_/X _11328_/Y _10669_/X vssd1 vssd1 vccd1 vccd1 _13904_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14048_ _14411_/CLK _14048_/D vssd1 vssd1 vccd1 vccd1 _14048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12979__A _13010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ _06875_/A _06875_/B _06875_/C vssd1 vssd1 vccd1 vccd1 _07105_/A sky130_fd_sc_hd__nor3_2
XFILLER_41_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08540_ _09941_/B vssd1 vssd1 vccd1 vccd1 _08547_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_36_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08471_ _08590_/A _08471_/B _08471_/C vssd1 vssd1 vccd1 vccd1 _08590_/B sky130_fd_sc_hd__nand3_1
XFILLER_39_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07422_ _07431_/A _07422_/B vssd1 vssd1 vccd1 vccd1 _07422_/X sky130_fd_sc_hd__or2_1
XFILLER_91_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07353_ _07349_/X _07350_/X _07351_/X _07352_/X vssd1 vssd1 vccd1 vccd1 _07353_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07284_ _07521_/D vssd1 vssd1 vccd1 vccd1 _07519_/A sky130_fd_sc_hd__buf_2
X_09023_ _09023_/A _09023_/B _09023_/C vssd1 vssd1 vccd1 vccd1 _09025_/C sky130_fd_sc_hd__nand3_2
XFILLER_15_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07048__A _07087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09925_ _09922_/Y _10186_/A _09924_/X vssd1 vssd1 vccd1 vccd1 _10394_/A sky130_fd_sc_hd__a21o_2
XANTENNA__12889__A _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__A _11848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _10305_/B vssd1 vssd1 vccd1 vccd1 _10186_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _08941_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08810_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09787_ _09968_/A vssd1 vssd1 vccd1 vccd1 _10485_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13248__A2 _13215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ _06999_/A vssd1 vssd1 vccd1 vccd1 _14310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08738_ _08738_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _08740_/B sky130_fd_sc_hd__and2_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _08608_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08669_/X sky130_fd_sc_hd__and2b_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _11207_/A vssd1 vssd1 vccd1 vccd1 _10700_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11675_/X _11680_/B _11680_/C _11680_/D vssd1 vssd1 vccd1 vccd1 _11681_/A
+ sky130_fd_sc_hd__and4b_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _10631_/A _10644_/B vssd1 vssd1 vccd1 vccd1 _10633_/A sky130_fd_sc_hd__or2b_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13350_ _14353_/Q _13332_/X _13349_/X _13343_/X vssd1 vssd1 vccd1 vccd1 _14353_/D
+ sky130_fd_sc_hd__o211a_1
X_10562_ _13963_/Q _10562_/B vssd1 vssd1 vccd1 vccd1 _10562_/X sky130_fd_sc_hd__or2_1
XANTENNA__13708__A0 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12301_ _12304_/A vssd1 vssd1 vccd1 vccd1 _12301_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13281_ _14417_/Q _13306_/A _13280_/X vssd1 vssd1 vccd1 vccd1 _13281_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10493_ _10493_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10495_/B sky130_fd_sc_hd__xnor2_1
XFILLER_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12232_ _12233_/A vssd1 vssd1 vccd1 vccd1 _12232_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12931__A1 _14159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ input92/X vssd1 vssd1 vccd1 vccd1 _12913_/A sky130_fd_sc_hd__buf_6
XFILLER_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11114_ _11065_/Y _11114_/B _11114_/C vssd1 vssd1 vccd1 vccd1 _11114_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12094_ _12146_/A vssd1 vssd1 vccd1 vccd1 _12095_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11045_ _11262_/A _11134_/B _10963_/B _10963_/C vssd1 vssd1 vccd1 vccd1 _11048_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12695__A0 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10170__A1 _08836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12996_ _12997_/A vssd1 vssd1 vccd1 vccd1 _12996_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09901__A _10435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11947_ _11947_/A vssd1 vssd1 vccd1 vccd1 _11947_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11878_ hold36/X _11872_/X _11876_/X _11877_/Y _11874_/X vssd1 vssd1 vccd1 vccd1
+ _13748_/D sky130_fd_sc_hd__o221a_1
XFILLER_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13617_ _13617_/A vssd1 vssd1 vccd1 vccd1 _14429_/D sky130_fd_sc_hd__clkbuf_1
X_10829_ _10828_/B _10828_/C _10828_/A vssd1 vssd1 vccd1 vccd1 _10829_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12039__A _12060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13548_ _13548_/A vssd1 vssd1 vccd1 vccd1 _14409_/D sky130_fd_sc_hd__clkbuf_1
X_13479_ input88/X _14390_/Q _13494_/S vssd1 vssd1 vccd1 vccd1 _13480_/B sky130_fd_sc_hd__mux2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08252__A _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07971_ _09153_/B vssd1 vssd1 vccd1 vccd1 _08547_/A sky130_fd_sc_hd__clkbuf_2
X_09710_ _09708_/B _09708_/Y _09692_/Y _09709_/X vssd1 vssd1 vccd1 vccd1 _09710_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_68_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06922_ _14463_/Q _14287_/Q vssd1 vssd1 vccd1 vccd1 _06922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09641_ _09641_/A vssd1 vssd1 vccd1 vccd1 _09641_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09572_ _09569_/X _09570_/Y _09518_/A _09518_/Y vssd1 vssd1 vccd1 vccd1 _09573_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_71_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08523_ _08828_/A vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__buf_2
XFILLER_82_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08454_ _09134_/A vssd1 vssd1 vccd1 vccd1 _08980_/A sky130_fd_sc_hd__buf_2
XANTENNA__10464__A2 _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08427__A _08983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07405_ _07769_/S vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__buf_2
XFILLER_91_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08385_ _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _08387_/C sky130_fd_sc_hd__nand2_1
XFILLER_17_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11413__A1 _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ _07363_/A vssd1 vssd1 vccd1 vccd1 _07336_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07093__A1 _14298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07267_ _14165_/Q _14166_/Q _11663_/B _14240_/Q vssd1 vssd1 vccd1 vccd1 _07267_/X
+ sky130_fd_sc_hd__or4b_1
XANTENNA__08290__B1 _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09006_ _09072_/B _09005_/C _09005_/A vssd1 vssd1 vccd1 vccd1 _09007_/C sky130_fd_sc_hd__a21o_1
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07198_ _14278_/Q _07197_/X _07201_/S vssd1 vssd1 vccd1 vccd1 _07199_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10519__A3 _10516_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11300__B _11300_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09790__B1 _09783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09908_ _10039_/B _10065_/B vssd1 vssd1 vccd1 vccd1 _10153_/B sky130_fd_sc_hd__nor2_2
XANTENNA__12677__A0 _12936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09839_ _10004_/A _10383_/A vssd1 vssd1 vccd1 vccd1 _09968_/B sky130_fd_sc_hd__nand2_2
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12850_ _12650_/X _14131_/Q _12853_/S vssd1 vssd1 vccd1 vccd1 _12851_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_27_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11801_ _14234_/Q _13037_/A _11800_/X _14110_/Q vssd1 vssd1 vccd1 vccd1 _11801_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12781_ _14110_/Q _12771_/X _12779_/X _12780_/X _12207_/X vssd1 vssd1 vccd1 vccd1
+ _14110_/D sky130_fd_sc_hd__o221a_1
XANTENNA__12558__S _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__A1 _09091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11101__B1 _11100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _13766_/Q _11732_/B vssd1 vssd1 vccd1 vccd1 _11732_/Y sky130_fd_sc_hd__nand2_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14451_/CLK _14451_/D vssd1 vssd1 vccd1 vccd1 _14451_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11920_/A _11663_/B vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__nand2_2
XFILLER_14_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _12610_/X _14368_/Q _13408_/S vssd1 vssd1 vccd1 vccd1 _13403_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10614_ _10614_/A _10614_/B _10614_/C vssd1 vssd1 vccd1 vccd1 _10614_/Y sky130_fd_sc_hd__nand3_1
X_14382_ _14464_/CLK _14382_/D vssd1 vssd1 vccd1 vccd1 _14382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11594_ _11652_/S vssd1 vssd1 vccd1 vccd1 _11611_/S sky130_fd_sc_hd__buf_2
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13333_ _14381_/Q _13328_/X _13315_/X _14461_/Q vssd1 vssd1 vccd1 vccd1 _13333_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10545_ _10562_/B vssd1 vssd1 vccd1 vccd1 _10545_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09168__A _09216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13264_ _14333_/Q _13240_/X _13263_/X _13254_/X vssd1 vssd1 vccd1 vccd1 _14333_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10476_ _10485_/A _10477_/B vssd1 vssd1 vccd1 vccd1 _10498_/C sky130_fd_sc_hd__or2_1
XANTENNA_output176_A _14323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ _11990_/B _13059_/A _12699_/C _13835_/Q vssd1 vssd1 vccd1 vccd1 _12215_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13195_ _13332_/A vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_29_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12146_ _12146_/A vssd1 vssd1 vccd1 vccd1 _12146_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12077_ _13804_/Q _12000_/A _12021_/A _13820_/Q vssd1 vssd1 vccd1 vccd1 _12078_/B
+ sky130_fd_sc_hd__a22o_1
X_11028_ _13915_/Q vssd1 vssd1 vccd1 vccd1 _11054_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06898__A1 _14323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09053__D _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13093__A0 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14275_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12979_ _13010_/A vssd1 vssd1 vccd1 vccd1 _13004_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09836__A1 _09824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13153__A _13153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12840__A0 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08170_ _08170_/A _08170_/B _08170_/C vssd1 vssd1 vccd1 vccd1 _08170_/Y sky130_fd_sc_hd__nor3_2
XFILLER_119_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07121_ _07090_/X _07120_/X _14387_/Q vssd1 vssd1 vccd1 vccd1 _07122_/S sky130_fd_sc_hd__o21a_1
X_07052_ _14415_/Q _07059_/B _14447_/Q vssd1 vssd1 vccd1 vccd1 _07052_/X sky130_fd_sc_hd__and3b_1
Xoutput101 _14060_/Q vssd1 vssd1 vccd1 vccd1 addr1[0] sky130_fd_sc_hd__buf_2
Xoutput112 _11753_/X vssd1 vssd1 vccd1 vccd1 io_wbs_ack sky130_fd_sc_hd__buf_2
Xoutput123 _11850_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[19] sky130_fd_sc_hd__buf_2
Xoutput134 _11867_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[29] sky130_fd_sc_hd__buf_2
Xoutput145 _14301_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[0] sky130_fd_sc_hd__buf_2
Xoutput156 _14311_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[1] sky130_fd_sc_hd__buf_2
XFILLER_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput167 _14321_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[2] sky130_fd_sc_hd__buf_2
Xoutput178 _14167_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_spi_sclk_o sky130_fd_sc_hd__buf_2
XANTENNA__13328__A _13328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ _08002_/A _08658_/B _08004_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _07968_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12232__A _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06905_ _06902_/X _14322_/Q _06905_/S vssd1 vssd1 vccd1 vccd1 _06906_/A sky130_fd_sc_hd__mux2_1
X_07885_ _07885_/A _07885_/B vssd1 vssd1 vccd1 vccd1 _07886_/A sky130_fd_sc_hd__or2_1
XFILLER_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09624_ _09470_/B _09470_/C _09623_/X _09454_/Y vssd1 vssd1 vccd1 vccd1 _09624_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14100__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09555_ _09555_/A _09555_/B _09555_/C vssd1 vssd1 vccd1 vccd1 _09558_/A sky130_fd_sc_hd__nand3_1
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08506_ _09349_/A _09807_/A vssd1 vssd1 vccd1 vccd1 _08693_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09486_ _09485_/A _09485_/C _09485_/B vssd1 vssd1 vccd1 vccd1 _09488_/B sky130_fd_sc_hd__a21o_1
XFILLER_19_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08437_ _13865_/Q vssd1 vssd1 vccd1 vccd1 _09207_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13818__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07996__A _13870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ _14017_/Q vssd1 vssd1 vccd1 vccd1 _09165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07319_ _07319_/A vssd1 vssd1 vccd1 vccd1 _07464_/A sky130_fd_sc_hd__clkbuf_4
X_08299_ _08113_/A _08329_/B _08298_/Y vssd1 vssd1 vccd1 vccd1 _08301_/B sky130_fd_sc_hd__a21oi_1
X_10330_ _10354_/A _10330_/B vssd1 vssd1 vccd1 vccd1 _10332_/A sky130_fd_sc_hd__xnor2_2
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10261_ _10619_/A _10626_/B vssd1 vssd1 vccd1 vccd1 _10261_/X sky130_fd_sc_hd__or2_1
X_12000_ _12000_/A vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10192_ _10197_/A _10197_/B _09915_/X vssd1 vssd1 vccd1 vccd1 _10199_/B sky130_fd_sc_hd__a21oi_1
XFILLER_8_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _13982_/CLK _13951_/D _12371_/Y vssd1 vssd1 vccd1 vccd1 _13951_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11981__A _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12902_ _13062_/A _12902_/B vssd1 vssd1 vccd1 vccd1 _12942_/B sky130_fd_sc_hd__or2_2
XFILLER_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13882_ _14198_/CLK _13882_/D _12285_/Y vssd1 vssd1 vccd1 vccd1 _13882_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12833_ _12853_/S vssd1 vssd1 vccd1 vccd1 _12846_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10597__A _10597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ _12828_/A _13042_/B vssd1 vssd1 vccd1 vccd1 _12776_/A sky130_fd_sc_hd__nor2_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _11715_/A vssd1 vssd1 vccd1 vccd1 _11716_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11205__B _11305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ input74/X _14057_/Q _12695_/S vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__mux2_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14434_ _14467_/CLK _14434_/D vssd1 vssd1 vccd1 vccd1 _14434_/Q sky130_fd_sc_hd__dfxtp_1
X_11646_ _11646_/A _11554_/Y vssd1 vssd1 vccd1 vccd1 _11647_/B sky130_fd_sc_hd__or2b_1
Xinput14 dout1[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput25 dout1[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_2
X_14365_ _14365_/CLK _14365_/D vssd1 vssd1 vccd1 vccd1 _14365_/Q sky130_fd_sc_hd__dfxtp_2
Xinput36 io_wbs_adr[12] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
X_11577_ _11601_/A _11602_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__a21boi_4
XANTENNA__12317__A _12317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput47 io_wbs_adr[22] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
Xinput58 io_wbs_adr[3] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
X_13316_ _14377_/Q _13307_/X _13315_/X _14457_/Q vssd1 vssd1 vccd1 vccd1 _13316_/X
+ sky130_fd_sc_hd__a22o_1
Xinput69 io_wbs_datwr[12] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_1
X_10528_ _10528_/A vssd1 vssd1 vccd1 vccd1 _10528_/X sky130_fd_sc_hd__buf_2
X_14296_ _14411_/CLK _14296_/D _13162_/Y vssd1 vssd1 vccd1 vccd1 _14296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13247_ _14410_/Q _13230_/X _13246_/X vssd1 vssd1 vccd1 vccd1 _13247_/X sky130_fd_sc_hd__a21o_1
X_10459_ _10411_/A _10459_/B vssd1 vssd1 vccd1 vccd1 _10459_/X sky130_fd_sc_hd__and2b_1
X_13178_ _13178_/A vssd1 vssd1 vccd1 vccd1 _13183_/A sky130_fd_sc_hd__buf_2
XFILLER_112_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06969__B _14281_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _13815_/Q _12117_/X _12128_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _13815_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13302__A1 _14341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07670_ _07670_/A _07670_/B vssd1 vssd1 vccd1 vccd1 _07744_/A sky130_fd_sc_hd__xnor2_2
XFILLER_42_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13066__A0 _12633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09340_ _09340_/A _09340_/B vssd1 vssd1 vccd1 vccd1 _09340_/X sky130_fd_sc_hd__or2_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11616__A1 _11614_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ _09271_/A _09271_/B _09271_/C vssd1 vssd1 vccd1 vccd1 _09273_/A sky130_fd_sc_hd__or3_4
XFILLER_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ _08223_/B _08223_/C _08243_/A vssd1 vssd1 vccd1 vccd1 _08224_/A sky130_fd_sc_hd__a21oi_1
XFILLER_105_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08153_ _08198_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08154_/B sky130_fd_sc_hd__or2_1
XFILLER_119_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07104_ _14264_/Q _07085_/X _07103_/X _14360_/Q vssd1 vssd1 vccd1 vccd1 _07104_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08084_ _08122_/A vssd1 vssd1 vccd1 vccd1 _08084_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07035_ _14417_/Q _07059_/B _14449_/Q vssd1 vssd1 vccd1 vccd1 _07035_/X sky130_fd_sc_hd__and3b_1
XFILLER_115_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08440__A _08982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _08986_/A _08986_/B _08986_/C vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__nand3_1
XFILLER_76_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07937_ _13869_/Q vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__buf_2
XFILLER_21_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07868_ _07868_/A _07868_/B vssd1 vssd1 vccd1 vccd1 _07869_/B sky130_fd_sc_hd__nand2_1
XFILLER_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ _09607_/A _09607_/B _09607_/C vssd1 vssd1 vccd1 vccd1 _09675_/A sky130_fd_sc_hd__and3_1
XFILLER_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07799_ _13947_/Q vssd1 vssd1 vccd1 vccd1 _10931_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_73_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11607__A1 _11606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ _09538_/A _09538_/B vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__xor2_1
XFILLER_58_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09421__D _10613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09469_ _09452_/X _09453_/Y _09423_/A _09423_/Y vssd1 vssd1 vccd1 vccd1 _09470_/D
+ sky130_fd_sc_hd__o211ai_1
XFILLER_40_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11500_ _11014_/B _11489_/X _11499_/X _11285_/A _11490_/X vssd1 vssd1 vccd1 vccd1
+ _11500_/X sky130_fd_sc_hd__o221a_1
XANTENNA__13521__A _13592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12480_ _13998_/Q _12460_/X _12478_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _13998_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _11431_/A vssd1 vssd1 vccd1 vccd1 _11493_/B sky130_fd_sc_hd__inv_2
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12137__A input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14150_ _14152_/CLK _14150_/D vssd1 vssd1 vccd1 vccd1 _14150_/Q sky130_fd_sc_hd__dfxtp_1
X_11362_ _11362_/A vssd1 vssd1 vccd1 vccd1 _11392_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10594__A1 _10565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ _13101_/A vssd1 vssd1 vccd1 vccd1 _14251_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13667__S _13670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__xor2_1
X_14081_ _14217_/CLK _14081_/D _12726_/Y vssd1 vssd1 vccd1 vccd1 _14081_/Q sky130_fd_sc_hd__dfrtp_4
X_11293_ _11327_/A _11331_/A _11328_/A vssd1 vssd1 vccd1 vccd1 _11324_/C sky130_fd_sc_hd__o21bai_1
XANTENNA__08539__A1 _08966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ _13032_/A vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input52_A io_wbs_adr[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10244_ _10244_/A _10244_/B vssd1 vssd1 vccd1 vccd1 _10250_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08350__A _13866_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10175_ _10160_/Y _10175_/B vssd1 vssd1 vccd1 vccd1 _10176_/A sky130_fd_sc_hd__and2b_1
XFILLER_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output139_A _11813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A1 _14341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13934_ _14102_/CLK _13934_/D _12350_/Y vssd1 vssd1 vccd1 vccd1 _13934_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13865_ _13867_/CLK _13865_/D _12265_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12816_ hold7/X _12772_/X _12803_/A _14146_/Q _12809_/X vssd1 vssd1 vccd1 vccd1 _12816_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13796_ _14400_/CLK _13796_/D vssd1 vssd1 vccd1 vccd1 _13796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12753_/A vssd1 vssd1 vccd1 vccd1 _12752_/A sky130_fd_sc_hd__buf_2
XFILLER_72_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _12678_/A _12678_/B vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__and2_1
XFILLER_30_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14417_ _14417_/CLK _14417_/D vssd1 vssd1 vccd1 vccd1 _14417_/Q sky130_fd_sc_hd__dfxtp_1
X_11629_ _11629_/A vssd1 vssd1 vccd1 vccd1 _13847_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12047__A _13609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14348_ _14348_/CLK _14348_/D vssd1 vssd1 vccd1 vccd1 _14348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07450__A1 _14084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14279_ _14281_/CLK _14279_/D _13140_/Y vssd1 vssd1 vccd1 vccd1 _14279_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11534__A0 _10206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08811_/A _08811_/B _08811_/C vssd1 vssd1 vccd1 vccd1 _08840_/X sky130_fd_sc_hd__a21o_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08771_/A _08771_/B _08771_/C vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_0_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14256_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07722_ hold1/X _07754_/B vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__and2_1
XFILLER_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11837__B2 _14121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__B _09803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09091__A _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _07716_/A _07716_/B _14145_/Q vssd1 vssd1 vccd1 vccd1 _07653_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07584_ _07595_/A vssd1 vssd1 vccd1 vccd1 _07593_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_81_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14019__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ _09346_/A _09321_/C _09321_/B vssd1 vssd1 vccd1 vccd1 _09324_/C sky130_fd_sc_hd__a21o_1
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13341__A _13341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09254_ _09276_/A _09276_/B _09276_/C vssd1 vssd1 vccd1 vccd1 _09254_/Y sky130_fd_sc_hd__nor3_2
XANTENNA__08435__A _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ _09769_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08217_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12014__B2 _13827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ _09184_/B _09184_/C _09184_/A vssd1 vssd1 vccd1 vccd1 _09185_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08136_ _08208_/C vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_88_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07993__B _09999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _08002_/A _08132_/D _07999_/B _07997_/X vssd1 vssd1 vccd1 vccd1 _08124_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_49_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07018_ _14419_/Q _07017_/Y _07009_/X vssd1 vssd1 vccd1 vccd1 _07018_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08969_ _09044_/A _09998_/A vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11980_ _12233_/A vssd1 vssd1 vccd1 vccd1 _11980_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ _10931_/A vssd1 vssd1 vccd1 vccd1 _11169_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_5_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13650_ input91/X _14439_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13651_/B sky130_fd_sc_hd__mux2_1
X_10862_ _10675_/X _10860_/X _10861_/Y vssd1 vssd1 vccd1 vccd1 _13937_/D sky130_fd_sc_hd__o21ai_1
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12789__C1 _12207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12601_ _12615_/A _12601_/B vssd1 vssd1 vccd1 vccd1 _12602_/A sky130_fd_sc_hd__and2_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _13590_/A _13581_/B vssd1 vssd1 vccd1 vccd1 _13582_/A sky130_fd_sc_hd__and2_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ _10889_/B _10889_/C _10889_/A vssd1 vssd1 vccd1 vccd1 _10884_/C sky130_fd_sc_hd__o21ai_1
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12532_ _12532_/A vssd1 vssd1 vccd1 vccd1 _14013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08345__A _13866_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ _13994_/Q _12460_/X _12462_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _13994_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11414_ _11525_/A _11525_/B vssd1 vssd1 vccd1 vccd1 _11521_/A sky130_fd_sc_hd__or2_1
X_14202_ _14211_/CLK _14202_/D _12994_/Y vssd1 vssd1 vccd1 vccd1 _14202_/Q sky130_fd_sc_hd__dfrtp_1
X_12394_ _12397_/A vssd1 vssd1 vccd1 vccd1 _12394_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10567__A1 _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ _14149_/CLK _14133_/D vssd1 vssd1 vccd1 vccd1 _14133_/Q sky130_fd_sc_hd__dfxtp_1
X_11345_ _11345_/A _11345_/B vssd1 vssd1 vccd1 vccd1 _11345_/X sky130_fd_sc_hd__and2_1
XFILLER_4_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14064_ _14065_/CLK _14064_/D _12706_/Y vssd1 vssd1 vccd1 vccd1 _14064_/Q sky130_fd_sc_hd__dfrtp_1
X_11276_ _11276_/A _11276_/B vssd1 vssd1 vccd1 vccd1 _11277_/B sky130_fd_sc_hd__nor2_1
XFILLER_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08080__A _08146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13015_ _13016_/A vssd1 vssd1 vccd1 vccd1 _13015_/Y sky130_fd_sc_hd__inv_2
X_10227_ _10227_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10232_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10158_ _10172_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10175_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12330__A _12348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10089_ _10127_/A _10087_/X _10088_/X vssd1 vssd1 vccd1 vccd1 _10333_/A sky130_fd_sc_hd__o21ai_4
XFILLER_43_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13917_ _13920_/CLK _13917_/D _12329_/Y vssd1 vssd1 vccd1 vccd1 _13917_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__07499__B2 _07399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13848_ _14028_/CLK _13848_/D _12242_/Y vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfrtp_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13779_ _14427_/CLK _13779_/D _11976_/Y vssd1 vssd1 vccd1 vccd1 _13779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09941_ _09941_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__or2_2
XANTENNA__11507__B1 _10686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09872_ _09872_/A _09872_/B vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__nor2_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08923__A1 _09188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08823_/A vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__buf_6
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13336__A _13336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08754_ _08828_/B _08629_/A _09882_/A _08828_/A vssd1 vssd1 vccd1 vccd1 _08756_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_22_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12240__A _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _14075_/Q _07619_/Y _07703_/X _07704_/Y vssd1 vssd1 vccd1 vccd1 _14075_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _08683_/X _10009_/A _08605_/X _08604_/X _08767_/B vssd1 vssd1 vccd1 vccd1
+ _08687_/C sky130_fd_sc_hd__a32oi_4
XANTENNA__12483__A1 _14034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08151__A2 _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07636_ _07675_/A _07676_/A _07675_/B vssd1 vssd1 vccd1 vccd1 _07674_/B sky130_fd_sc_hd__a21boi_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07567_ _14098_/Q input15/X _07571_/S vssd1 vssd1 vccd1 vccd1 _07568_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10695__A _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09306_ _09294_/A _09294_/B _09294_/C vssd1 vssd1 vccd1 vccd1 _09393_/C sky130_fd_sc_hd__a21o_1
XFILLER_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07498_ _14188_/Q _14187_/Q _07534_/B vssd1 vssd1 vccd1 vccd1 _07498_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07111__B1 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__A _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09237_ _08867_/A _09824_/A _09236_/A _09236_/C vssd1 vssd1 vccd1 vccd1 _09239_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _09216_/A _09168_/B _09168_/C vssd1 vssd1 vccd1 vccd1 _09171_/A sky130_fd_sc_hd__or3_1
XANTENNA__09403__A2 _09397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07414__A1 _07399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ _09590_/A _08119_/B _08119_/C vssd1 vssd1 vccd1 vccd1 _08120_/B sky130_fd_sc_hd__and3_1
X_09099_ _09097_/A _09097_/C _09097_/B vssd1 vssd1 vccd1 vccd1 _09100_/C sky130_fd_sc_hd__a21o_1
XANTENNA__07414__B2 _14208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11130_ _11119_/X _11127_/C _11129_/Y _10851_/B _11038_/A vssd1 vssd1 vccd1 vccd1
+ _13913_/D sky130_fd_sc_hd__a32o_1
XANTENNA__09167__A1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11062_/B sky130_fd_sc_hd__or2_1
XFILLER_95_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10012_ _10382_/B _10006_/B _10015_/A vssd1 vssd1 vccd1 vccd1 _10244_/A sky130_fd_sc_hd__o21ai_2
XFILLER_62_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12150__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__B _09493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input15_A dout1[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12474__A1 _14032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11963_ _11965_/A vssd1 vssd1 vccd1 vccd1 _11963_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13702_ _13712_/A _13702_/B vssd1 vssd1 vccd1 vccd1 _13703_/A sky130_fd_sc_hd__and2_1
XFILLER_45_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10914_ _13910_/Q _10913_/X _10953_/A vssd1 vssd1 vccd1 vccd1 _10914_/X sky130_fd_sc_hd__mux2_1
X_11894_ _11897_/B _11894_/B vssd1 vssd1 vccd1 vccd1 _11894_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13633_ _13633_/A vssd1 vssd1 vccd1 vccd1 _14434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10845_ _11100_/A vssd1 vssd1 vccd1 vccd1 _10845_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_73_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10776_ _07804_/B _10663_/Y _10936_/A _10670_/Y _10748_/B vssd1 vssd1 vccd1 vccd1
+ _10905_/B sky130_fd_sc_hd__o221ai_4
X_13564_ _13573_/A _13564_/B vssd1 vssd1 vccd1 vccd1 _13565_/A sky130_fd_sc_hd__and2_1
XFILLER_13_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12515_ input77/X vssd1 vssd1 vccd1 vccd1 _12515_/X sky130_fd_sc_hd__buf_4
X_13495_ _13502_/A _13495_/B vssd1 vssd1 vccd1 vccd1 _13496_/A sky130_fd_sc_hd__and2_1
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12446_ _08946_/A _12439_/X _12442_/X _14042_/Q vssd1 vssd1 vccd1 vccd1 _12446_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ _12378_/A vssd1 vssd1 vccd1 vccd1 _12377_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11328_ _11328_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11328_/Y sky130_fd_sc_hd__xnor2_1
X_14116_ _14258_/CLK _14116_/D vssd1 vssd1 vccd1 vccd1 _14116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11259_ _11269_/A _11269_/B vssd1 vssd1 vccd1 vccd1 _11347_/A sky130_fd_sc_hd__nand2_1
X_14047_ _14363_/CLK _14047_/D vssd1 vssd1 vccd1 vccd1 _14047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09634__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06916__B1 _06877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12060__A _12060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08470_ _08470_/A _08470_/B vssd1 vssd1 vccd1 vccd1 _08471_/C sky130_fd_sc_hd__xnor2_1
XFILLER_78_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07421_ _14205_/Q _14207_/Q _07442_/S vssd1 vssd1 vccd1 vccd1 _07422_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12217__A1 _12209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07352_ _07491_/A vssd1 vssd1 vccd1 vccd1 _07352_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07283_ _14165_/D _14166_/D vssd1 vssd1 vccd1 vccd1 _07521_/D sky130_fd_sc_hd__or2_1
XANTENNA__10243__A3 _10645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ _09022_/A _09022_/B vssd1 vssd1 vccd1 vccd1 _09023_/C sky130_fd_sc_hd__or2_1
XFILLER_102_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12925__C1 _12920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09924_ _10004_/A _10004_/B vssd1 vssd1 vccd1 vccd1 _09924_/X sky130_fd_sc_hd__and2_1
XFILLER_113_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A dout1[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _09482_/B _09848_/X _09847_/X vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__a21o_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _08805_/C _08805_/B _08850_/A vssd1 vssd1 vccd1 vccd1 _08811_/B sky130_fd_sc_hd__a21bo_1
XFILLER_65_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06998_ _06995_/X _14310_/Q _06998_/S vssd1 vssd1 vccd1 vccd1 _06999_/A sky130_fd_sc_hd__mux2_1
XANTENNA__07580__A0 _14092_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09786_ _09786_/A vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__inv_2
XFILLER_67_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08737_ _08617_/A _08616_/B _08616_/C vssd1 vssd1 vccd1 vccd1 _08738_/B sky130_fd_sc_hd__a21o_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13653__A0 input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12456__A1 _14028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08668_ _08667_/B _08667_/C _08667_/A vssd1 vssd1 vccd1 vccd1 _08668_/X sky130_fd_sc_hd__a21o_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07619_ _07765_/S vssd1 vssd1 vccd1 vccd1 _07619_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13405__A0 _12681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _08595_/X _08599_/B vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__and2b_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10629__S _10629_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10630_ _10630_/A vssd1 vssd1 vccd1 vccd1 _13954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10561_ _10561_/A _10561_/B vssd1 vssd1 vccd1 vccd1 _10561_/Y sky130_fd_sc_hd__nor2_2
X_12300_ _12304_/A vssd1 vssd1 vccd1 vccd1 _12300_/Y sky130_fd_sc_hd__inv_2
X_13280_ _14449_/Q _13250_/X _13245_/A _14401_/Q vssd1 vssd1 vccd1 vccd1 _13280_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10492_ _10492_/A _10492_/B vssd1 vssd1 vccd1 vccd1 _10493_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08623__A _08623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ _12231_/A vssd1 vssd1 vccd1 vccd1 _13839_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12162_ _13826_/Q _12146_/X _12160_/X _12161_/X vssd1 vssd1 vccd1 vccd1 _13826_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11113_ _11010_/B _11110_/X _11111_/X _11112_/Y vssd1 vssd1 vccd1 vccd1 _13920_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11984__A input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12093_ _12900_/A _12092_/Y vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__nor2b_4
XFILLER_2_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11044_ _13944_/Q _11044_/B _10963_/B _10963_/C vssd1 vssd1 vccd1 vccd1 _11048_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12695__A1 _14057_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__A0 _14096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12447__A1 _14026_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ _12997_/A vssd1 vssd1 vccd1 vccd1 _12995_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09312__A1 _08823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09312__B2 _08445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11946_ _11947_/A vssd1 vssd1 vccd1 vccd1 _11946_/Y sky130_fd_sc_hd__inv_2
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _13748_/Q _13747_/Q vssd1 vssd1 vccd1 vccd1 _11877_/Y sky130_fd_sc_hd__nor2_1
X_13616_ _13625_/A _13616_/B vssd1 vssd1 vccd1 vccd1 _13617_/A sky130_fd_sc_hd__and2_1
X_10828_ _10828_/A _10828_/B _10828_/C vssd1 vssd1 vccd1 vccd1 _10828_/Y sky130_fd_sc_hd__nand3_1
XFILLER_60_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13547_ _13556_/A _13547_/B vssd1 vssd1 vccd1 vccd1 _13548_/A sky130_fd_sc_hd__and2_1
X_10759_ _10769_/A vssd1 vssd1 vccd1 vccd1 _10765_/A sky130_fd_sc_hd__inv_2
XFILLER_12_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09629__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13478_ _13522_/S vssd1 vssd1 vccd1 vccd1 _13494_/S sky130_fd_sc_hd__clkbuf_2
X_12429_ _12429_/A _13202_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _12440_/B sky130_fd_sc_hd__and3_1
XFILLER_114_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07149__A _11663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07970_ _14019_/Q vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__buf_2
XFILLER_114_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06921_ _06921_/A vssd1 vssd1 vccd1 vccd1 _14320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09640_ _09638_/A _09636_/Y _09634_/Y _09635_/Y vssd1 vssd1 vccd1 vccd1 _09640_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10303__A _10420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ _09518_/A _09518_/Y _09569_/X _09570_/Y vssd1 vssd1 vccd1 vccd1 _09573_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_36_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08522_ _09844_/A vssd1 vssd1 vccd1 vccd1 _09000_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09811__B _09811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08453_ _08592_/B _08452_/C _08452_/B vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__a21o_1
XFILLER_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07404_ _11746_/S vssd1 vssd1 vccd1 vccd1 _07404_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08384_ _08384_/A _08384_/B vssd1 vssd1 vccd1 vccd1 _08387_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07335_ _14222_/Q _07311_/X _07316_/X _07334_/X vssd1 vssd1 vccd1 vccd1 _14222_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07266_ _13951_/Q _07769_/S vssd1 vssd1 vccd1 vccd1 _07266_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08443__A _13863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09005_ _09005_/A _09072_/B _09005_/C vssd1 vssd1 vccd1 vccd1 _09007_/B sky130_fd_sc_hd__nand3_1
XFILLER_3_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07197_ _14094_/Q _07185_/X _07186_/X vssd1 vssd1 vccd1 vccd1 _07197_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09907_ _10039_/B _10065_/B vssd1 vssd1 vccd1 vccd1 _10171_/B sky130_fd_sc_hd__xor2_4
XANTENNA__13747__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12677__A1 _14052_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_2_0_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09838_ _09838_/A vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__buf_2
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09769_ _09769_/A _09769_/B vssd1 vssd1 vccd1 vccd1 _09770_/B sky130_fd_sc_hd__xnor2_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11800_ _12768_/A vssd1 vssd1 vccd1 vccd1 _11800_/X sky130_fd_sc_hd__buf_2
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _14135_/Q _12776_/X _12760_/X vssd1 vssd1 vccd1 vccd1 _12780_/X sky130_fd_sc_hd__a21o_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11101__B2 _11079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _11716_/A _11729_/Y _11730_/X _11714_/A _13767_/Q vssd1 vssd1 vccd1 vccd1
+ _13767_/D sky130_fd_sc_hd__a32o_1
XFILLER_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _14450_/CLK _14450_/D vssd1 vssd1 vccd1 vccd1 _14450_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11662_ hold6/X vssd1 vssd1 vccd1 vccd1 _11920_/A sky130_fd_sc_hd__buf_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13401_/A vssd1 vssd1 vccd1 vccd1 _14367_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11979__A _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10613_ _10613_/A _10613_/B _10613_/C vssd1 vssd1 vccd1 vccd1 _10614_/C sky130_fd_sc_hd__or3_1
X_14381_ _14465_/CLK _14381_/D vssd1 vssd1 vccd1 vccd1 _14381_/Q sky130_fd_sc_hd__dfxtp_1
X_11593_ _11615_/A vssd1 vssd1 vccd1 vccd1 _11652_/S sky130_fd_sc_hd__clkbuf_2
X_13332_ _13332_/A vssd1 vssd1 vccd1 vccd1 _13332_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input82_A io_wbs_datwr[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ _10544_/A vssd1 vssd1 vccd1 vccd1 _13965_/D sky130_fd_sc_hd__clkbuf_1
X_13263_ _14365_/Q _13208_/X _13262_/X _13258_/X vssd1 vssd1 vccd1 vccd1 _13263_/X
+ sky130_fd_sc_hd__a211o_1
X_10475_ _10498_/B _10475_/B vssd1 vssd1 vccd1 vccd1 _10477_/B sky130_fd_sc_hd__nand2_1
XFILLER_109_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12214_ _13059_/A _12699_/C vssd1 vssd1 vccd1 vccd1 _12226_/B sky130_fd_sc_hd__nand2_1
X_13194_ _13194_/A _13209_/A _13194_/C vssd1 vssd1 vccd1 vccd1 _13332_/A sky130_fd_sc_hd__and3_4
XANTENNA_output169_A _14294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _13821_/Q _12133_/X _12143_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _13821_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12603__A _12611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12076_ _12076_/A vssd1 vssd1 vccd1 vccd1 _13803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11027_ _11056_/A _11056_/B vssd1 vssd1 vccd1 vccd1 _11120_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08528__A _09241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ _12978_/A vssd1 vssd1 vccd1 vccd1 _12978_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09836__A2 _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07432__A _11746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _12046_/A vssd1 vssd1 vccd1 vccd1 _12933_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07120_ _14435_/Q _07134_/B _14467_/Q vssd1 vssd1 vccd1 vccd1 _07120_/X sky130_fd_sc_hd__and3b_1
XANTENNA__10603__B1 _10613_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07051_ _07090_/A vssd1 vssd1 vccd1 vccd1 _07051_/X sky130_fd_sc_hd__clkbuf_2
Xoutput102 _14061_/Q vssd1 vssd1 vccd1 vccd1 addr1[1] sky130_fd_sc_hd__buf_2
Xoutput113 _11786_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[0] sky130_fd_sc_hd__buf_2
Xoutput124 _11791_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[1] sky130_fd_sc_hd__buf_2
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput135 _11803_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[2] sky130_fd_sc_hd__buf_2
Xoutput146 _14302_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[10] sky130_fd_sc_hd__buf_2
XFILLER_82_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput157 _14312_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[20] sky130_fd_sc_hd__buf_2
XFILLER_114_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput168 _14322_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[30] sky130_fd_sc_hd__buf_2
XANTENNA__13609__A _13609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput179 _14169_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_spi_sdo_o sky130_fd_sc_hd__buf_2
XFILLER_86_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12513__A _12517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07953_ _09793_/A vssd1 vssd1 vccd1 vccd1 _08658_/B sky130_fd_sc_hd__buf_6
XFILLER_68_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06904_ _06894_/X _06903_/X _14386_/Q vssd1 vssd1 vccd1 vccd1 _06905_/S sky130_fd_sc_hd__o21a_1
X_07884_ _07884_/A vssd1 vssd1 vccd1 vccd1 _13980_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09623_ _09452_/X _09453_/Y _09423_/A _09423_/Y vssd1 vssd1 vccd1 vccd1 _09623_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09822__A _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09554_ _09554_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11095__B1 _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ _09869_/A vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__buf_2
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07838__A1 _14027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09485_ _09485_/A _09485_/B _09485_/C vssd1 vssd1 vccd1 vccd1 _09488_/A sky130_fd_sc_hd__nand3_1
X_08436_ _08789_/A vssd1 vssd1 vccd1 vccd1 _08982_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08367_ _08716_/B vssd1 vssd1 vccd1 vccd1 _08842_/A sky130_fd_sc_hd__buf_6
XFILLER_108_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07318_ _07471_/A vssd1 vssd1 vccd1 vccd1 _07521_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_20_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08298_ _08298_/A _08298_/B vssd1 vssd1 vccd1 vccd1 _08298_/Y sky130_fd_sc_hd__nor2_1
X_07249_ _14079_/Q _13879_/Q _07252_/S vssd1 vssd1 vccd1 vccd1 _07249_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10260_ _10260_/A _10260_/B vssd1 vssd1 vccd1 vccd1 _10626_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10191_ _10191_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10199_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12423__A input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13950_ _13950_/CLK _13950_/D _12370_/Y vssd1 vssd1 vccd1 vccd1 _13950_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12901_ _12928_/A vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13881_ _14275_/CLK _13881_/D _12284_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13254__A _13254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _13072_/A vssd1 vssd1 vccd1 vccd1 _12847_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_28_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08348__A _14021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12828_/A _12900_/A vssd1 vssd1 vccd1 vccd1 _12801_/A sky130_fd_sc_hd__nor2_2
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11714_/A vssd1 vssd1 vccd1 vccd1 _11714_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10833__B1 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12694_/A vssd1 vssd1 vccd1 vccd1 _14056_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14465_/CLK _14433_/D vssd1 vssd1 vccd1 vccd1 _14433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11645_ _11645_/A vssd1 vssd1 vccd1 vccd1 _13843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 dout1[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14364_ _14365_/CLK _14364_/D vssd1 vssd1 vccd1 vccd1 _14364_/Q sky130_fd_sc_hd__dfxtp_2
Xinput26 dout1[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
X_11576_ _14053_/Q _13965_/Q vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput37 io_wbs_adr[13] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 io_wbs_adr[23] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
Xinput59 io_wbs_adr[4] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_2
X_13315_ _13315_/A vssd1 vssd1 vccd1 vccd1 _13315_/X sky130_fd_sc_hd__clkbuf_2
X_10527_ _13967_/Q _07924_/X _10522_/X _10526_/X vssd1 vssd1 vccd1 vccd1 _13967_/D
+ sky130_fd_sc_hd__a22o_1
X_14295_ _14410_/CLK _14295_/D _13161_/Y vssd1 vssd1 vccd1 vccd1 _14295_/Q sky130_fd_sc_hd__dfrtp_4
X_13246_ _14442_/Q _13336_/A _13245_/X _14394_/Q vssd1 vssd1 vccd1 vccd1 _13246_/X
+ sky130_fd_sc_hd__a22o_1
X_10458_ _10564_/A _10564_/B _10418_/X _10461_/A vssd1 vssd1 vccd1 vccd1 _10458_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08557__A2 _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13429__A _13504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13177_ _13177_/A vssd1 vssd1 vccd1 vccd1 _13177_/Y sky130_fd_sc_hd__inv_2
X_10389_ _10391_/B _10391_/C _10391_/A vssd1 vssd1 vccd1 vccd1 _10404_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12128_ input73/X _12130_/B vssd1 vssd1 vccd1 vccd1 _12128_/X sky130_fd_sc_hd__or2_1
XFILLER_96_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12059_ _12059_/A vssd1 vssd1 vccd1 vccd1 _12059_/X sky130_fd_sc_hd__buf_2
XFILLER_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14418__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__B _14261_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09270_ _09114_/A _09114_/C _09114_/B vssd1 vssd1 vccd1 vccd1 _09271_/C sky130_fd_sc_hd__o21ba_2
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08221_ _08221_/A _08221_/B _08221_/C vssd1 vssd1 vccd1 vccd1 _08226_/B sky130_fd_sc_hd__and3_1
XFILLER_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08705__B _09132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08152_ _08198_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08223_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07103_ _14408_/Q _07102_/Y _07087_/X vssd1 vssd1 vccd1 vccd1 _07103_/X sky130_fd_sc_hd__a21o_1
X_08083_ _08325_/A _08052_/Y _08160_/C _08082_/Y vssd1 vssd1 vccd1 vccd1 _08122_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_119_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07034_ _14273_/Q _07007_/X _07033_/X _14369_/Q vssd1 vssd1 vccd1 vccd1 _07034_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08440__B _08794_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07337__A _14104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _08449_/B _09848_/B _09804_/A _09233_/A vssd1 vssd1 vccd1 vccd1 _08986_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_102_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07056__B _14270_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ _09123_/C vssd1 vssd1 vccd1 vccd1 _09233_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_69_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14098__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ _07859_/Y _07865_/X _07890_/A _13984_/Q vssd1 vssd1 vccd1 vccd1 _13984_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_84_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09606_ _09603_/X _09604_/Y _09592_/B _09592_/Y vssd1 vssd1 vccd1 vccd1 _09607_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_84_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07798_ _07798_/A vssd1 vssd1 vccd1 vccd1 _10676_/A sky130_fd_sc_hd__buf_2
XFILLER_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09537_ _09537_/A _09537_/B vssd1 vssd1 vccd1 vccd1 _09538_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12804__A1 _14157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09468_ _09468_/A _09468_/B vssd1 vssd1 vccd1 vccd1 _09470_/C sky130_fd_sc_hd__nand2_1
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08419_ _09206_/B vssd1 vssd1 vccd1 vccd1 _10215_/A sky130_fd_sc_hd__buf_4
XANTENNA__13935__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09399_ _09399_/A _09399_/B vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__nor2_2
XANTENNA__11322__A _11322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11430_ _11288_/A _11010_/B _11436_/S vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11361_ _13893_/Q _13951_/D _11358_/X _11360_/Y vssd1 vssd1 vccd1 vccd1 _13893_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13100_ _13106_/A _13100_/B vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__and2_1
X_10312_ _10288_/A _10288_/B _10311_/Y vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__a21oi_1
X_11292_ _11324_/B _11292_/B vssd1 vssd1 vccd1 vccd1 _11328_/A sky130_fd_sc_hd__nand2_1
X_14080_ _14283_/CLK _14080_/D _12725_/Y vssd1 vssd1 vccd1 vccd1 _14080_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__08539__A2 _08658_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13031_ _13037_/B _13059_/B vssd1 vssd1 vccd1 vccd1 _13032_/A sky130_fd_sc_hd__nand2_2
XFILLER_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10243_ _10638_/B _10645_/A _10645_/B _10241_/X _10637_/A vssd1 vssd1 vccd1 vccd1
+ _10626_/A sky130_fd_sc_hd__o311a_2
XANTENNA__12153__A input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_117_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10174_ _10174_/A _10174_/B vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_input45_A io_wbs_adr[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11992__A input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13933_ _13947_/CLK _13933_/D _12349_/Y vssd1 vssd1 vccd1 vccd1 _13933_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13864_ _13867_/CLK _13864_/D _12264_/Y vssd1 vssd1 vccd1 vccd1 _13864_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__13048__A1 _14235_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12815_ _14120_/Q _12800_/X _12814_/X _12805_/X vssd1 vssd1 vccd1 vccd1 _14120_/D
+ sky130_fd_sc_hd__o211a_1
X_13795_ _14335_/CLK _13795_/D vssd1 vssd1 vccd1 vccd1 _13795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _12746_/A vssd1 vssd1 vccd1 vccd1 _12746_/Y sky130_fd_sc_hd__inv_2
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12677_ _12936_/A _14052_/Q _12685_/S vssd1 vssd1 vccd1 vccd1 _12678_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14416_ _14449_/CLK _14416_/D vssd1 vssd1 vccd1 vccd1 _14416_/Q sky130_fd_sc_hd__dfxtp_1
X_11628_ _13847_/Q _11627_/Y _11632_/S vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_3_1_0_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_io_wbs_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14347_ _14354_/CLK _14347_/D vssd1 vssd1 vccd1 vccd1 _14347_/Q sky130_fd_sc_hd__dfxtp_1
X_11559_ _11548_/X _11639_/B _11638_/A vssd1 vssd1 vccd1 vccd1 _11634_/C sky130_fd_sc_hd__a21oi_1
XFILLER_116_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08541__A _08547_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14278_ _14281_/CLK _14278_/D _13139_/Y vssd1 vssd1 vccd1 vccd1 _14278_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13229_ _14326_/Q _13196_/X _13227_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _14326_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _08770_/A _08770_/B vssd1 vssd1 vccd1 vccd1 _08771_/C sky130_fd_sc_hd__xnor2_1
XFILLER_112_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07721_ _07723_/A vssd1 vssd1 vccd1 vccd1 _07754_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09091__B _09091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _14071_/Q _07660_/A _14072_/Q vssd1 vssd1 vccd1 vccd1 _07716_/B sky130_fd_sc_hd__a21oi_2
XFILLER_92_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_41_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07583_ _07583_/A vssd1 vssd1 vccd1 vccd1 _14091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09322_ _09225_/A _09225_/C _09225_/B vssd1 vssd1 vccd1 vccd1 _09324_/B sky130_fd_sc_hd__a21bo_1
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08716__A _08716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09253_ _09276_/A _09276_/C _09276_/B vssd1 vssd1 vccd1 vccd1 _09253_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08435__B _10215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08204_ _08215_/A vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__clkbuf_2
X_09184_ _09184_/A _09184_/B _09184_/C vssd1 vssd1 vccd1 vccd1 _09184_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__13211__A1 _14356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08135_ _08135_/A vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08066_ _08140_/B _08066_/B vssd1 vssd1 vccd1 vccd1 _08124_/A sky130_fd_sc_hd__nor2_1
XFILLER_108_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07017_ _14451_/Q _14275_/Q vssd1 vssd1 vccd1 vccd1 _07017_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10959__S0 _11175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12701__A _12703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _09962_/B vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__buf_6
XANTENNA__06952__A1 _14316_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07919_ _07918_/X _13971_/Q _07919_/S vssd1 vssd1 vccd1 vccd1 _07920_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11828__A2 _11855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08899_ _08899_/A vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__buf_4
XFILLER_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10930_ _10951_/A _11158_/S vssd1 vssd1 vccd1 vccd1 _10971_/A sky130_fd_sc_hd__or2_1
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10861_ _13937_/Q _11110_/A vssd1 vssd1 vccd1 vccd1 _10861_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12926_/A _14033_/Q _12600_/S vssd1 vssd1 vccd1 vccd1 _12601_/B sky130_fd_sc_hd__mux2_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ _12688_/X _14419_/Q _13593_/S vssd1 vssd1 vccd1 vccd1 _13581_/B sky130_fd_sc_hd__mux2_1
XFILLER_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10792_ _10884_/B _10792_/B vssd1 vssd1 vccd1 vccd1 _10889_/A sky130_fd_sc_hd__and2_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12534_/A _12531_/B vssd1 vssd1 vccd1 vccd1 _12532_/A sky130_fd_sc_hd__and2_1
XANTENNA__12148__A input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12462_ _14029_/Q _12438_/X _12461_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _12462_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09406__B1 _09404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14201_ _14215_/CLK _14201_/D _12993_/Y vssd1 vssd1 vccd1 vccd1 _14201_/Q sky130_fd_sc_hd__dfrtp_1
X_11413_ _11269_/A _11038_/A _11415_/A vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11987__A input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ _12397_/A vssd1 vssd1 vccd1 vccd1 _12393_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _14250_/CLK _14132_/D vssd1 vssd1 vccd1 vccd1 _14132_/Q sky130_fd_sc_hd__dfxtp_2
X_11344_ _11344_/A _11344_/B _11344_/C vssd1 vssd1 vccd1 vccd1 _11345_/B sky130_fd_sc_hd__nand3_1
XANTENNA__14263__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14063_ _14065_/CLK _14063_/D _12705_/Y vssd1 vssd1 vccd1 vccd1 _14063_/Q sky130_fd_sc_hd__dfrtp_2
X_11275_ _11344_/B _11344_/C _11344_/A vssd1 vssd1 vccd1 vccd1 _11345_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11516__A1 _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ _13016_/A vssd1 vssd1 vccd1 vccd1 _13014_/Y sky130_fd_sc_hd__inv_2
X_10226_ _10226_/A _10190_/A vssd1 vssd1 vccd1 vccd1 _10232_/A sky130_fd_sc_hd__or2b_1
XANTENNA_output151_A _14307_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10157_ _10157_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09192__A _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ _10126_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _10088_/X sky130_fd_sc_hd__or2_1
XFILLER_47_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13916_ _13920_/CLK _13916_/D _12328_/Y vssd1 vssd1 vccd1 vccd1 _13916_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13847_ _14198_/CLK _13847_/D _12241_/Y vssd1 vssd1 vccd1 vccd1 _13847_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13778_ _14348_/CLK _13778_/D _11975_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08999__A2 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12729_ _12753_/A vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__buf_2
XANTENNA__08255__B _08255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09940_ _10197_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _09950_/A sky130_fd_sc_hd__xnor2_2
X_09871_ _10126_/B _10083_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _09872_/B sky130_fd_sc_hd__a21oi_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07187__A1 _14097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08923__A2 _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ _08821_/A _08821_/C _08821_/B vssd1 vssd1 vccd1 vccd1 _08831_/C sky130_fd_sc_hd__a21o_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08753_ _14009_/Q _09000_/B vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07704_ _07548_/S _07651_/X _07702_/X _07619_/Y vssd1 vssd1 vccd1 vccd1 _07704_/Y
+ sky130_fd_sc_hd__a31oi_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _08684_/A vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__buf_6
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09830__A _10435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ _14128_/Q _14063_/Q vssd1 vssd1 vccd1 vccd1 _07675_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07566_ _07566_/A vssd1 vssd1 vccd1 vccd1 _14099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07350__A _14102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ _09305_/A _09305_/B vssd1 vssd1 vccd1 vccd1 _09393_/B sky130_fd_sc_hd__xnor2_2
XFILLER_107_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07497_ _14187_/Q _07452_/A vssd1 vssd1 vccd1 vccd1 _07501_/A sky130_fd_sc_hd__or2b_1
XFILLER_55_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09236_ _09236_/A _09236_/B _09236_/C vssd1 vssd1 vccd1 vccd1 _09239_/A sky130_fd_sc_hd__nand3_1
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14286__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ _08580_/B _09811_/A _09811_/B _09493_/A vssd1 vssd1 vccd1 vccd1 _09168_/C
+ sky130_fd_sc_hd__a22oi_4
XFILLER_108_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08118_ _08119_/B _08119_/C _09683_/A vssd1 vssd1 vccd1 vccd1 _08120_/A sky130_fd_sc_hd__a21oi_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _09098_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09100_/B sky130_fd_sc_hd__and2_1
XANTENNA__08181__A _09696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08049_ _08146_/A _08050_/B vssd1 vssd1 vccd1 vccd1 _08119_/C sky130_fd_sc_hd__or2_1
X_11060_ _11120_/B _11120_/C _11059_/X vssd1 vssd1 vccd1 vccd1 _11117_/C sky130_fd_sc_hd__a21bo_1
XFILLER_1_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12171__A1 _13829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11746__S _11746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _10011_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__or2b_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11962_ _11965_/A vssd1 vssd1 vccd1 vccd1 _11962_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13701_ input75/X _14454_/Q _13704_/S vssd1 vssd1 vccd1 vccd1 _13702_/B sky130_fd_sc_hd__mux2_1
X_10913_ _13909_/Q _13910_/Q _11171_/S vssd1 vssd1 vccd1 vccd1 _10913_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11893_ _13753_/Q _11893_/B vssd1 vssd1 vccd1 vccd1 _11894_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13632_ _13644_/A _13632_/B vssd1 vssd1 vccd1 vccd1 _13633_/A sky130_fd_sc_hd__and2_1
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ _10844_/A vssd1 vssd1 vccd1 vccd1 _13940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13563_ _12668_/X _14414_/Q _13576_/S vssd1 vssd1 vccd1 vccd1 _13564_/B sky130_fd_sc_hd__mux2_1
X_10775_ _10648_/A _11184_/S _10757_/B _10770_/A vssd1 vssd1 vccd1 vccd1 _10780_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12514_ _12514_/A vssd1 vssd1 vccd1 vccd1 _14008_/D sky130_fd_sc_hd__clkbuf_2
X_13494_ _12654_/X _14395_/Q _13494_/S vssd1 vssd1 vccd1 vccd1 _13495_/B sky130_fd_sc_hd__mux2_1
X_12445_ _13990_/Q _12422_/X _12444_/X _12203_/X vssd1 vssd1 vccd1 vccd1 _13990_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11510__A _11510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11737__B2 _13825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12376_ _12378_/A vssd1 vssd1 vccd1 vccd1 _12376_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08091__A _08091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ _14239_/CLK _14115_/D vssd1 vssd1 vccd1 vccd1 _14115_/Q sky130_fd_sc_hd__dfxtp_1
X_11327_ _11327_/A _11331_/A vssd1 vssd1 vccd1 vccd1 _11328_/B sky130_fd_sc_hd__or2_1
XFILLER_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10126__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14046_ _14363_/CLK _14046_/D vssd1 vssd1 vccd1 vccd1 _14046_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14009__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ _11258_/A _11258_/B vssd1 vssd1 vccd1 vccd1 _11269_/B sky130_fd_sc_hd__xnor2_2
XFILLER_84_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07169__A1 _14102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12162__A1 _13826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10209_ _10209_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10211_/B sky130_fd_sc_hd__nor2_1
X_11189_ _11240_/B _11241_/A vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__and2_1
XFILLER_95_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07435__A _07462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06993__B _14278_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13172__A _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ _14227_/Q vssd1 vssd1 vccd1 vccd1 _07442_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_78_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07351_ _14218_/Q _14220_/Q _07360_/S vssd1 vssd1 vccd1 vccd1 _07351_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07282_ _07300_/B _14166_/Q _07312_/A _07307_/C vssd1 vssd1 vccd1 vccd1 _14166_/D
+ sky130_fd_sc_hd__a31o_1
X_09021_ _09022_/A _09022_/B vssd1 vssd1 vccd1 vccd1 _09023_/B sky130_fd_sc_hd__nand2_2
XFILLER_8_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09923_ _10091_/A _10305_/B vssd1 vssd1 vccd1 vccd1 _10004_/B sky130_fd_sc_hd__xnor2_1
XFILLER_59_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__xnor2_2
XFILLER_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12251__A _12251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _08850_/A _08805_/B _08805_/C vssd1 vssd1 vccd1 vccd1 _08811_/A sky130_fd_sc_hd__nand3b_2
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _10622_/A vssd1 vssd1 vccd1 vccd1 _10634_/A sky130_fd_sc_hd__buf_2
XANTENNA__13102__A0 _12650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06997_ _06973_/X _06996_/X _14374_/Q vssd1 vssd1 vccd1 vccd1 _06998_/S sky130_fd_sc_hd__o21a_1
XFILLER_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08736_ _08731_/A _08764_/A _08731_/C _08776_/A vssd1 vssd1 vccd1 vccd1 _08740_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_96_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _08667_/A _08667_/B _08667_/C vssd1 vssd1 vccd1 vccd1 _08970_/A sky130_fd_sc_hd__nand3_1
XFILLER_96_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _14256_/Q _14254_/Q _11927_/A vssd1 vssd1 vccd1 vccd1 _07765_/S sky130_fd_sc_hd__o21a_2
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _08823_/A _09811_/B _08629_/A _08595_/A vssd1 vssd1 vccd1 vccd1 _08599_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07549_ _07549_/A vssd1 vssd1 vccd1 vccd1 _14106_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07096__B1 _07087_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ _09718_/X _09724_/A _10558_/X _10622_/A vssd1 vssd1 vccd1 vccd1 _10561_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_10_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09219_ _08580_/B _09803_/B _09811_/A _09493_/A vssd1 vssd1 vccd1 vccd1 _09220_/C
+ sky130_fd_sc_hd__a22oi_1
XFILLER_33_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10491_ _10491_/A _10491_/B _10491_/C vssd1 vssd1 vccd1 vccd1 _10492_/B sky130_fd_sc_hd__and3_1
XANTENNA__08623__B _08623_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12230_ _12517_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12231_/A sky130_fd_sc_hd__and2_1
XFILLER_2_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12161_ _12203_/A vssd1 vssd1 vccd1 vccd1 _12161_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_2_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11112_ _11125_/A _11112_/B vssd1 vssd1 vccd1 vccd1 _11112_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12092_ _13113_/B _12828_/C vssd1 vssd1 vccd1 vccd1 _12092_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11043_ _11134_/A _11134_/B vssd1 vssd1 vccd1 vccd1 _11135_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12161__A _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13691__S _13704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12994_ _12997_/A vssd1 vssd1 vccd1 vccd1 _12994_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11945_ _11947_/A vssd1 vssd1 vccd1 vccd1 _11945_/Y sky130_fd_sc_hd__inv_2
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output114_A _11829_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _13748_/Q _13747_/Q vssd1 vssd1 vccd1 vccd1 _11876_/X sky130_fd_sc_hd__and2_1
XFILLER_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ input83/X _14429_/Q _13628_/S vssd1 vssd1 vccd1 vccd1 _13616_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10827_ _10700_/X _10701_/X _10825_/X _10826_/X vssd1 vssd1 vccd1 vccd1 _13944_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12080__B1 _12021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13546_ input93/X _14409_/Q _13559_/S vssd1 vssd1 vccd1 vccd1 _13547_/B sky130_fd_sc_hd__mux2_1
XFILLER_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10758_ _10758_/A vssd1 vssd1 vccd1 vccd1 _10769_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ _13477_/A vssd1 vssd1 vccd1 vccd1 _14389_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12336__A _12348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ _13945_/Q vssd1 vssd1 vccd1 vccd1 _11533_/S sky130_fd_sc_hd__buf_2
XANTENNA__11240__A _11240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12428_ _12624_/A _12900_/A vssd1 vssd1 vccd1 vccd1 _12485_/A sky130_fd_sc_hd__nor2_2
XANTENNA__13580__A0 _12688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08252__C _09088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12359_ _12360_/A vssd1 vssd1 vccd1 vccd1 _12359_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06920_ _06917_/X _14320_/Q _06920_/S vssd1 vssd1 vccd1 vccd1 _06921_/A sky130_fd_sc_hd__mux2_1
X_14029_ _14041_/CLK _14029_/D vssd1 vssd1 vccd1 vccd1 _14029_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_110_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold16_A hold16/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09570_ _09586_/B _09586_/C _09586_/A vssd1 vssd1 vccd1 vccd1 _09570_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_64_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08521_ _09811_/A vssd1 vssd1 vccd1 vccd1 _10007_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_91_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11415__A _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08452_ _08592_/B _08452_/B _08452_/C vssd1 vssd1 vccd1 vccd1 _08590_/A sky130_fd_sc_hd__nand3_1
XFILLER_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13399__A0 _12673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07403_ _07459_/A vssd1 vssd1 vccd1 vccd1 _11746_/S sky130_fd_sc_hd__buf_2
X_08383_ _08380_/X _08381_/Y _09678_/A _08379_/Y vssd1 vssd1 vccd1 vccd1 _09698_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12071__B1 _12060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ _07321_/X _07332_/X _07333_/X _07329_/X vssd1 vssd1 vccd1 vccd1 _07334_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07265_ _13837_/Q _13836_/Q vssd1 vssd1 vccd1 vccd1 _07769_/S sky130_fd_sc_hd__nor2_1
XFILLER_118_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12246__A _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ _09072_/A _09003_/C _09000_/Y vssd1 vssd1 vccd1 vccd1 _09005_/C sky130_fd_sc_hd__a21bo_1
X_07196_ _07196_/A vssd1 vssd1 vccd1 vccd1 _14279_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07250__A0 _14263_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09790__A2 _07924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09906_ _09906_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _10065_/B sky130_fd_sc_hd__xnor2_4
XFILLER_28_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _10004_/A _09838_/A vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__or2_4
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09768_ _10578_/A _08252_/B _09764_/X _10393_/A vssd1 vssd1 vccd1 vccd1 _09769_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08719_/A _08743_/A _08719_/C vssd1 vssd1 vccd1 vccd1 _08723_/B sky130_fd_sc_hd__nand3_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09699_ _09698_/A _09698_/B _09698_/C vssd1 vssd1 vccd1 vccd1 _09699_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _13827_/Q _11730_/B vssd1 vssd1 vccd1 vccd1 _11730_/X sky130_fd_sc_hd__or2_1
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10860__A1 _11322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11661_ _11682_/C vssd1 vssd1 vccd1 vccd1 _11661_/X sky130_fd_sc_hd__clkbuf_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _13409_/A _13400_/B vssd1 vssd1 vccd1 vccd1 _13401_/A sky130_fd_sc_hd__and2_1
X_10612_ _13957_/Q _10550_/X _10606_/X _10611_/X vssd1 vssd1 vccd1 vccd1 _13957_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_23_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14380_ _14465_/CLK _14380_/D vssd1 vssd1 vccd1 vccd1 _14380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11592_ _11592_/A _11592_/B vssd1 vssd1 vccd1 vccd1 _11592_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_70_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _14348_/Q _13311_/X _13330_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _14348_/D
+ sky130_fd_sc_hd__o211a_1
X_10543_ _13965_/Q _10542_/X _10585_/S vssd1 vssd1 vccd1 vccd1 _10544_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12156__A input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input75_A io_wbs_datwr[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ _14413_/Q _13230_/X _13261_/X vssd1 vssd1 vccd1 vccd1 _13262_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ _10474_/A _10473_/A vssd1 vssd1 vccd1 vccd1 _10475_/B sky130_fd_sc_hd__or2b_1
XANTENNA__09168__C _09168_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_io_wbs_clk clkbuf_3_7_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_io_wbs_clk/X
+ sky130_fd_sc_hd__clkbuf_2
X_12213_ _12213_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _12699_/C sky130_fd_sc_hd__nor2_1
XFILLER_68_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13193_ _13193_/A vssd1 vssd1 vccd1 vccd1 _13193_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07241__A0 _14266_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ _12203_/A vssd1 vssd1 vccd1 vccd1 _12144_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12075_ _12081_/A _12075_/B vssd1 vssd1 vccd1 vccd1 _12076_/A sky130_fd_sc_hd__and2_1
XFILLER_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11026_ _11026_/A _11026_/B vssd1 vssd1 vccd1 vccd1 _11056_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12977_ _12978_/A vssd1 vssd1 vccd1 vccd1 _12977_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08528__B _09241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ input98/X vssd1 vssd1 vccd1 vccd1 _12046_/A sky130_fd_sc_hd__inv_2
XFILLER_61_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_33_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11859_ _11859_/A vssd1 vssd1 vccd1 vccd1 _11859_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13529_ _12827_/X _14404_/Q _13542_/S vssd1 vssd1 vccd1 vccd1 _13530_/B sky130_fd_sc_hd__mux2_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07050_ _14271_/Q _07046_/X _07049_/X _14367_/Q vssd1 vssd1 vccd1 vccd1 _07050_/X
+ sky130_fd_sc_hd__o211a_1
Xoutput103 _14062_/Q vssd1 vssd1 vccd1 vccd1 addr1[2] sky130_fd_sc_hd__buf_2
Xoutput114 _11829_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[10] sky130_fd_sc_hd__buf_2
XFILLER_114_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput125 _11851_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[20] sky130_fd_sc_hd__buf_2
Xoutput136 _11869_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[30] sky130_fd_sc_hd__buf_2
Xoutput147 _14303_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[11] sky130_fd_sc_hd__buf_2
XFILLER_47_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07232__A0 _14084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput158 _14313_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[21] sky130_fd_sc_hd__buf_2
Xoutput169 _14294_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[31] sky130_fd_sc_hd__buf_2
XFILLER_115_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07952_ _08312_/A vssd1 vssd1 vccd1 vccd1 _08002_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06903_ _14434_/Q _07085_/A _14466_/Q vssd1 vssd1 vccd1 vccd1 _06903_/X sky130_fd_sc_hd__and3b_1
XFILLER_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07883_ _07882_/Y _13980_/Q _07912_/S vssd1 vssd1 vccd1 vccd1 _07884_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10033__B _10090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09622_ _09622_/A _09622_/B vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09553_ _09550_/Y _09594_/A _09553_/C _09553_/D vssd1 vssd1 vccd1 vccd1 _09594_/B
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__09288__A1 _08794_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08504_ _14012_/Q vssd1 vssd1 vccd1 vccd1 _09349_/A sky130_fd_sc_hd__buf_2
X_09484_ _09478_/A _09478_/B _09478_/C vssd1 vssd1 vccd1 vccd1 _09485_/C sky130_fd_sc_hd__a21o_1
XFILLER_19_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08435_ _08435_/A _10215_/A _08592_/A _08435_/D vssd1 vssd1 vccd1 vccd1 _08592_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_93_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13360__A _13447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08366_ _08366_/A _08366_/B _09601_/A vssd1 vssd1 vccd1 vccd1 _09678_/B sky130_fd_sc_hd__nand3_2
XANTENNA__08454__A _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07317_ _07333_/S vssd1 vssd1 vccd1 vccd1 _11925_/S sky130_fd_sc_hd__inv_2
X_08297_ _09683_/A _08298_/B vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07248_ _07248_/A vssd1 vssd1 vccd1 vccd1 _14264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07179_ _14099_/Q _07167_/X _07168_/X vssd1 vssd1 vccd1 vccd1 _07179_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09285__A _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _10190_/A _10226_/A vssd1 vssd1 vccd1 vccd1 _10194_/A sky130_fd_sc_hd__xnor2_1
XFILLER_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12423__B input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12900_ _12900_/A _12900_/B vssd1 vssd1 vccd1 vccd1 _12928_/A sky130_fd_sc_hd__nor2_2
XFILLER_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13880_ _14275_/CLK _13880_/D _12283_/Y vssd1 vssd1 vccd1 vccd1 _13880_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12831_ _12831_/A vssd1 vssd1 vccd1 vccd1 _14125_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12951_/A _12762_/B _12762_/C vssd1 vssd1 vccd1 vccd1 _12828_/A sky130_fd_sc_hd__or3_4
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11713_/A vssd1 vssd1 vccd1 vccd1 _13771_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12696_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _12694_/A sky130_fd_sc_hd__and2_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14464_/CLK _14432_/D vssd1 vssd1 vccd1 vccd1 _14432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ hold30/A _11643_/Y _11652_/S vssd1 vssd1 vccd1 vccd1 _11645_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14363_ _14363_/CLK _14363_/D vssd1 vssd1 vccd1 vccd1 _14363_/Q sky130_fd_sc_hd__dfxtp_2
Xinput16 dout1[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11575_ _11541_/Y _11606_/A _11605_/B vssd1 vssd1 vccd1 vccd1 _11602_/A sky130_fd_sc_hd__o21ai_4
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput27 dout1[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
X_13314_ _14344_/Q _13311_/X _13313_/X _13301_/X vssd1 vssd1 vccd1 vccd1 _14344_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput38 io_wbs_adr[14] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
Xinput49 io_wbs_adr[24] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
X_10526_ _10597_/A _10524_/X _10525_/Y _10562_/B vssd1 vssd1 vccd1 vccd1 _10526_/X
+ sky130_fd_sc_hd__o31a_4
XFILLER_109_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14294_ _14322_/CLK _14294_/D _13159_/Y vssd1 vssd1 vccd1 vccd1 _14294_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13535__A0 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ _13245_/A vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10457_ _10457_/A _10546_/A vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__or2_1
X_13176_ _13177_/A vssd1 vssd1 vccd1 vccd1 _13176_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10388_ _10388_/A _10388_/B vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__xnor2_1
XFILLER_96_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12127_ hold31/A _12117_/X _12126_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _13814_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09923__A _10091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ _12058_/A vssd1 vssd1 vccd1 vccd1 _13798_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11009_ _13920_/Q vssd1 vssd1 vccd1 vccd1 _11010_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_77_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08220_ _08221_/B _08221_/C _08221_/A vssd1 vssd1 vccd1 vccd1 _08226_/A sky130_fd_sc_hd__a21oi_1
XFILLER_61_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08705__C _09206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08151_ _08317_/A _09786_/A _08071_/X _08150_/X vssd1 vssd1 vccd1 vccd1 _08153_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09442__A1 _09553_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09442__B2 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07102_ _14440_/Q _14264_/Q vssd1 vssd1 vccd1 vccd1 _07102_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11073__A_N _11002_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08082_ _08081_/A _08081_/B _08081_/C vssd1 vssd1 vccd1 vccd1 _08082_/Y sky130_fd_sc_hd__a21oi_1
X_07033_ _14417_/Q _07032_/Y _07009_/X vssd1 vssd1 vccd1 vccd1 _07033_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07205__A0 _14092_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08984_ _09296_/D vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__buf_2
XFILLER_114_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09833__A _10436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07935_ _13870_/Q vssd1 vssd1 vccd1 vccd1 _09123_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12501__A1 _14039_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07866_ _07919_/S vssd1 vssd1 vccd1 vccd1 _07890_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09605_ _09592_/B _09592_/Y _09603_/X _09604_/Y vssd1 vssd1 vccd1 vccd1 _09607_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07797_ _10946_/A vssd1 vssd1 vccd1 vccd1 _07798_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09536_ _09536_/A _09536_/B vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__xnor2_2
XFILLER_58_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10815__A1 _10705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ _09468_/A _09468_/B vssd1 vssd1 vccd1 vccd1 _09470_/B sky130_fd_sc_hd__or2_1
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08418_ _09881_/A vssd1 vssd1 vccd1 vccd1 _09206_/B sky130_fd_sc_hd__buf_2
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08184__A _09055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ _09329_/A _09329_/Y _09396_/Y _09397_/X vssd1 vssd1 vccd1 vccd1 _09641_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08349_ _14023_/Q vssd1 vssd1 vccd1 vccd1 _09361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11360_ _13951_/D _11536_/A vssd1 vssd1 vccd1 vccd1 _11360_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13517__A0 _12561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10311_ _10311_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10311_/Y sky130_fd_sc_hd__nor2_1
X_11291_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11292_/B sky130_fd_sc_hd__or2_1
XFILLER_106_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030_ _13115_/A vssd1 vssd1 vccd1 vccd1 _13030_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07528__A _07528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ _10120_/A _10120_/B _10120_/C vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__a21o_1
XFILLER_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10173_ _10173_/A _10173_/B vssd1 vssd1 vccd1 vccd1 _10174_/B sky130_fd_sc_hd__xnor2_1
XFILLER_65_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input38_A io_wbs_adr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13265__A _13265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13932_ _13947_/CLK _13932_/D _12347_/Y vssd1 vssd1 vccd1 vccd1 _13932_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13863_ _13867_/CLK _13863_/D _12263_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12814_ hold10/A _12801_/X _12803_/X _14145_/Q _12809_/X vssd1 vssd1 vccd1 vccd1
+ _12814_/X sky130_fd_sc_hd__a221o_1
XFILLER_90_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13794_ _14335_/CLK _13794_/D vssd1 vssd1 vccd1 vccd1 _13794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _12746_/A vssd1 vssd1 vccd1 vccd1 _12745_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12676_/A vssd1 vssd1 vccd1 vccd1 _14051_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14415_ _14449_/CLK _14415_/D vssd1 vssd1 vccd1 vccd1 _14415_/Q sky130_fd_sc_hd__dfxtp_1
X_11627_ _11627_/A _11627_/B vssd1 vssd1 vccd1 vccd1 _11627_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_8_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13220__A2 _13216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14346_ _14465_/CLK _14346_/D vssd1 vssd1 vccd1 vccd1 _14346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11558_ _14044_/Q _13956_/Q vssd1 vssd1 vccd1 vccd1 _11638_/A sky130_fd_sc_hd__and2_1
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13508__A0 _12673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10509_ _10520_/B _10501_/Y _10506_/Y _10508_/X vssd1 vssd1 vccd1 vccd1 _10511_/B
+ sky130_fd_sc_hd__o211ai_1
X_14277_ _14281_/CLK _14277_/D _13138_/Y vssd1 vssd1 vccd1 vccd1 _14277_/Q sky130_fd_sc_hd__dfrtp_4
X_11489_ _11513_/A vssd1 vssd1 vccd1 vccd1 _11489_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _13254_/A vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13159_/A vssd1 vssd1 vccd1 vccd1 _13159_/Y sky130_fd_sc_hd__inv_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07720_ _07730_/S vssd1 vssd1 vccd1 vccd1 _07720_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08269__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07651_ _14075_/Q _07651_/B vssd1 vssd1 vccd1 vccd1 _07651_/X sky130_fd_sc_hd__xor2_2
XFILLER_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07582_ _14091_/Q input7/X _07582_/S vssd1 vssd1 vccd1 vccd1 _07583_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ _09346_/A _09321_/B _09321_/C vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__nand3_1
XFILLER_34_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12519__A _12536_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08716__B _08716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _09333_/B _09252_/B vssd1 vssd1 vccd1 vccd1 _09276_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11470__A1 _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08203_ _08213_/B _08203_/B _08203_/C vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__or3_2
XANTENNA__11142__B _11142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09183_ _09180_/Y _09181_/X _09106_/C _09106_/Y vssd1 vssd1 vccd1 vccd1 _09184_/C
+ sky130_fd_sc_hd__a211o_1
X_08134_ _08208_/B _09963_/B _08132_/D _08249_/A vssd1 vssd1 vccd1 vccd1 _08134_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_107_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08065_ _08135_/A _08289_/A _08140_/A _08061_/Y vssd1 vssd1 vccd1 vccd1 _08066_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_108_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07016_ _07016_/A vssd1 vssd1 vccd1 vccd1 _14308_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07729__A1 _14159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07067__B _07098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08967_ _08967_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _08967_/X sky130_fd_sc_hd__or2b_1
XFILLER_5_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07918_ _07918_/A _07918_/B vssd1 vssd1 vccd1 vccd1 _07918_/X sky130_fd_sc_hd__xor2_1
XFILLER_69_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08898_ _08934_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08921_/A sky130_fd_sc_hd__nor2_1
XFILLER_5_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08179__A _09402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07849_ _14033_/Q _13979_/Q vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__and2_1
XFILLER_95_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10860_ _11322_/A _10853_/C _10858_/X _10859_/Y vssd1 vssd1 vccd1 vccd1 _10860_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__12789__A1 _14112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09519_ _09518_/A _09518_/C _09518_/B vssd1 vssd1 vccd1 vccd1 _09519_/X sky130_fd_sc_hd__a21o_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _13931_/Q _10791_/B vssd1 vssd1 vccd1 vccd1 _10792_/B sky130_fd_sc_hd__or2_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12530_ _12917_/A _08983_/B _12537_/S vssd1 vssd1 vccd1 vccd1 _12531_/B sky130_fd_sc_hd__mux2_1
XFILLER_13_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12461_ _08983_/B _12439_/X _12454_/X _14045_/Q vssd1 vssd1 vccd1 vccd1 _12461_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14200_ _14215_/CLK _14200_/D _12991_/Y vssd1 vssd1 vccd1 vccd1 _14200_/Q sky130_fd_sc_hd__dfrtp_1
X_11412_ _11529_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11525_/A sky130_fd_sc_hd__or2_1
XANTENNA__08064__D _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11987__B input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ _12410_/A vssd1 vssd1 vccd1 vccd1 _12397_/A sky130_fd_sc_hd__buf_2
X_14131_ _14250_/CLK _14131_/D vssd1 vssd1 vccd1 vccd1 _14131_/Q sky130_fd_sc_hd__dfxtp_1
X_11343_ _11276_/A _10904_/X _11342_/Y _07784_/X vssd1 vssd1 vccd1 vccd1 _13899_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08090__B1 _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09457__B _09457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12164__A _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14062_ _14065_/CLK _14062_/D _12703_/Y vssd1 vssd1 vccd1 vccd1 _14062_/Q sky130_fd_sc_hd__dfrtp_2
X_11274_ _11341_/B _11274_/B vssd1 vssd1 vccd1 vccd1 _11344_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13694__S _13704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13013_ _13016_/A vssd1 vssd1 vccd1 vccd1 _13013_/Y sky130_fd_sc_hd__inv_2
X_10225_ _10279_/B _10225_/B vssd1 vssd1 vccd1 vccd1 _10236_/A sky130_fd_sc_hd__xnor2_2
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09473__A _14021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ _10156_/A _10171_/B vssd1 vssd1 vccd1 vccd1 _10172_/A sky130_fd_sc_hd__nand2_1
XANTENNA_output144_A _11827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__buf_2
X_10087_ _10126_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _10087_/X sky130_fd_sc_hd__and2_1
XFILLER_43_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13915_ _13915_/CLK _13915_/D _12327_/Y vssd1 vssd1 vccd1 vccd1 _13915_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_69_io_wbs_clk clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14163_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__12229__A0 _12906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13846_ _14028_/CLK _13846_/D _12239_/Y vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfrtp_1
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13777_ _14348_/CLK _13777_/D _11974_/Y vssd1 vssd1 vccd1 vccd1 _13777_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_16_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10989_ _13925_/Q vssd1 vssd1 vccd1 vccd1 _11082_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12728_ _13010_/A vssd1 vssd1 vccd1 vccd1 _12753_/A sky130_fd_sc_hd__clkbuf_2
X_12659_ _13072_/A vssd1 vssd1 vccd1 vccd1 _12678_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08552__A _08716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14329_ _14396_/CLK _14329_/D vssd1 vssd1 vccd1 vccd1 _14329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09870_ _09870_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _10092_/B sky130_fd_sc_hd__xnor2_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08821_/A _08821_/B _08821_/C vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__nand3_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08758_/A _08758_/C _08758_/B vssd1 vssd1 vccd1 vccd1 _08785_/B sky130_fd_sc_hd__a21o_1
XFILLER_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07703_ _14148_/Q _07548_/S _07702_/X hold37/X vssd1 vssd1 vccd1 vccd1 _07703_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_39_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08683_ _08937_/B vssd1 vssd1 vccd1 vccd1 _08683_/X sky130_fd_sc_hd__buf_8
XFILLER_54_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07634_ _07628_/Y _07679_/A _07678_/B vssd1 vssd1 vccd1 vccd1 _07676_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07565_ _14099_/Q input16/X _07571_/S vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12249__A _12251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09304_ _09304_/A _09303_/X vssd1 vssd1 vccd1 vccd1 _09305_/B sky130_fd_sc_hd__or2b_1
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07496_ _14189_/Q _07495_/X _07493_/X vssd1 vssd1 vccd1 vccd1 _14189_/D sky130_fd_sc_hd__a21bo_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09235_ _09233_/B _09553_/D _09058_/B _09508_/A vssd1 vssd1 vccd1 vccd1 _09236_/C
+ sky130_fd_sc_hd__a22o_1
X_09166_ _09297_/A _09875_/A vssd1 vssd1 vccd1 vccd1 _09168_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08117_ _09590_/A vssd1 vssd1 vccd1 vccd1 _09683_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09097_ _09097_/A _09097_/B _09097_/C vssd1 vssd1 vccd1 vccd1 _09100_/A sky130_fd_sc_hd__nand3_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08048_ _08295_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08050_/B sky130_fd_sc_hd__xnor2_1
XFILLER_116_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10010_ _09895_/A _10127_/A _10048_/B _10048_/A vssd1 vssd1 vccd1 vccd1 _10397_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09999_ _09999_/A _09999_/B vssd1 vssd1 vccd1 vccd1 _09999_/Y sky130_fd_sc_hd__nand2_2
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11961_ _11965_/A vssd1 vssd1 vccd1 vccd1 _11961_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13700_ _13700_/A vssd1 vssd1 vccd1 vccd1 _14453_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10912_ _10912_/A vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__buf_2
XFILLER_45_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11892_ _13812_/Q _11882_/X _11890_/X _11891_/Y _11885_/X vssd1 vssd1 vccd1 vccd1
+ _13752_/D sky130_fd_sc_hd__o221a_1
XFILLER_45_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13631_ input89/X _14434_/Q _13634_/S vssd1 vssd1 vccd1 vccd1 _13632_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10843_ _13940_/Q _10842_/X _10871_/S vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09627__A1 _09360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12159__A input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11434__A1 _11007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13562_ _13634_/S vssd1 vssd1 vccd1 vccd1 _13576_/S sky130_fd_sc_hd__clkbuf_2
X_10774_ _13931_/Q _10791_/B vssd1 vssd1 vccd1 vccd1 _10884_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12513_ _12517_/A _12513_/B vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__and2_1
XANTENNA__11998__A _12008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13493_ _13493_/A vssd1 vssd1 vccd1 vccd1 _14394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ _14025_/Q _12438_/X _12443_/X _12435_/X vssd1 vssd1 vccd1 vccd1 _12444_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12375_ _12378_/A vssd1 vssd1 vccd1 vccd1 _12375_/Y sky130_fd_sc_hd__inv_2
X_14114_ _14250_/CLK _14114_/D vssd1 vssd1 vccd1 vccd1 _14114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_99_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11326_ _11294_/A _11319_/X _11325_/Y _11322_/X vssd1 vssd1 vccd1 vccd1 _13905_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14045_ _14363_/CLK _14045_/D vssd1 vssd1 vccd1 vccd1 _14045_/Q sky130_fd_sc_hd__dfxtp_1
X_11257_ _11355_/B _11262_/C _11252_/A vssd1 vssd1 vccd1 vccd1 _11258_/B sky130_fd_sc_hd__a21oi_1
XFILLER_69_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10208_ _10208_/A _10208_/B _10208_/C vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__and3_1
XFILLER_68_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11188_ _11142_/A _11185_/X _11187_/X vssd1 vssd1 vccd1 vccd1 _11241_/A sky130_fd_sc_hd__o21ai_2
XFILLER_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10139_ _10139_/A _10139_/B vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__xnor2_1
XFILLER_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09931__A _10090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13829_ _14335_/CLK _13829_/D vssd1 vssd1 vccd1 vccd1 _13829_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11425__A1 _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ _14102_/Q _07336_/X vssd1 vssd1 vccd1 vccd1 _07350_/X sky130_fd_sc_hd__or2b_1
X_07281_ _07274_/A _07312_/B _07307_/A vssd1 vssd1 vccd1 vccd1 _14165_/D sky130_fd_sc_hd__a21o_1
X_09020_ _09071_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09022_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08282__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12925__A1 _14157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12689__A0 _12688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09922_ _10091_/A vssd1 vssd1 vccd1 vccd1 _09922_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_53_io_wbs_clk_A clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09853_ _09959_/A _09959_/B vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__xnor2_2
XFILLER_113_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08804_ _08774_/B _08762_/C _08762_/A vssd1 vssd1 vccd1 vccd1 _08805_/B sky130_fd_sc_hd__o21ai_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _10578_/A vssd1 vssd1 vccd1 vccd1 _10622_/A sky130_fd_sc_hd__clkbuf_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06996_ _14422_/Q _07020_/B _14454_/Q vssd1 vssd1 vccd1 vccd1 _06996_/X sky130_fd_sc_hd__and3b_1
XFILLER_26_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08735_ _08735_/A _08735_/B _08735_/C vssd1 vssd1 vccd1 vccd1 _08776_/A sky130_fd_sc_hd__and3_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08666_ _08665_/A _08665_/B _08665_/C vssd1 vssd1 vccd1 vccd1 _08667_/C sky130_fd_sc_hd__a21o_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08457__A _08796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ hold12/A _14254_/Q vssd1 vssd1 vccd1 vccd1 _11927_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08597_ _09207_/C vssd1 vssd1 vccd1 vccd1 _08629_/A sky130_fd_sc_hd__buf_2
XFILLER_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11416__A1 _11032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07548_ _14106_/Q input24/X _07548_/S vssd1 vssd1 vccd1 vccd1 _07549_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07479_ _07483_/A _07479_/B vssd1 vssd1 vccd1 vccd1 _07479_/X sky130_fd_sc_hd__or2_1
XFILLER_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09218_ _09491_/A _09218_/B vssd1 vssd1 vccd1 vccd1 _09220_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08192__A _08403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10490_ _10491_/A _10491_/B _10491_/C vssd1 vssd1 vccd1 vccd1 _10492_/A sky130_fd_sc_hd__a21oi_1
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09149_ _09148_/A _09148_/C _09148_/B vssd1 vssd1 vccd1 vccd1 _09151_/B sky130_fd_sc_hd__o21ai_2
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ _12911_/A _12160_/B vssd1 vssd1 vccd1 vccd1 _12160_/X sky130_fd_sc_hd__or2_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11111_ _11111_/A _11111_/B _11115_/B vssd1 vssd1 vccd1 vccd1 _11111_/X sky130_fd_sc_hd__or3_1
X_12091_ _12823_/C vssd1 vssd1 vccd1 vccd1 _12828_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_1_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11042_ _13911_/Q vssd1 vssd1 vccd1 vccd1 _11134_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11058__A _11058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input20_A dout1[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12993_ _12997_/A vssd1 vssd1 vccd1 vccd1 _12993_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11944_ _11947_/A vssd1 vssd1 vccd1 vccd1 _11944_/Y sky130_fd_sc_hd__inv_2
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08367__A _08716_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11875_ hold24/X _11872_/X _11873_/Y _11874_/X vssd1 vssd1 vccd1 vccd1 _13747_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13614_ _13614_/A vssd1 vssd1 vccd1 vccd1 _13628_/S sky130_fd_sc_hd__buf_2
XANTENNA__12604__A0 _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10826_ _10826_/A vssd1 vssd1 vccd1 vccd1 _10826_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13545_ _13634_/S vssd1 vssd1 vccd1 vccd1 _13559_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10757_ _11184_/S _10757_/B vssd1 vssd1 vccd1 vccd1 _10757_/X sky130_fd_sc_hd__or2_1
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ _13485_/A _13476_/B vssd1 vssd1 vccd1 vccd1 _13477_/A sky130_fd_sc_hd__and2_1
XFILLER_51_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ _10688_/A vssd1 vssd1 vccd1 vccd1 _13946_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13770__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12427_ _12624_/A _13079_/A vssd1 vssd1 vccd1 vccd1 _12486_/A sky130_fd_sc_hd__nor2_2
XFILLER_12_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09348__D _13872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ _12360_/A vssd1 vssd1 vccd1 vccd1 _12358_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11309_ _11309_/A _11309_/B vssd1 vssd1 vccd1 vccd1 _11309_/X sky130_fd_sc_hd__xor2_1
XFILLER_99_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12289_ _12291_/A vssd1 vssd1 vccd1 vccd1 _12289_/Y sky130_fd_sc_hd__inv_2
X_14028_ _14028_/CLK _14028_/D vssd1 vssd1 vccd1 vccd1 _14028_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07011__A1 _14276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13096__A0 _12641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08520_ _08828_/B vssd1 vssd1 vccd1 vccd1 _08978_/B sky130_fd_sc_hd__buf_4
XANTENNA__12843__A0 _12641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08451_ _08435_/A _10215_/A _08592_/A _08435_/D vssd1 vssd1 vccd1 vccd1 _08452_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ _07528_/A _07402_/B vssd1 vssd1 vccd1 vccd1 _07402_/X sky130_fd_sc_hd__or2_1
XANTENNA__08427__D _09091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08382_ _09678_/A _08379_/Y _08380_/X _08381_/Y vssd1 vssd1 vccd1 vccd1 _09698_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_91_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07333_ _14221_/Q _14223_/Q _07333_/S vssd1 vssd1 vccd1 vccd1 _07333_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07264_ _14058_/Q _07459_/A vssd1 vssd1 vccd1 vccd1 _07264_/Y sky130_fd_sc_hd__nand2_1
X_09003_ _09000_/Y _09072_/A _09003_/C vssd1 vssd1 vccd1 vccd1 _09072_/B sky130_fd_sc_hd__nand3b_1
XFILLER_118_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07195_ _14279_/Q _07194_/X _07201_/S vssd1 vssd1 vccd1 vccd1 _07196_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12262__A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09905_ _09905_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__xor2_2
XFILLER_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07002__A1 _14277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _09824_/A _09857_/A _09835_/X vssd1 vssd1 vccd1 vccd1 _09838_/A sky130_fd_sc_hd__o21a_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06979_ _14424_/Q _06978_/Y _06970_/X vssd1 vssd1 vccd1 vccd1 _06979_/X sky130_fd_sc_hd__a21o_1
X_09767_ _10367_/A vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _08719_/A _08719_/C _08743_/A vssd1 vssd1 vccd1 vccd1 _08723_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12834__A0 _12515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _09698_/A _09698_/B _09698_/C vssd1 vssd1 vccd1 vccd1 _09698_/X sky130_fd_sc_hd__or3_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08187__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _09804_/A vssd1 vssd1 vccd1 vccd1 _08836_/B sky130_fd_sc_hd__buf_6
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _13773_/Q _13771_/Q vssd1 vssd1 vccd1 vccd1 _11682_/C sky130_fd_sc_hd__and2b_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13793__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07069__A1 _14301_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10611_ _10634_/A _10610_/Y _09788_/X vssd1 vssd1 vccd1 vccd1 _10611_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11591_ _11591_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11592_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13330_ _14428_/Q _13327_/X _13329_/X _13320_/X vssd1 vssd1 vccd1 vccd1 _13330_/X
+ sky130_fd_sc_hd__a211o_1
X_10542_ _10537_/Y _10538_/X _10541_/Y _10528_/X vssd1 vssd1 vccd1 vccd1 _10542_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13261_ _14445_/Q _13250_/X _13245_/X _14397_/Q vssd1 vssd1 vccd1 vccd1 _13261_/X
+ sky130_fd_sc_hd__a22o_1
X_10473_ _10473_/A _10474_/A vssd1 vssd1 vccd1 vccd1 _10498_/B sky130_fd_sc_hd__or2b_1
XFILLER_108_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ _13358_/A vssd1 vssd1 vccd1 vccd1 _13059_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11995__B _12211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ _13193_/A vssd1 vssd1 vccd1 vccd1 _13192_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input68_A io_wbs_datwr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ input80/X _12143_/B vssd1 vssd1 vccd1 vccd1 _12143_/X sky130_fd_sc_hd__or2_1
XANTENNA__12770__C1 _12498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12172__A input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07266__A _13951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ _13803_/Q _12059_/X _12060_/X _13819_/Q vssd1 vssd1 vccd1 vccd1 _12075_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07529__C1 _14192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11025_ _11244_/A _11029_/A _11029_/B vssd1 vssd1 vccd1 vccd1 _11026_/B sky130_fd_sc_hd__a21oi_1
XFILLER_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12900__A _12900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11628__A1 _11627_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12825__B1 _11745_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ _12978_/A vssd1 vssd1 vccd1 vccd1 _12976_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08097__A _08789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08528__C _09074_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11927_ _11927_/A vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__inv_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13731__A _13731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11858_ _14349_/Q _11864_/B vssd1 vssd1 vccd1 vccd1 _11859_/A sky130_fd_sc_hd__and2_1
XFILLER_14_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12053__A1 _13797_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ _13937_/Q _10809_/B vssd1 vssd1 vccd1 vccd1 _10810_/B sky130_fd_sc_hd__nor2_1
X_11789_ _14325_/Q _13194_/A _12192_/A _13834_/Q _11788_/X vssd1 vssd1 vccd1 vccd1
+ _11790_/B sky130_fd_sc_hd__a221o_1
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13528_ _13634_/S vssd1 vssd1 vccd1 vccd1 _13542_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10603__A2 _10613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07480__A1 _14078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13459_ _13459_/A vssd1 vssd1 vccd1 vccd1 _14384_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_115_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput104 _14063_/Q vssd1 vssd1 vccd1 vccd1 addr1[3] sky130_fd_sc_hd__buf_2
Xoutput115 _11832_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[11] sky130_fd_sc_hd__buf_2
XFILLER_86_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput126 _11852_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[21] sky130_fd_sc_hd__buf_2
Xoutput137 _11871_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[31] sky130_fd_sc_hd__buf_2
XANTENNA__13178__A _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput148 _14304_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[12] sky130_fd_sc_hd__buf_2
Xoutput159 _14314_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[22] sky130_fd_sc_hd__buf_2
XFILLER_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07951_ _09362_/A vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__buf_2
XFILLER_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11316__B1 _10851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06902_ _14290_/Q _06873_/X _06901_/X _14386_/Q vssd1 vssd1 vccd1 vccd1 _06902_/X
+ sky130_fd_sc_hd__o211a_1
X_07882_ _07882_/A _07882_/B vssd1 vssd1 vccd1 vccd1 _07882_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_96_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13069__A0 _12579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09621_ _09575_/X _09578_/Y _09576_/X _09577_/X vssd1 vssd1 vccd1 vccd1 _09622_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10031__A1_N _10421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ _09152_/A _09233_/C _09550_/Y _09594_/A vssd1 vssd1 vccd1 vccd1 _09554_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_71_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08503_ _08503_/A _08503_/B _08503_/C vssd1 vssd1 vccd1 vccd1 _08517_/A sky130_fd_sc_hd__nand3_1
XFILLER_93_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09483_ _09483_/A _09483_/B vssd1 vssd1 vccd1 vccd1 _09485_/B sky130_fd_sc_hd__xor2_1
XFILLER_102_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08434_ _08449_/B _09873_/A _08449_/C _09233_/A vssd1 vssd1 vccd1 vccd1 _08435_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13641__A _13644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08365_ _08366_/B _09601_/A _08366_/A vssd1 vssd1 vccd1 vccd1 _09678_/A sky130_fd_sc_hd__a21o_2
XANTENNA__08248__B1 _08208_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12257__A _12259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ _07348_/A vssd1 vssd1 vccd1 vccd1 _07316_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08296_ _08323_/A _08323_/B _08295_/Y vssd1 vssd1 vccd1 vccd1 _08298_/B sky130_fd_sc_hd__o21a_1
XFILLER_109_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07247_ _14264_/Q _07246_/X _07253_/S vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__mux2_1
X_07178_ _07178_/A vssd1 vssd1 vccd1 vccd1 _14284_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__B _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12504__C1 _12498_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12720__A _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09819_ _09233_/C _09857_/B _09818_/X vssd1 vssd1 vccd1 vccd1 _09826_/A sky130_fd_sc_hd__a21oi_1
XFILLER_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ _13184_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _12831_/A sky130_fd_sc_hd__or2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12429_/A _11988_/A _12773_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _12761_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11712_ _11715_/A _11714_/A _13771_/Q vssd1 vssd1 vccd1 vccd1 _11713_/A sky130_fd_sc_hd__mux2_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ input73/X _14056_/Q _12695_/S vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__mux2_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _14464_/CLK _14431_/D vssd1 vssd1 vccd1 vccd1 _14431_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11643_/A _11643_/B vssd1 vssd1 vccd1 vccd1 _11643_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12167__A _12917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14362_ _14410_/CLK _14362_/D vssd1 vssd1 vccd1 vccd1 _14362_/Q sky130_fd_sc_hd__dfxtp_2
X_11574_ _14052_/Q _13964_/Q vssd1 vssd1 vccd1 vccd1 _11605_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 dout1[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
XFILLER_11_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput28 dout1[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_1
Xinput39 io_wbs_adr[15] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
X_13313_ _14424_/Q _13306_/X _13312_/X _13299_/X vssd1 vssd1 vccd1 vccd1 _13313_/X
+ sky130_fd_sc_hd__a211o_1
X_10525_ _10524_/A _10524_/B _10524_/C vssd1 vssd1 vccd1 vccd1 _10525_/Y sky130_fd_sc_hd__a21oi_1
X_14293_ _14322_/CLK _14293_/D _13158_/Y vssd1 vssd1 vccd1 vccd1 _14293_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13244_ _14329_/Q _13240_/X _13243_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _14329_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10456_ _10456_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10546_/A sky130_fd_sc_hd__nand2_1
XANTENNA_output174_A _14299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__D1 _08944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ _13177_/A vssd1 vssd1 vccd1 vccd1 _13175_/Y sky130_fd_sc_hd__inv_2
X_10387_ _09801_/A _10421_/B _09801_/B vssd1 vssd1 vccd1 vccd1 _10388_/B sky130_fd_sc_hd__a21boi_1
XFILLER_112_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _12942_/A _12130_/B vssd1 vssd1 vccd1 vccd1 _12126_/X sky130_fd_sc_hd__or2_1
XFILLER_111_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12057_ _12065_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _12058_/A sky130_fd_sc_hd__and2_1
XFILLER_42_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09923__B _10305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11008_ _11008_/A _11008_/B vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__xor2_1
XFILLER_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12959_ _12960_/A vssd1 vssd1 vccd1 vccd1 _12959_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08150_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08150_/X sky130_fd_sc_hd__and2_1
XFILLER_105_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08705__D _09873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09442__A2 _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07101_ _07101_/A vssd1 vssd1 vccd1 vccd1 _14297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ _08081_/A _08081_/B _08081_/C vssd1 vssd1 vccd1 vccd1 _08160_/C sky130_fd_sc_hd__and3_1
XFILLER_88_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12805__A _12817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07032_ _14449_/Q _14273_/Q vssd1 vssd1 vccd1 vccd1 _07032_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _08983_/A _08983_/B _08983_/C _10007_/A vssd1 vssd1 vccd1 vccd1 _08986_/B
+ sky130_fd_sc_hd__nand4_4
XFILLER_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ _09145_/B vssd1 vssd1 vccd1 vccd1 _09084_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12540__A _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ _07858_/Y _07868_/B _07857_/Y _07874_/S vssd1 vssd1 vccd1 vccd1 _07865_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_84_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09604_ _09676_/B _09676_/C _09676_/A vssd1 vssd1 vccd1 vccd1 _09604_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_113_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07796_ _13948_/Q vssd1 vssd1 vccd1 vccd1 _10946_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09535_ _09535_/A _09535_/B vssd1 vssd1 vccd1 vccd1 _09536_/B sky130_fd_sc_hd__or2_1
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09466_ _09522_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09468_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08417_ _13866_/Q vssd1 vssd1 vccd1 vccd1 _09881_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12017__B2 _13828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09397_ _09396_/C _09396_/B _09360_/Y vssd1 vssd1 vccd1 vccd1 _09397_/X sky130_fd_sc_hd__a21bo_2
XFILLER_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08348_ _14021_/Q _09479_/D vssd1 vssd1 vccd1 vccd1 _09555_/C sky130_fd_sc_hd__and2_1
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10579__A1 _10644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08279_ _09777_/A _08233_/B _08278_/X vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__o21a_1
XFILLER_4_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10310_ _10310_/A _10310_/B vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11290_ _11330_/B _11334_/A _11330_/A vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__a21oi_1
XFILLER_118_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10241_ _10638_/B _10636_/A vssd1 vssd1 vccd1 vccd1 _10241_/X sky130_fd_sc_hd__or2_1
XFILLER_106_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10172_ _10172_/A _10172_/B vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__nand2_2
XFILLER_65_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13931_ _13982_/CLK _13931_/D _12346_/Y vssd1 vssd1 vccd1 vccd1 _13931_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_59_io_wbs_clk clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14411_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13862_ _13897_/CLK _13862_/D _12259_/Y vssd1 vssd1 vccd1 vccd1 _13862_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_75_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12813_ _14119_/Q _12800_/X _12812_/X _12805_/X vssd1 vssd1 vccd1 vccd1 _14119_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13793_ _14335_/CLK _13793_/D vssd1 vssd1 vccd1 vccd1 _13793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12746_/A vssd1 vssd1 vccd1 vccd1 _12744_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07132__B1 _06970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12678_/A _12675_/B vssd1 vssd1 vccd1 vccd1 _12676_/A sky130_fd_sc_hd__and2_1
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14414_ _14449_/CLK _14414_/D vssd1 vssd1 vccd1 vccd1 _14414_/Q sky130_fd_sc_hd__dfxtp_1
X_11626_ _11545_/Y _11626_/B vssd1 vssd1 vccd1 vccd1 _11627_/B sky130_fd_sc_hd__and2b_1
XFILLER_11_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14345_ _14348_/CLK _14345_/D vssd1 vssd1 vccd1 vccd1 _14345_/Q sky130_fd_sc_hd__dfxtp_1
X_11557_ _14043_/Q _13955_/Q _11556_/X vssd1 vssd1 vccd1 vccd1 _11639_/B sky130_fd_sc_hd__o21a_1
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10508_ _10508_/A _10508_/B vssd1 vssd1 vccd1 vccd1 _10508_/X sky130_fd_sc_hd__or2_1
X_11488_ _11482_/A _11487_/X _10686_/X vssd1 vssd1 vccd1 vccd1 _11488_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14276_ _14281_/CLK _14276_/D _13137_/Y vssd1 vssd1 vccd1 vccd1 _14276_/Q sky130_fd_sc_hd__dfrtp_4
X_13227_ _14358_/Q _13215_/X _13226_/X _13222_/X vssd1 vssd1 vccd1 vccd1 _13227_/X
+ sky130_fd_sc_hd__a211o_1
X_10439_ _10439_/A _10439_/B vssd1 vssd1 vccd1 vccd1 _10472_/S sky130_fd_sc_hd__nor2_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13158_ _13159_/A vssd1 vssd1 vccd1 vccd1 _13158_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12932_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12109_/X sky130_fd_sc_hd__or2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13089_ _13089_/A _13089_/B vssd1 vssd1 vccd1 vccd1 _13090_/A sky130_fd_sc_hd__and2_1
XANTENNA__12360__A _12360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_58_io_wbs_clk_A clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07650_ _14074_/Q _07656_/A vssd1 vssd1 vccd1 vccd1 _07651_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07581_ _07581_/A vssd1 vssd1 vccd1 vccd1 _14092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13191__A _13193_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ _09316_/A _09316_/B _09316_/C vssd1 vssd1 vccd1 vccd1 _09321_/C sky130_fd_sc_hd__a21o_1
XFILLER_81_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08285__A _09001_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08716__C _08925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09251_ _09248_/X _09249_/Y _09137_/A _09140_/A vssd1 vssd1 vccd1 vccd1 _09252_/B
+ sky130_fd_sc_hd__o211ai_1
X_08202_ _08243_/C _08202_/B vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__nand2_2
X_09182_ _09106_/C _09106_/Y _09180_/Y _09181_/X vssd1 vssd1 vccd1 vccd1 _09184_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08133_ _09822_/A vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_105_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08064_ _08140_/A _08061_/Y _08135_/A _09822_/A vssd1 vssd1 vccd1 vccd1 _08140_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07015_ _07011_/X _14308_/Q _07015_/S vssd1 vssd1 vccd1 vccd1 _07016_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09844__A _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08966_ _08966_/A _10486_/S _08966_/C vssd1 vssd1 vccd1 vccd1 _08966_/X sky130_fd_sc_hd__and3_1
XFILLER_103_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07364__A _14099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07917_ _07917_/A vssd1 vssd1 vccd1 vccd1 _13972_/D sky130_fd_sc_hd__clkbuf_1
X_08897_ _08897_/A _08897_/B vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__xnor2_1
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07848_ _07848_/A _07848_/B vssd1 vssd1 vccd1 vccd1 _07886_/B sky130_fd_sc_hd__and2_1
XFILLER_112_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07779_ _07779_/A _11585_/S _10585_/S vssd1 vssd1 vccd1 vccd1 _07780_/A sky130_fd_sc_hd__or3_1
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09518_ _09518_/A _09518_/B _09518_/C vssd1 vssd1 vccd1 vccd1 _09518_/Y sky130_fd_sc_hd__nand3_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10790_ _10894_/A _10894_/B _10894_/C vssd1 vssd1 vccd1 vccd1 _10889_/C sky130_fd_sc_hd__a21oi_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07114__B1 _14359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_60_io_wbs_clk_A clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09449_ _09449_/A _09448_/X vssd1 vssd1 vccd1 vccd1 _09450_/B sky130_fd_sc_hd__or2b_1
XANTENNA__08862__B1 _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12460_ _12460_/A vssd1 vssd1 vccd1 vccd1 _12460_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11411_ _13895_/Q _11048_/A _11415_/A vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__mux2_1
X_12391_ _12391_/A vssd1 vssd1 vccd1 vccd1 _12391_/Y sky130_fd_sc_hd__inv_2
X_11342_ _11342_/A _11342_/B vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__nor2_1
X_14130_ _14152_/CLK _14130_/D vssd1 vssd1 vccd1 vccd1 _14130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09457__C _13874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11273_ _11273_/A _11273_/B vssd1 vssd1 vccd1 vccd1 _11274_/B sky130_fd_sc_hd__or2_1
XFILLER_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14061_ _14065_/CLK _14061_/D _12702_/Y vssd1 vssd1 vccd1 vccd1 _14061_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08917__A1 _08683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _10213_/Y _10221_/X _10222_/Y _10223_/Y vssd1 vssd1 vccd1 vccd1 _10224_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_106_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input50_A io_wbs_adr[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13012_ _13016_/A vssd1 vssd1 vccd1 vccd1 _13012_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10155_ _10182_/A vssd1 vssd1 vccd1 vccd1 _10155_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10086_ _10138_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _10086_/X sky130_fd_sc_hd__or2_1
XFILLER_94_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13674__A0 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12477__A1 _08632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13914_ _13915_/CLK _13914_/D _12326_/Y vssd1 vssd1 vccd1 vccd1 _13914_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _14028_/CLK _13845_/D _12238_/Y vssd1 vssd1 vccd1 vccd1 _13845_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13776_ _14348_/CLK _13776_/D _11973_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Q sky130_fd_sc_hd__dfrtp_2
X_10988_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11093_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _12727_/A vssd1 vssd1 vccd1 vccd1 _12727_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12658_ _13428_/A vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__buf_4
XFILLER_102_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11609_ _11609_/A _11609_/B vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12589_ _12589_/A vssd1 vssd1 vccd1 vccd1 _14029_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12355__A _12379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14328_ _14396_/CLK _14328_/D vssd1 vssd1 vccd1 vccd1 _14328_/Q sky130_fd_sc_hd__dfxtp_1
X_14259_ _14259_/CLK _14259_/D _13115_/Y vssd1 vssd1 vccd1 vccd1 _14259_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08820_/A _08820_/B _08820_/C vssd1 vssd1 vccd1 vccd1 _08834_/A sky130_fd_sc_hd__nand3_1
XFILLER_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12090__A _12211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08751_ _08787_/B _08787_/C _08787_/A vssd1 vssd1 vccd1 vccd1 _08758_/B sky130_fd_sc_hd__o21bai_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07702_ _14147_/Q _07706_/A _07651_/X _14148_/Q _07701_/X vssd1 vssd1 vccd1 vccd1
+ _07702_/X sky130_fd_sc_hd__a221o_2
XFILLER_39_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08682_ _08682_/A _08610_/B vssd1 vssd1 vccd1 vccd1 _08687_/B sky130_fd_sc_hd__or2b_1
XFILLER_94_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07633_ _14127_/Q _14062_/Q vssd1 vssd1 vccd1 vccd1 _07678_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07564_ _07564_/A vssd1 vssd1 vccd1 vccd1 _14100_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_0_0_io_wbs_clk clkbuf_2_1_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_io_wbs_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09303_ _09302_/A _09302_/C _09302_/B vssd1 vssd1 vccd1 vccd1 _09303_/X sky130_fd_sc_hd__a21o_1
XFILLER_110_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07495_ _14188_/Q _14187_/Q _07452_/A vssd1 vssd1 vccd1 vccd1 _07495_/X sky130_fd_sc_hd__or3b_1
XFILLER_16_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _09234_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__and2_1
XFILLER_22_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09165_ _09165_/A _09217_/B _09165_/C _09881_/A vssd1 vssd1 vccd1 vccd1 _09216_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08116_ _09465_/A _08116_/B vssd1 vssd1 vccd1 vccd1 _09590_/A sky130_fd_sc_hd__xor2_4
XANTENNA__12943__A2 _12928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__A _14100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09096_ _09090_/A _09090_/C _09090_/B vssd1 vssd1 vccd1 vccd1 _09097_/C sky130_fd_sc_hd__a21o_1
XANTENNA__08072__A1 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08047_ _08622_/A _09800_/A _07994_/A _07985_/B vssd1 vssd1 vccd1 vccd1 _08115_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07078__B _14267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14182__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14470__182 vssd1 vssd1 vccd1 vccd1 _14470__182/HI io_oeb[2] sky130_fd_sc_hd__conb_1
XFILLER_89_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10513__A _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _09998_/A vssd1 vssd1 vccd1 vccd1 _09998_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08949_ _08949_/A _08949_/B vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11960_ _11971_/A vssd1 vssd1 vccd1 vccd1 _11965_/A sky130_fd_sc_hd__buf_2
XFILLER_91_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08918__A _08944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13408__A0 _12561_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ _13926_/Q vssd1 vssd1 vccd1 vccd1 _10912_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11891_ _11893_/B vssd1 vssd1 vccd1 vccd1 _11891_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13630_ _13630_/A vssd1 vssd1 vccd1 vccd1 _14433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10842_ _13982_/Q _10841_/Y _10875_/S vssd1 vssd1 vccd1 vccd1 _10842_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13561_ _13561_/A vssd1 vssd1 vccd1 vccd1 _14413_/D sky130_fd_sc_hd__clkbuf_1
X_10773_ _10773_/A _10773_/B vssd1 vssd1 vccd1 vccd1 _10791_/B sky130_fd_sc_hd__xnor2_1
XFILLER_34_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ _12218_/X _08966_/A _12520_/S vssd1 vssd1 vccd1 vccd1 _12513_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input98_A io_wbs_rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13492_ _13502_/A _13492_/B vssd1 vssd1 vccd1 vccd1 _13493_/A sky130_fd_sc_hd__and2_1
XFILLER_100_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12443_ _08683_/X _12439_/X _12442_/X _14041_/Q vssd1 vssd1 vccd1 vccd1 _12443_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12374_ _12378_/A vssd1 vssd1 vccd1 vccd1 _12374_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ _14239_/CLK _14113_/D vssd1 vssd1 vccd1 vccd1 _14113_/Q sky130_fd_sc_hd__dfxtp_1
X_11325_ _11325_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11325_/Y sky130_fd_sc_hd__nor2_1
X_11256_ _11256_/A vssd1 vssd1 vccd1 vccd1 _11355_/B sky130_fd_sc_hd__clkbuf_2
X_14044_ _14363_/CLK _14044_/D vssd1 vssd1 vccd1 vccd1 _14044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10207_ _10216_/A _10216_/B vssd1 vssd1 vccd1 vccd1 _10211_/A sky130_fd_sc_hd__nor2_1
X_11187_ _11181_/A _11186_/X _11173_/X _10975_/A vssd1 vssd1 vccd1 vccd1 _11187_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_45_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07574__A0 _14095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10138_ _10138_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _10139_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11238__B _11282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13647__A0 input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10069_ _10069_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08828__A _08828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08547__B _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13828_ _14335_/CLK _13828_/D vssd1 vssd1 vccd1 vccd1 _13828_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_16_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13759_ _13820_/CLK _13759_/D _11950_/Y vssd1 vssd1 vccd1 vccd1 _13759_/Q sky130_fd_sc_hd__dfrtp_1
X_07280_ _07280_/A vssd1 vssd1 vccd1 vccd1 _07307_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12085__A _12517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09921_ _09921_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _09956_/A sky130_fd_sc_hd__xor2_2
XANTENNA__12689__A1 _14055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09852_ _10127_/A _10205_/A _09896_/A vssd1 vssd1 vccd1 vccd1 _09959_/B sky130_fd_sc_hd__o21a_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07565__A0 _14099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10333__A _10333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _08803_/A _08803_/B _08814_/B _08803_/D vssd1 vssd1 vccd1 vccd1 _08850_/A
+ sky130_fd_sc_hd__or4_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _10597_/A _09783_/B _09783_/C vssd1 vssd1 vccd1 vccd1 _09783_/X sky130_fd_sc_hd__or3_4
XFILLER_85_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ _14278_/Q _06968_/X _06994_/X _14374_/Q vssd1 vssd1 vccd1 vccd1 _06995_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13644__A _13644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08734_ _08734_/A _08734_/B vssd1 vssd1 vccd1 vccd1 _08735_/C sky130_fd_sc_hd__xnor2_1
XFILLER_27_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11113__A1 _11010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07642__A _14132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _08665_/A _08665_/B _08665_/C vssd1 vssd1 vccd1 vccd1 _08667_/B sky130_fd_sc_hd__nand3_2
XANTENNA__12861__A1 _14133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07616_ _07616_/A vssd1 vssd1 vccd1 vccd1 _14076_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _13866_/Q vssd1 vssd1 vccd1 vccd1 _09811_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07547_ _07547_/A vssd1 vssd1 vccd1 vccd1 _14107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11821__C1 _11820_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ _14194_/Q _14196_/Q _07482_/S vssd1 vssd1 vccd1 vccd1 _07479_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08473__A _13860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09217_ _09543_/A _09217_/B _09296_/D _09217_/D vssd1 vssd1 vccd1 vccd1 _09295_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__08623__D _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _09148_/A _09148_/B _09148_/C vssd1 vssd1 vccd1 vccd1 _09151_/A sky130_fd_sc_hd__or3_1
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09079_ _09079_/A _09079_/B _09079_/C vssd1 vssd1 vccd1 vccd1 _09081_/B sky130_fd_sc_hd__nand3_1
XFILLER_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11110_ _11110_/A vssd1 vssd1 vccd1 vccd1 _11110_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12090_ _12211_/A input65/X vssd1 vssd1 vccd1 vccd1 _12823_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07817__A _14036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11041_ _11041_/A vssd1 vssd1 vccd1 vccd1 _11127_/B sky130_fd_sc_hd__inv_2
XFILLER_39_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07556__A0 _14103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11352__B2 _07784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12992_ _13004_/A vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__buf_2
XFILLER_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A dout1[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ _11947_/A vssd1 vssd1 vccd1 vccd1 _11943_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11874_ hold38/A vssd1 vssd1 vccd1 vccd1 _11874_/X sky130_fd_sc_hd__buf_2
XFILLER_60_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13613_ _13613_/A vssd1 vssd1 vccd1 vccd1 _14428_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12604__A1 _14034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ _10700_/X _10705_/B _10828_/A _10828_/C _10824_/Y vssd1 vssd1 vccd1 vccd1
+ _10825_/X sky130_fd_sc_hd__o221a_1
XFILLER_41_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13544_ _13544_/A vssd1 vssd1 vccd1 vccd1 _14408_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12080__A2 _12000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ _11152_/S _10755_/Y _10716_/B vssd1 vssd1 vccd1 vccd1 _10773_/A sky130_fd_sc_hd__a21oi_1
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13475_ _13084_/X _14389_/Q _13475_/S vssd1 vssd1 vccd1 vccd1 _13476_/B sky130_fd_sc_hd__mux2_1
X_10687_ _13985_/Q _10686_/X _10690_/S vssd1 vssd1 vccd1 vccd1 _10688_/A sky130_fd_sc_hd__mux2_1
X_12426_ _12426_/A vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__clkinv_2
X_12357_ _12360_/A vssd1 vssd1 vccd1 vccd1 _12357_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12633__A input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11308_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11309_/B sky130_fd_sc_hd__xor2_2
XFILLER_113_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12288_ _12291_/A vssd1 vssd1 vccd1 vccd1 _12288_/Y sky130_fd_sc_hd__inv_2
X_14027_ _14028_/CLK _14027_/D vssd1 vssd1 vccd1 vccd1 _14027_/Q sky130_fd_sc_hd__dfxtp_2
X_11239_ _13900_/Q vssd1 vssd1 vccd1 vccd1 _11279_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11343__B2 _07784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09942__A _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07462__A _07462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08450_ _08503_/B _08503_/C _08503_/A vssd1 vssd1 vccd1 vccd1 _08452_/B sky130_fd_sc_hd__a21bo_1
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07401_ _14208_/Q _14210_/Q _07415_/S vssd1 vssd1 vccd1 vccd1 _07402_/B sky130_fd_sc_hd__mux2_1
X_08381_ _08380_/A _08380_/B _08380_/C vssd1 vssd1 vccd1 vccd1 _08381_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07332_ _14105_/Q _07323_/X vssd1 vssd1 vccd1 vccd1 _07332_/X sky130_fd_sc_hd__or2b_1
XFILLER_108_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12071__A2 _12059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07263_ _07263_/A _13836_/Q vssd1 vssd1 vccd1 vccd1 _07459_/A sky130_fd_sc_hd__and2_1
XANTENNA__10328__A _10421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09002_ _08555_/B _08794_/B _09091_/B _09001_/A vssd1 vssd1 vccd1 vccd1 _09003_/C
+ sky130_fd_sc_hd__a22o_1
X_07194_ _14095_/Q _07185_/X _07186_/X vssd1 vssd1 vccd1 vccd1 _07194_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13639__A _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09904_ _08547_/D _09885_/X _09884_/X vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__o21ai_4
XFILLER_99_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input5_A dout1[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ _08291_/C _09553_/D _09241_/D vssd1 vssd1 vccd1 vccd1 _09835_/X sky130_fd_sc_hd__a21o_1
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_115_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10998__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09766_ _09766_/A vssd1 vssd1 vccd1 vccd1 _10367_/A sky130_fd_sc_hd__clkbuf_2
X_06978_ _14456_/Q _14280_/Q vssd1 vssd1 vccd1 vccd1 _06978_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08717_ _08742_/A _08803_/A vssd1 vssd1 vccd1 vccd1 _08743_/A sky130_fd_sc_hd__and2_1
XFILLER_55_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11098__B1 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09697_ _09697_/A _09697_/B vssd1 vssd1 vccd1 vccd1 _09727_/A sky130_fd_sc_hd__or2_1
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07091__B _07098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14370__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _09217_/D vssd1 vssd1 vccd1 vccd1 _09804_/A sky130_fd_sc_hd__buf_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _08579_/A vssd1 vssd1 vccd1 vccd1 _08580_/B sky130_fd_sc_hd__buf_4
XANTENNA__12718__A _12721_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10610_/A _10610_/B vssd1 vssd1 vccd1 vccd1 _10610_/Y sky130_fd_sc_hd__xnor2_1
X_11590_ _11585_/S _11587_/X _11588_/Y _11589_/X vssd1 vssd1 vccd1 vccd1 _13856_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_70_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10541_ _10541_/A _10541_/B vssd1 vssd1 vccd1 vccd1 _10541_/Y sky130_fd_sc_hd__xnor2_4
X_13260_ _14332_/Q _13240_/X _13259_/X _13254_/X vssd1 vssd1 vccd1 vccd1 _14332_/D
+ sky130_fd_sc_hd__o211a_1
X_10472_ _10493_/A _10471_/Y _10472_/S vssd1 vssd1 vccd1 vccd1 _10474_/A sky130_fd_sc_hd__mux2_1
X_12211_ _12211_/A input65/X vssd1 vssd1 vccd1 vccd1 _13358_/A sky130_fd_sc_hd__and2_2
X_13191_ _13193_/A vssd1 vssd1 vccd1 vccd1 _13191_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ _13820_/Q _12133_/X _12141_/X _12131_/X vssd1 vssd1 vccd1 vccd1 _13820_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12073_ _12073_/A vssd1 vssd1 vccd1 vccd1 _13802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11024_ _10970_/C _11035_/A _11252_/A vssd1 vssd1 vccd1 vccd1 _11029_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09762__A _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13284__A _13306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08378__A _08385_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12975_ _12978_/A vssd1 vssd1 vccd1 vccd1 _12975_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08097__B _08097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10420__B _10420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08528__D _09206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11926_ _11926_/A vssd1 vssd1 vccd1 vccd1 _14169_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _11857_/A vssd1 vssd1 vccd1 vccd1 _11857_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10808_ _10863_/B _10869_/A _10863_/A vssd1 vssd1 vccd1 vccd1 _10858_/C sky130_fd_sc_hd__o21ai_1
XFILLER_32_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11788_ _13784_/Q _11823_/A _12773_/A _14109_/Q vssd1 vssd1 vccd1 vccd1 _11788_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13527_ _13614_/A vssd1 vssd1 vccd1 vccd1 _13634_/S sky130_fd_sc_hd__clkbuf_4
X_10739_ _13948_/Q vssd1 vssd1 vccd1 vccd1 _10923_/S sky130_fd_sc_hd__inv_2
XFILLER_51_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13458_ _13461_/A _13458_/B vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__and2_1
XFILLER_12_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12409_ _12409_/A vssd1 vssd1 vccd1 vccd1 _12409_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput105 _14064_/Q vssd1 vssd1 vccd1 vccd1 addr1[4] sky130_fd_sc_hd__buf_2
X_13389_ _13392_/A _13389_/B vssd1 vssd1 vccd1 vccd1 _13390_/A sky130_fd_sc_hd__and2_1
XANTENNA__12363__A _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput116 _11836_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[12] sky130_fd_sc_hd__buf_2
XFILLER_12_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput127 _11853_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[22] sky130_fd_sc_hd__buf_2
XFILLER_114_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput138 _11807_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[3] sky130_fd_sc_hd__buf_2
XFILLER_86_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput149 _14305_/Q vssd1 vssd1 vccd1 vccd1 wfg_drive_pat_dout_o[13] sky130_fd_sc_hd__buf_2
XFILLER_115_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14243__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09400__A1_N _09999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07950_ _14021_/Q vssd1 vssd1 vccd1 vccd1 _09362_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06991__A1 _14311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__A1 _11119_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ _14434_/Q _06900_/Y _06877_/X vssd1 vssd1 vccd1 vccd1 _06901_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09672__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07881_ _07819_/Y _07881_/B vssd1 vssd1 vccd1 vccd1 _07882_/B sky130_fd_sc_hd__and2b_1
XFILLER_110_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11707__A hold6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _09667_/A _09666_/A vssd1 vssd1 vccd1 vccd1 _10576_/A sky130_fd_sc_hd__or2_1
XANTENNA__14393__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09551_ _14020_/Q _14019_/Q _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09594_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_97_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12816__A1 hold7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12816__B2 _14146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08502_ _08590_/B _08502_/B _08502_/C vssd1 vssd1 vccd1 vccd1 _08537_/A sky130_fd_sc_hd__nand3_1
XFILLER_97_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12624__D_N _12441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07299__A2 _14192_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09482_ _09482_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09483_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08433_ _08791_/A vssd1 vssd1 vccd1 vccd1 _09233_/A sky130_fd_sc_hd__buf_2
XFILLER_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08248__A1 _09762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _08366_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13241__B2 _14393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _07452_/A vssd1 vssd1 vccd1 vccd1 _07348_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_65_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_20_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08295_ _08295_/A _08295_/B vssd1 vssd1 vccd1 vccd1 _08295_/Y sky130_fd_sc_hd__nand2_1
X_07246_ _14080_/Q _13880_/Q _07252_/S vssd1 vssd1 vccd1 vccd1 _07246_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09847__A _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07177_ _14284_/Q _07176_/X _07183_/S vssd1 vssd1 vccd1 vccd1 _07178_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10505__B _10505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__B _14266_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09818_ _09818_/A _09818_/B vssd1 vssd1 vccd1 vccd1 _09818_/X sky130_fd_sc_hd__and2_1
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_49_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14348_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_28_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12807__A1 _14158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09749_ _09749_/A _09749_/B _09749_/C vssd1 vssd1 vccd1 vccd1 _09750_/B sky130_fd_sc_hd__or3_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12760_ _12809_/A vssd1 vssd1 vccd1 vccd1 _12760_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08926__A _09055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11920_/A _11882_/A vssd1 vssd1 vccd1 vccd1 _11714_/A sky130_fd_sc_hd__and2_2
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07830__A _14026_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12691_/A vssd1 vssd1 vccd1 vccd1 _14055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14464_/CLK _14430_/D vssd1 vssd1 vccd1 vccd1 _14430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _14043_/Q _13955_/Q vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14361_ _14410_/CLK _14361_/D vssd1 vssd1 vccd1 vccd1 _14361_/Q sky130_fd_sc_hd__dfxtp_1
X_11573_ _11609_/A _11610_/A _11609_/B vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__a21boi_4
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 dout1[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input80_A io_wbs_datwr[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ _14376_/Q _13307_/X _13294_/X _14456_/Q vssd1 vssd1 vccd1 vccd1 _13312_/X
+ sky130_fd_sc_hd__a22o_1
Xinput29 dout1[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
X_10524_ _10524_/A _10524_/B _10524_/C vssd1 vssd1 vccd1 vccd1 _10524_/X sky130_fd_sc_hd__and3_1
X_14292_ _14453_/CLK _14292_/D _13157_/Y vssd1 vssd1 vccd1 vccd1 _14292_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14266__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13243_ _14409_/Q _13199_/X _13241_/X _13242_/X vssd1 vssd1 vccd1 vccd1 _13243_/X
+ sky130_fd_sc_hd__a211o_1
X_10455_ _10455_/A _10455_/B _10455_/C vssd1 vssd1 vccd1 vccd1 _10456_/B sky130_fd_sc_hd__nand3_1
XFILLER_109_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08947__C1 _08683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ _13177_/A vssd1 vssd1 vccd1 vccd1 _13174_/Y sky130_fd_sc_hd__inv_2
X_10386_ _10386_/A _10400_/A vssd1 vssd1 vccd1 vccd1 _10388_/A sky130_fd_sc_hd__xor2_1
XANTENNA_output167_A _14321_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ input72/X vssd1 vssd1 vccd1 vccd1 _12942_/A sky130_fd_sc_hd__buf_6
XFILLER_97_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12911__A _12911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12056_ _13798_/Q _12038_/X _12039_/X hold31/A vssd1 vssd1 vccd1 vccd1 _12057_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_81_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11007_ _11070_/B _11007_/B vssd1 vssd1 vccd1 vccd1 _11104_/B sky130_fd_sc_hd__and2b_1
XFILLER_93_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ _12960_/A vssd1 vssd1 vccd1 vccd1 _12958_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11909_ _11911_/B vssd1 vssd1 vccd1 vccd1 _11909_/Y sky130_fd_sc_hd__inv_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ _12932_/A _12896_/B vssd1 vssd1 vccd1 vccd1 _12889_/X sky130_fd_sc_hd__or2_1
XANTENNA__12358__A _12360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13223__A1 hold33/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07100_ _07097_/X _14297_/Q _07100_/S vssd1 vssd1 vccd1 vccd1 _07101_/A sky130_fd_sc_hd__mux2_1
X_08080_ _08146_/A _08163_/B vssd1 vssd1 vccd1 vccd1 _08081_/C sky130_fd_sc_hd__xor2_1
XANTENNA__08650__A1 _08435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08571__A _08571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07031_ _07031_/A vssd1 vssd1 vccd1 vccd1 _14306_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12093__A _12900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08982_ _08982_/A _08982_/B vssd1 vssd1 vccd1 vccd1 _08986_/A sky130_fd_sc_hd__and2_1
X_07933_ _14022_/Q vssd1 vssd1 vccd1 vccd1 _09145_/B sky130_fd_sc_hd__buf_2
XFILLER_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07864_ _07878_/A vssd1 vssd1 vccd1 vccd1 _07874_/S sky130_fd_sc_hd__buf_2
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10512__A2 _10524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ _09676_/A _09676_/B _09676_/C vssd1 vssd1 vccd1 vccd1 _09603_/X sky130_fd_sc_hd__and3_1
XFILLER_83_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07795_ _10950_/S vssd1 vssd1 vccd1 vccd1 _11164_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09534_ _08982_/A _09510_/B _09510_/C _09459_/A vssd1 vssd1 vccd1 vccd1 _09536_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08746__A _09200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09465_ _09465_/A _09465_/B vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12268__A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08416_ _09188_/A vssd1 vssd1 vccd1 vccd1 _08966_/A sky130_fd_sc_hd__buf_6
XFILLER_58_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09396_ _09360_/Y _09396_/B _09396_/C vssd1 vssd1 vccd1 vccd1 _09396_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__14289__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08347_ _13868_/Q vssd1 vssd1 vccd1 vccd1 _09479_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__09577__A _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08481__A _09865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ _09777_/B _08278_/B vssd1 vssd1 vccd1 vccd1 _08278_/X sky130_fd_sc_hd__or2_1
X_07229_ _14085_/Q _13885_/Q _07235_/S vssd1 vssd1 vccd1 vccd1 _07229_/X sky130_fd_sc_hd__mux2_2
XANTENNA__11528__A1 _08944_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ _10187_/X _10237_/X _10238_/Y _10239_/Y vssd1 vssd1 vccd1 vccd1 _10645_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_105_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10171_ _10171_/A _10171_/B vssd1 vssd1 vccd1 vccd1 _10172_/B sky130_fd_sc_hd__or2_1
XFILLER_78_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07825__A _14030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13930_ _13987_/CLK _13930_/D _12345_/Y vssd1 vssd1 vccd1 vccd1 _13930_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13861_ _13867_/CLK _13861_/D _12258_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12812_ hold1/A _12801_/X _12803_/X _14144_/Q _12809_/X vssd1 vssd1 vccd1 vccd1 _12812_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__13562__A _13634_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13792_ _13809_/CLK _13792_/D vssd1 vssd1 vccd1 vccd1 _13792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08656__A _08656_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _12746_/A vssd1 vssd1 vccd1 vccd1 _12743_/Y sky130_fd_sc_hd__inv_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11082__A _11082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12673_/X _14051_/Q _12685_/S vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__mux2_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _14449_/CLK _14413_/D vssd1 vssd1 vccd1 vccd1 _14413_/Q sky130_fd_sc_hd__dfxtp_1
X_11625_ _11625_/A vssd1 vssd1 vccd1 vccd1 _13848_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12906__A _12906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344_ _14348_/CLK _14344_/D vssd1 vssd1 vccd1 vccd1 _14344_/Q sky130_fd_sc_hd__dfxtp_1
X_11556_ _14043_/Q _13955_/Q _11643_/A vssd1 vssd1 vccd1 vccd1 _11556_/X sky130_fd_sc_hd__a21o_1
X_10507_ _10520_/A _10507_/B vssd1 vssd1 vccd1 vccd1 _10508_/B sky130_fd_sc_hd__and2_1
X_14275_ _14275_/CLK _14275_/D _13136_/Y vssd1 vssd1 vccd1 vccd1 _14275_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_109_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11487_ _11487_/A _11487_/B vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__and2_1
XANTENNA__11519__A1 _11054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13226_ _14406_/Q _13216_/X _13225_/X vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__a21o_1
XFILLER_48_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10438_ _10438_/A _10438_/B _10438_/C vssd1 vssd1 vccd1 vccd1 _10439_/B sky130_fd_sc_hd__nor3_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ _13159_/A vssd1 vssd1 vccd1 vccd1 _13157_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12641__A input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _10369_/A _10369_/B _10369_/C vssd1 vssd1 vccd1 vccd1 _10370_/B sky130_fd_sc_hd__and3_1
XFILLER_3_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ input68/X vssd1 vssd1 vccd1 vccd1 _12932_/A sky130_fd_sc_hd__buf_4
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _12633_/X hold26/A _13096_/S vssd1 vssd1 vccd1 vccd1 _13089_/B sky130_fd_sc_hd__mux2_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12039_ _12060_/A vssd1 vssd1 vccd1 vccd1 _12039_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07580_ _14092_/Q input8/X _07582_/S vssd1 vssd1 vccd1 vccd1 _07581_/A sky130_fd_sc_hd__mux2_1
XFILLER_81_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12088__A _13470_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09250_ _09137_/A _09140_/A _09248_/X _09249_/Y vssd1 vssd1 vccd1 vccd1 _09333_/B
+ sky130_fd_sc_hd__a211o_1
X_08201_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08202_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _09194_/B _09180_/B _09180_/C _09180_/D vssd1 vssd1 vccd1 vccd1 _09181_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08132_ _08132_/A _08208_/B _08289_/A _08132_/D vssd1 vssd1 vccd1 vccd1 _08213_/A
+ sky130_fd_sc_hd__and4_1
X_08063_ _09543_/C vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__clkbuf_4
X_07014_ _07012_/X _07013_/X _14372_/Q vssd1 vssd1 vccd1 vccd1 _07015_/S sky130_fd_sc_hd__o21a_1
XFILLER_108_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06937__A1 _14318_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08965_ _08965_/A _08692_/A vssd1 vssd1 vccd1 vccd1 _08965_/X sky130_fd_sc_hd__or2b_1
XFILLER_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07916_ _07915_/X _13972_/Q _07919_/S vssd1 vssd1 vccd1 vccd1 _07917_/A sky130_fd_sc_hd__mux2_1
X_08896_ _08896_/A _10171_/A _08948_/D vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__nand3_1
XFILLER_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09860__A _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07847_ _07847_/A _07847_/B _07847_/C vssd1 vssd1 vccd1 vccd1 _07848_/B sky130_fd_sc_hd__or3_1
XFILLER_84_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08476__A _13860_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07778_ _10629_/S vssd1 vssd1 vccd1 vccd1 _10585_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_72_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ _09501_/X _09502_/Y _09471_/A _09471_/Y vssd1 vssd1 vccd1 vccd1 _09518_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07114__A1 _07090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09489_/B _09447_/C _09447_/A vssd1 vssd1 vccd1 vccd1 _09448_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08862__A1 _08978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08862__B2 _08978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09379_ _13870_/Q vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11410_ _11355_/A _11134_/A _11415_/A vssd1 vssd1 vccd1 vccd1 _11529_/A sky130_fd_sc_hd__mux2_1
X_12390_ _12391_/A vssd1 vssd1 vccd1 vccd1 _12390_/Y sky130_fd_sc_hd__inv_2
X_11341_ _11341_/A _11341_/B _11345_/A vssd1 vssd1 vccd1 vccd1 _11342_/B sky130_fd_sc_hd__and3_1
XFILLER_119_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14060_ _14075_/CLK _14060_/D _12701_/Y vssd1 vssd1 vccd1 vccd1 _14060_/Q sky130_fd_sc_hd__dfrtp_2
X_11272_ _11347_/A _11347_/B _11348_/A vssd1 vssd1 vccd1 vccd1 _11344_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__12174__A1 _13830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13371__A0 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13011_ _13116_/A vssd1 vssd1 vccd1 vccd1 _13016_/A sky130_fd_sc_hd__buf_2
XANTENNA__08917__A2 _08941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ _10213_/B _10213_/C _10213_/A vssd1 vssd1 vccd1 vccd1 _10223_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11921__A1 _13822_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A io_wbs_adr[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10154_ _10159_/A _10159_/B _10153_/Y vssd1 vssd1 vccd1 vccd1 _10182_/A sky130_fd_sc_hd__o21ai_1
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10085_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__xor2_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__buf_2
XFILLER_75_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13913_ _13915_/CLK _13913_/D _12325_/Y vssd1 vssd1 vccd1 vccd1 _13913_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10488__B2 _09998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13844_ _14028_/CLK _13844_/D _12237_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13775_ _14451_/CLK _13775_/D _11972_/Y vssd1 vssd1 vccd1 vccd1 _13775_/Q sky130_fd_sc_hd__dfrtp_2
X_10987_ _10987_/A _10987_/B vssd1 vssd1 vccd1 vccd1 _11092_/B sky130_fd_sc_hd__xnor2_1
XFILLER_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12726_ _12727_/A vssd1 vssd1 vccd1 vccd1 _12726_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12657_ _12657_/A vssd1 vssd1 vccd1 vccd1 _14047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11540__A _14053_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ _11608_/A vssd1 vssd1 vccd1 vccd1 _13852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08605__B2 _08978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ _12594_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _12589_/A sky130_fd_sc_hd__and2_1
XFILLER_50_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14327_ _14396_/CLK _14327_/D vssd1 vssd1 vccd1 vccd1 _14327_/Q sky130_fd_sc_hd__dfxtp_1
X_11539_ _14054_/Q _13966_/Q vssd1 vssd1 vccd1 vccd1 _11539_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14258_ _14258_/CLK _14258_/D vssd1 vssd1 vccd1 vccd1 _14258_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12165__A1 _13827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13362__A0 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13209_ _13209_/A _13358_/B vssd1 vssd1 vccd1 vccd1 _13341_/A sky130_fd_sc_hd__nand2_8
XFILLER_112_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14189_ _14256_/CLK _14189_/D _12977_/Y vssd1 vssd1 vccd1 vccd1 _14189_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12371__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06919__A1 _06894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12090__B input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08750_/A _08750_/B _09865_/B _13860_/Q vssd1 vssd1 vccd1 vccd1 _08787_/A
+ sky130_fd_sc_hd__and4_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07701_ _07653_/X _07699_/X _07706_/A _14147_/Q _07700_/Y vssd1 vssd1 vccd1 vccd1
+ _07701_/X sky130_fd_sc_hd__o221a_1
XFILLER_94_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08681_ _08681_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08687_/A sky130_fd_sc_hd__or2b_1
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ _07684_/B _07685_/B _07684_/A vssd1 vssd1 vccd1 vccd1 _07679_/A sky130_fd_sc_hd__o21ba_1
XFILLER_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07563_ _14100_/Q input17/X _07571_/S vssd1 vssd1 vccd1 vccd1 _07564_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09302_ _09302_/A _09302_/B _09302_/C vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__and3_1
XFILLER_34_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07494_ _07489_/X _07492_/Y _07493_/X _14190_/Q vssd1 vssd1 vccd1 vccd1 _14190_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_34_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _09233_/A _09233_/B _09233_/C _09233_/D vssd1 vssd1 vccd1 vccd1 _09236_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_21_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09164_ _09164_/A _09079_/A vssd1 vssd1 vccd1 vccd1 _09173_/A sky130_fd_sc_hd__or2b_1
XFILLER_108_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ _08198_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08119_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09095_ _09095_/A _09095_/B vssd1 vssd1 vccd1 vccd1 _09097_/B sky130_fd_sc_hd__xnor2_2
X_08046_ _09482_/A vssd1 vssd1 vccd1 vccd1 _08622_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13377__A _13411_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13105__A0 _12654_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09997_ _10393_/A _09997_/B vssd1 vssd1 vccd1 vccd1 _10032_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09309__C1 _09308_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _08944_/X _08948_/B _10206_/A _08948_/D vssd1 vssd1 vccd1 vccd1 _08948_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_76_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09590__A _09590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08879_ _08879_/A _08879_/B vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08918__B _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ _11140_/B vssd1 vssd1 vccd1 vccd1 _11142_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_57_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07395__B_N _07363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11890_ _13751_/Q _11888_/B _13752_/Q vssd1 vssd1 vccd1 vccd1 _11890_/X sky130_fd_sc_hd__o21a_1
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10841_ _10841_/A _10841_/B vssd1 vssd1 vccd1 vccd1 _10841_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_44_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13560_ _13573_/A _13560_/B vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__and2_1
X_10772_ _10770_/Y _10761_/C _10771_/Y _10757_/X _10765_/B vssd1 vssd1 vccd1 vccd1
+ _10773_/B sky130_fd_sc_hd__o32a_1
XFILLER_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12511_ _12562_/S vssd1 vssd1 vccd1 vccd1 _12520_/S sky130_fd_sc_hd__clkbuf_2
X_13491_ _12650_/X _14394_/Q _13494_/S vssd1 vssd1 vccd1 vccd1 _13492_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12442_ _12476_/A vssd1 vssd1 vccd1 vccd1 _12442_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12373_ _12379_/A vssd1 vssd1 vccd1 vccd1 _12378_/A sky130_fd_sc_hd__buf_2
X_14112_ _14152_/CLK _14112_/D vssd1 vssd1 vccd1 vccd1 _14112_/Q sky130_fd_sc_hd__dfxtp_2
X_11324_ _11324_/A _11324_/B _11324_/C vssd1 vssd1 vccd1 vccd1 _11325_/B sky130_fd_sc_hd__and3_1
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09765__A _10302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14043_ _14363_/CLK _14043_/D vssd1 vssd1 vccd1 vccd1 _14043_/Q sky130_fd_sc_hd__dfxtp_1
X_11255_ _13896_/Q vssd1 vssd1 vccd1 vccd1 _11269_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10704__A _11244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10206_ _10206_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10216_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11186_ _11171_/X _11170_/X _11186_/S vssd1 vssd1 vccd1 vccd1 _11186_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10137_ _10162_/A _10162_/B _10136_/X vssd1 vssd1 vccd1 vccd1 _10141_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10068_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__and2_1
XFILLER_85_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08547__C _08824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ _14335_/CLK _13827_/D vssd1 vssd1 vccd1 vccd1 _13827_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_90_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13758_ _13820_/CLK _13758_/D _11949_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Q sky130_fd_sc_hd__dfrtp_1
X_12709_ _12709_/A vssd1 vssd1 vccd1 vccd1 _12709_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10585__S _10585_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ _13689_/A vssd1 vssd1 vccd1 vccd1 _14450_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12366__A _12366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09378__C _13870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13583__A0 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ _09990_/B _09920_/B vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__xnor2_2
XFILLER_116_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10614__A _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09851_ _09895_/A _09895_/B vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__or2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08802_ _08801_/A _08801_/B _08801_/C vssd1 vssd1 vccd1 vccd1 _08803_/D sky130_fd_sc_hd__a21oi_1
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09781_/A _10515_/B _09781_/C vssd1 vssd1 vccd1 vccd1 _09783_/C sky130_fd_sc_hd__a21oi_1
XFILLER_26_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06994_ _14422_/Q _06993_/Y _06970_/X vssd1 vssd1 vccd1 vccd1 _06994_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08905_/A _10009_/A vssd1 vssd1 vccd1 vccd1 _08734_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11113__A2 _11110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08664_ _08664_/A _08664_/B vssd1 vssd1 vccd1 vccd1 _08665_/C sky130_fd_sc_hd__xnor2_1
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07615_ _14076_/Q input1/X _07615_/S vssd1 vssd1 vccd1 vccd1 _07616_/A sky130_fd_sc_hd__mux2_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _08595_/A _08791_/B _09844_/A _09844_/B vssd1 vssd1 vccd1 vccd1 _08595_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12074__B1 _12060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07546_ _14107_/Q input25/X _07548_/S vssd1 vssd1 vccd1 vccd1 _07547_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10624__A1 _13955_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07477_ _07452_/X _07475_/X _07476_/X _07462_/X _14196_/Q vssd1 vssd1 vccd1 vccd1
+ _14196_/D sky130_fd_sc_hd__a32o_1
XANTENNA__09490__A1 _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08293__A2 _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12276__A _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09216_ _09216_/A _09171_/A vssd1 vssd1 vccd1 vccd1 _09225_/A sky130_fd_sc_hd__or2b_1
XFILLER_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09147_ _09472_/B _09199_/D _09941_/A _09361_/A vssd1 vssd1 vccd1 vccd1 _09148_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07253__A0 _14262_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ _09164_/A _09076_/C _09076_/B vssd1 vssd1 vccd1 vccd1 _09079_/C sky130_fd_sc_hd__o21ai_1
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08029_ _14016_/Q vssd1 vssd1 vccd1 vccd1 _09378_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__09552__A2_N _09233_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11040_ _11050_/A _11050_/B vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07556__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_72_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_40_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07833__A _14025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12991_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11942_ _11971_/A vssd1 vssd1 vccd1 vccd1 _11947_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_45_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _13747_/Q vssd1 vssd1 vccd1 vccd1 _11873_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _13625_/A _13612_/B vssd1 vssd1 vccd1 vccd1 _13613_/A sky130_fd_sc_hd__and2_1
XFILLER_38_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10824_ _13943_/Q _13942_/Q _10708_/B vssd1 vssd1 vccd1 vccd1 _10824_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13543_ _13556_/A _13543_/B vssd1 vssd1 vccd1 vccd1 _13544_/A sky130_fd_sc_hd__and2_1
X_10755_ _10777_/B _11155_/S vssd1 vssd1 vccd1 vccd1 _10755_/Y sky130_fd_sc_hd__nor2_1
X_13474_ _12209_/X _13475_/S _13473_/Y vssd1 vssd1 vccd1 vccd1 _14388_/D sky130_fd_sc_hd__o21a_1
X_10686_ _11467_/A vssd1 vssd1 vccd1 vccd1 _10686_/X sky130_fd_sc_hd__clkbuf_2
X_14477__189 vssd1 vssd1 vccd1 vccd1 _14477__189/HI io_oeb[9] sky130_fd_sc_hd__conb_1
X_12425_ _14007_/Q _12425_/B vssd1 vssd1 vccd1 vccd1 _12425_/X sky130_fd_sc_hd__or2_1
XFILLER_51_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07244__A0 _14265_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _12360_/A vssd1 vssd1 vccd1 vccd1 _12356_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11307_ _11216_/A _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11308_/B sky130_fd_sc_hd__a21bo_1
X_12287_ _12291_/A vssd1 vssd1 vccd1 vccd1 _12287_/Y sky130_fd_sc_hd__inv_2
X_14026_ _14028_/CLK _14026_/D vssd1 vssd1 vccd1 vccd1 _14026_/Q sky130_fd_sc_hd__dfxtp_2
X_11238_ _11282_/A _11282_/B vssd1 vssd1 vccd1 vccd1 _11333_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11169_ _13925_/Q _10912_/A _11169_/S vssd1 vssd1 vccd1 vccd1 _11169_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14022__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13480__A _13485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07400_ _07464_/A vssd1 vssd1 vccd1 vccd1 _07528_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08380_ _08380_/A _08380_/B _08380_/C vssd1 vssd1 vccd1 vccd1 _08380_/X sky130_fd_sc_hd__and3_1
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07331_ _14223_/Q _07311_/X _07316_/X _07330_/X vssd1 vssd1 vccd1 vccd1 _14223_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12096__A input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07262_ _13837_/Q vssd1 vssd1 vccd1 vccd1 _07263_/A sky130_fd_sc_hd__inv_2
X_09001_ _09001_/A _09001_/B _09152_/B _09091_/B vssd1 vssd1 vccd1 vccd1 _09072_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_117_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07193_ _07193_/A vssd1 vssd1 vccd1 vccd1 _14280_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09224__A1 _09223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__A0 _14083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09903_ _09903_/A vssd1 vssd1 vccd1 vccd1 _09903_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09834_ _09834_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _10004_/A sky130_fd_sc_hd__xnor2_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10542__B1 _10541_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14453_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_115_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09765_ _10302_/A vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06977_ _06977_/A vssd1 vssd1 vccd1 vccd1 _14313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08716_ _08716_/A _08716_/B _08925_/C _10057_/A vssd1 vssd1 vccd1 vccd1 _08803_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_6_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11098__B2 _11082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09696_ _09696_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09697_/B sky130_fd_sc_hd__and2_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _08587_/A _08585_/X _08586_/A vssd1 vssd1 vccd1 vccd1 _08667_/A sky130_fd_sc_hd__a21o_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11903__A _11906_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08578_ _09491_/A _09882_/A vssd1 vssd1 vccd1 vccd1 _08578_/Y sky130_fd_sc_hd__nand2_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _14184_/Q _07526_/X _07528_/X _14192_/D vssd1 vssd1 vccd1 vccd1 _14176_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _10540_/A _10540_/B vssd1 vssd1 vccd1 vccd1 _10541_/B sky130_fd_sc_hd__or2_2
XFILLER_109_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ _10471_/A vssd1 vssd1 vccd1 vccd1 _10471_/Y sky130_fd_sc_hd__inv_2
X_12210_ _13359_/A vssd1 vssd1 vccd1 vccd1 _12210_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07226__A0 _14086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__A _14028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ _13193_/A vssd1 vssd1 vccd1 vccd1 _13190_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_78_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14179_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_12141_ input79/X _12143_/B vssd1 vssd1 vccd1 vccd1 _12141_/X sky130_fd_sc_hd__or2_1
XFILLER_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12072_ _12081_/A _12072_/B vssd1 vssd1 vccd1 vccd1 _12073_/A sky130_fd_sc_hd__and2_1
XFILLER_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11023_ _13916_/Q vssd1 vssd1 vccd1 vccd1 _11056_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_103_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09762__B _09762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08659__A _13870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11085__A _11092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ _12978_/A vssd1 vssd1 vccd1 vccd1 _12974_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11925_ _14193_/Q _11924_/X _11925_/S vssd1 vssd1 vccd1 vccd1 _11926_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12909__A _12909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07701__B2 _14147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11856_ _14348_/Q _11864_/B vssd1 vssd1 vccd1 vccd1 _11857_/A sky130_fd_sc_hd__and2_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10807_ _10858_/B _10807_/B vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__and2_1
X_11787_ _13990_/Q _11809_/A _11770_/X _14233_/Q vssd1 vssd1 vccd1 vccd1 _11790_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13526_ _13526_/A _13637_/B vssd1 vssd1 vccd1 vccd1 _13614_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10738_ _13937_/Q _10809_/B vssd1 vssd1 vccd1 vccd1 _10853_/B sky130_fd_sc_hd__and2_1
XANTENNA__13538__A0 input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10148__B _10149_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13457_ input86/X _14384_/Q _13460_/S vssd1 vssd1 vccd1 vccd1 _13458_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10669_ _10826_/A vssd1 vssd1 vccd1 vccd1 _10669_/X sky130_fd_sc_hd__buf_4
XFILLER_51_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12408_ _12409_/A vssd1 vssd1 vccd1 vccd1 _12408_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13388_ _12660_/X _14364_/Q _13391_/S vssd1 vssd1 vccd1 vccd1 _13389_/B sky130_fd_sc_hd__mux2_1
Xoutput106 _14065_/Q vssd1 vssd1 vccd1 vccd1 addr1[5] sky130_fd_sc_hd__buf_2
XFILLER_86_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput117 _11838_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[13] sky130_fd_sc_hd__buf_2
Xoutput128 _11854_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[23] sky130_fd_sc_hd__buf_2
X_12339_ _12341_/A vssd1 vssd1 vccd1 vccd1 _12339_/Y sky130_fd_sc_hd__inv_2
Xoutput139 _11813_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[4] sky130_fd_sc_hd__buf_2
XFILLER_114_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06900_ _14466_/Q _14290_/Q vssd1 vssd1 vccd1 vccd1 _06900_/Y sky130_fd_sc_hd__nand2_1
X_14009_ _14417_/CLK _14009_/D vssd1 vssd1 vccd1 vccd1 _14009_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_68_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07880_ _07880_/A vssd1 vssd1 vccd1 vccd1 _13981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09550_ _09479_/B _09123_/C _09818_/B _09153_/A vssd1 vssd1 vccd1 vccd1 _09550_/Y
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__12816__A2 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08501_ _08590_/A _08471_/B _08471_/C vssd1 vssd1 vccd1 vccd1 _08502_/C sky130_fd_sc_hd__a21o_1
XFILLER_36_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10827__B2 _10826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ _09481_/A _09481_/B vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__or2_1
XFILLER_58_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11723__A _11882_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08432_ _14014_/Q vssd1 vssd1 vccd1 vccd1 _08791_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08363_ _08366_/B _08363_/B _08363_/C vssd1 vssd1 vccd1 vccd1 _09601_/A sky130_fd_sc_hd__nand3_2
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08248__A2 _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13241__A2 _13201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07314_ _07374_/A vssd1 vssd1 vccd1 vccd1 _07452_/A sky130_fd_sc_hd__buf_2
X_08294_ _08295_/A _08295_/B vssd1 vssd1 vccd1 vccd1 _08323_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13529__A0 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07245_ _07245_/A vssd1 vssd1 vccd1 vccd1 _14265_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09847__B _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07176_ _14100_/Q _07167_/X _07168_/X vssd1 vssd1 vccd1 vccd1 _07176_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10763__A0 _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13701__A0 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09857_/B sky130_fd_sc_hd__xor2_4
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08198__B _08198_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09748_ _09725_/X _09741_/X _09745_/X _09741_/B _10530_/A vssd1 vssd1 vccd1 vccd1
+ _10524_/B sky130_fd_sc_hd__a221o_4
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09676_/B _09676_/Y _09677_/Y _09678_/X vssd1 vssd1 vccd1 vccd1 _09687_/A
+ sky130_fd_sc_hd__a211oi_4
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08926__B _08944_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ hold5/A _11710_/B vssd1 vssd1 vccd1 vccd1 _11715_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11491__A1 _11007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12696_/A _12690_/B vssd1 vssd1 vccd1 vccd1 _12691_/A sky130_fd_sc_hd__and2_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11641_/A vssd1 vssd1 vccd1 vccd1 _13844_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14360_ _14365_/CLK _14360_/D vssd1 vssd1 vccd1 vccd1 _14360_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11572_ _14051_/Q _13963_/Q vssd1 vssd1 vccd1 vccd1 _11609_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _13332_/A vssd1 vssd1 vccd1 vccd1 _13311_/X sky130_fd_sc_hd__clkbuf_2
Xinput19 dout1[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
X_10523_ _09751_/Y _10523_/B vssd1 vssd1 vccd1 vccd1 _10524_/C sky130_fd_sc_hd__and2b_1
X_14291_ _14322_/CLK _14291_/D _13156_/Y vssd1 vssd1 vccd1 vccd1 _14291_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12464__A _12485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13242_ _14361_/Q _13236_/X _13210_/X vssd1 vssd1 vccd1 vccd1 _13242_/X sky130_fd_sc_hd__a21o_1
XANTENNA_input73_A io_wbs_datwr[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _10455_/B _10455_/C _10455_/A vssd1 vssd1 vccd1 vccd1 _10456_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08947__B1 _08937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ _13177_/A vssd1 vssd1 vccd1 vccd1 _13173_/Y sky130_fd_sc_hd__inv_2
X_10385_ _10353_/A _10353_/B _10384_/X vssd1 vssd1 vccd1 vccd1 _10400_/A sky130_fd_sc_hd__o21a_1
XFILLER_112_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12124_ _13813_/Q _12117_/X _12123_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _13813_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11808__A _11855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _12055_/A vssd1 vssd1 vccd1 vccd1 _13797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11006_ _13921_/Q vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_78_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12957_ _12960_/A vssd1 vssd1 vccd1 vccd1 _12957_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08836__B _08836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11908_ _13757_/Q _11906_/B _13758_/Q vssd1 vssd1 vccd1 vccd1 _11908_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _14143_/Q _12885_/X _12887_/X _12879_/X vssd1 vssd1 vccd1 vccd1 _14143_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08555__C _09870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11839_ _14338_/Q _11855_/A _11830_/X _14122_/Q vssd1 vssd1 vccd1 vccd1 _11839_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13223__A2 _13215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _13518_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13510_/A sky130_fd_sc_hd__and2_1
XANTENNA__08650__A2 _08836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08571__B _08944_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07030_ _07026_/X _14306_/Q _07030_/S vssd1 vssd1 vccd1 vccd1 _07031_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10745__B1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14360__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ _08981_/A _08981_/B vssd1 vssd1 vccd1 vccd1 _08991_/A sky130_fd_sc_hd__xnor2_2
XFILLER_69_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07932_ _09145_/A vssd1 vssd1 vccd1 vccd1 _09084_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09363__B1 _09200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07863_ _13985_/Q _07863_/B vssd1 vssd1 vccd1 vccd1 _13985_/D sky130_fd_sc_hd__xnor2_1
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ _09601_/A _09601_/B _09601_/C vssd1 vssd1 vccd1 vccd1 _09676_/C sky130_fd_sc_hd__a21o_1
XFILLER_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07794_ _13949_/Q vssd1 vssd1 vccd1 vccd1 _10950_/S sky130_fd_sc_hd__buf_2
XFILLER_3_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09533_ _09499_/A _09498_/B _09496_/X vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07931__A _14023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12670__A0 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _09464_/A _09464_/B vssd1 vssd1 vccd1 vccd1 _09465_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08415_ _09044_/A vssd1 vssd1 vccd1 vccd1 _09188_/A sky130_fd_sc_hd__buf_4
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09395_ _09393_/A _09393_/Y _09390_/X _09392_/Y vssd1 vssd1 vccd1 vccd1 _09396_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_12_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08346_ _09424_/B _09217_/D _09843_/A _09424_/A vssd1 vssd1 vccd1 vccd1 _09555_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11599__S _11611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08277_ _08277_/A _08277_/B vssd1 vssd1 vccd1 vccd1 _08280_/A sky130_fd_sc_hd__nand2_1
X_07228_ _07228_/A vssd1 vssd1 vccd1 vccd1 _14270_/D sky130_fd_sc_hd__clkbuf_1
X_07159_ _14289_/Q _07158_/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07160_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10170_ _08836_/B _09847_/X _09848_/X vssd1 vssd1 vccd1 vccd1 _10279_/B sky130_fd_sc_hd__o21a_4
XANTENNA_clkbuf_leaf_11_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_105_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12489__B1 _12488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _13897_/CLK _13860_/D _12257_/Y vssd1 vssd1 vccd1 vccd1 _13860_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08937__A _08946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07841__A _14029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ _14118_/Q _12800_/X _12810_/X _12805_/X vssd1 vssd1 vccd1 vccd1 _14118_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13791_ _14396_/CLK _13791_/D vssd1 vssd1 vccd1 vccd1 _13791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__A0 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12746_/A vssd1 vssd1 vccd1 vccd1 _12742_/Y sky130_fd_sc_hd__inv_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ input68/X vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__buf_4
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13205__A2 _13201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14412_ _14449_/CLK _14412_/D vssd1 vssd1 vccd1 vccd1 _14412_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ hold28/A _11623_/Y _11632_/S vssd1 vssd1 vccd1 vccd1 _11625_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14343_ _14348_/CLK _14343_/D vssd1 vssd1 vccd1 vccd1 _14343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11555_ _11646_/A _11647_/A _11554_/Y vssd1 vssd1 vccd1 vccd1 _11643_/A sky130_fd_sc_hd__o21ai_1
XFILLER_6_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10506_ _10506_/A _10506_/B vssd1 vssd1 vccd1 vccd1 _10506_/Y sky130_fd_sc_hd__xnor2_1
X_14274_ _14275_/CLK _14274_/D _13134_/Y vssd1 vssd1 vccd1 vccd1 _14274_/Q sky130_fd_sc_hd__dfrtp_4
X_11486_ _11510_/A vssd1 vssd1 vccd1 vccd1 _11486_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13225_ _14438_/Q _13336_/A _13218_/X _14390_/Q vssd1 vssd1 vccd1 vccd1 _13225_/X
+ sky130_fd_sc_hd__a22o_1
X_10437_ _10438_/B _10438_/C _10438_/A vssd1 vssd1 vccd1 vccd1 _10439_/A sky130_fd_sc_hd__o21a_1
XANTENNA__12922__A _12922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ _13159_/A vssd1 vssd1 vccd1 vccd1 _13156_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _10369_/B _10369_/C _10369_/A vssd1 vssd1 vccd1 vccd1 _10377_/B sky130_fd_sc_hd__a21oi_1
XFILLER_98_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12107_ hold40/A _12095_/X _12106_/X _11931_/X vssd1 vssd1 vccd1 vccd1 _13809_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11538__A _14055_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13087_ _13087_/A vssd1 vssd1 vccd1 vccd1 _14247_/D sky130_fd_sc_hd__clkbuf_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _10407_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10374_/B sky130_fd_sc_hd__nand2_1
X_12038_ _12059_/A vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07751__A _14153_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12369__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13989_ _14441_/CLK _13989_/D vssd1 vssd1 vccd1 vccd1 _13989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08200_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08243_/C sky130_fd_sc_hd__or2_1
XFILLER_61_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09180_ _09194_/B _09180_/B _09180_/C _09180_/D vssd1 vssd1 vccd1 vccd1 _09180_/Y
+ sky130_fd_sc_hd__nand4_4
XANTENNA_clkbuf_0_io_wbs_clk_A io_wbs_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _08131_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _08215_/A sky130_fd_sc_hd__xnor2_2
XFILLER_105_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08062_ _13873_/Q vssd1 vssd1 vccd1 vccd1 _09543_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_31_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07013_ _14420_/Q _07020_/B _14452_/Q vssd1 vssd1 vccd1 vccd1 _07013_/X sky130_fd_sc_hd__and3b_1
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12832__A _13072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07926__A _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08964_ _08964_/A _08964_/B vssd1 vssd1 vccd1 vccd1 _08964_/Y sky130_fd_sc_hd__nand2_1
XFILLER_64_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07915_ _07915_/A _07915_/B vssd1 vssd1 vccd1 vccd1 _07915_/X sky130_fd_sc_hd__xor2_1
XFILLER_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08895_ _08895_/A _08895_/B vssd1 vssd1 vccd1 vccd1 _08948_/D sky130_fd_sc_hd__xnor2_1
XFILLER_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13663__A _13680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _07824_/Y _07893_/A _07892_/B vssd1 vssd1 vccd1 vccd1 _07847_/C sky130_fd_sc_hd__o21a_1
XFILLER_68_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_77_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__14256__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _10655_/A _07806_/B _07786_/A vssd1 vssd1 vccd1 vccd1 _10629_/S sky130_fd_sc_hd__and3b_4
XANTENNA__12279__A _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ _09516_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _09518_/B sky130_fd_sc_hd__xor2_2
XANTENNA__11446__A1 _10912_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08311__A1 _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__B2 _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09447_ _09447_/A _09489_/B _09447_/C vssd1 vssd1 vccd1 vccd1 _09449_/A sky130_fd_sc_hd__and3_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08862__A2 _08494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ _09378_/A _09378_/B _13870_/Q _13869_/Q vssd1 vssd1 vccd1 vccd1 _09441_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__08492__A _13862_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08329_ _08389_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08391_/C sky130_fd_sc_hd__xnor2_1
XFILLER_21_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ _11279_/A _11319_/X _11339_/Y _11322_/X vssd1 vssd1 vccd1 vccd1 _13900_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11271_ _11271_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11348_/A sky130_fd_sc_hd__xor2_1
X_13010_ _13010_/A vssd1 vssd1 vccd1 vccd1 _13116_/A sky130_fd_sc_hd__clkbuf_2
X_10222_ _10204_/B _10204_/C _10204_/A vssd1 vssd1 vccd1 vccd1 _10222_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13371__A1 _14359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__A _14026_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10185__A1 _10279_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07050__A1 _14271_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _10285_/B _10153_/B vssd1 vssd1 vccd1 vccd1 _10153_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10084_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10138_/A sky130_fd_sc_hd__nor2_1
XANTENNA_input36_A io_wbs_adr[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13912_ _13915_/CLK _13912_/D _12322_/Y vssd1 vssd1 vccd1 vccd1 _13912_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_43_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10488__A2 _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13843_ _14028_/CLK _13843_/D _12236_/Y vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dfrtp_1
XFILLER_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12634__A0 _12633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13774_ _14451_/CLK _13774_/D vssd1 vssd1 vccd1 vccd1 _13774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10986_ _10700_/X _10990_/A _10990_/B vssd1 vssd1 vccd1 vccd1 _10987_/B sky130_fd_sc_hd__o21a_1
XFILLER_15_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12725_ _12727_/A vssd1 vssd1 vccd1 vccd1 _12725_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12917__A _12917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12656_ _12656_/A _12656_/B vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__and2_1
XFILLER_54_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ _13852_/Q _11606_/Y _11611_/S vssd1 vssd1 vccd1 vccd1 _11608_/A sky130_fd_sc_hd__mux2_1
X_12587_ _12917_/A _14029_/Q _12600_/S vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14326_ _14396_/CLK _14326_/D vssd1 vssd1 vccd1 vccd1 _14326_/Q sky130_fd_sc_hd__dfxtp_1
X_11538_ _14055_/Q _13967_/Q vssd1 vssd1 vccd1 vccd1 _11591_/A sky130_fd_sc_hd__or2_1
XFILLER_8_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11967__S _13184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14257_ _14258_/CLK _14257_/D vssd1 vssd1 vccd1 vccd1 _14257_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10871__S _10871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11469_ _11082_/A _11460_/X _11461_/X vssd1 vssd1 vccd1 vccd1 _11469_/X sky130_fd_sc_hd__o21a_1
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13362__A1 _14356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ _13236_/A vssd1 vssd1 vccd1 vccd1 _13208_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ _14284_/CLK _14188_/D _12976_/Y vssd1 vssd1 vccd1 vccd1 _14188_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07041__A1 _14272_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13139_ _13140_/A vssd1 vssd1 vccd1 vccd1 _13139_/Y sky130_fd_sc_hd__inv_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_0_0_io_wbs_clk_A clkbuf_2_1_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_97_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09961__A _10091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07700_ _07700_/A _07700_/B vssd1 vssd1 vccd1 vccd1 _07700_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08680_ _09044_/A _10486_/S vssd1 vssd1 vccd1 vccd1 _08689_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07631_ _14126_/Q _14061_/Q vssd1 vssd1 vccd1 vccd1 _07684_/A sky130_fd_sc_hd__and2_1
XFILLER_54_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11428__A1 _11014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ _07595_/A vssd1 vssd1 vccd1 vccd1 _07571_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09301_ _09377_/A _09299_/C _09299_/B vssd1 vssd1 vccd1 vccd1 _09302_/C sky130_fd_sc_hd__o21ai_1
XFILLER_80_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07493_ _07276_/B _07534_/B _07399_/A vssd1 vssd1 vccd1 vccd1 _07493_/X sky130_fd_sc_hd__a21bo_1
XFILLER_62_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12827__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09232_ _09229_/X _09230_/Y _09198_/A _09198_/Y vssd1 vssd1 vccd1 vccd1 _09276_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09163_ _09161_/A _09161_/B _09161_/C vssd1 vssd1 vccd1 vccd1 _09198_/C sky130_fd_sc_hd__a21o_1
XFILLER_21_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08114_ _08295_/A vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13952__RESET_B _12372_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09094_ _09094_/A _09094_/B vssd1 vssd1 vccd1 vccd1 _09095_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08045_ _14018_/Q vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__buf_2
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10082__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ _09996_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _10610_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09309__B1 _09307_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08947_ _08944_/D _08946_/Y _08937_/C _08683_/X _08944_/C vssd1 vssd1 vccd1 vccd1
+ _08948_/B sky130_fd_sc_hd__o2111a_1
XFILLER_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08878_ _08844_/B _08844_/C _08844_/A vssd1 vssd1 vccd1 vccd1 _08879_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08487__A _09443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07391__A _14227_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07829_ _14027_/Q _13973_/Q vssd1 vssd1 vccd1 vccd1 _07909_/A sky130_fd_sc_hd__or2_1
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10840_ _10840_/A _10840_/B vssd1 vssd1 vccd1 vccd1 _10841_/B sky130_fd_sc_hd__or2_1
XFILLER_44_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07099__A1 _07090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _13950_/Q _13949_/Q vssd1 vssd1 vccd1 vccd1 _10771_/Y sky130_fd_sc_hd__nor2_2
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12510_ _13079_/A _12567_/B vssd1 vssd1 vccd1 vccd1 _12562_/S sky130_fd_sc_hd__or2_4
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13490_ _13490_/A vssd1 vssd1 vccd1 vccd1 _14393_/D sky130_fd_sc_hd__clkbuf_1
X_12441_ _12441_/A vssd1 vssd1 vccd1 vccd1 _12476_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12372_ _12372_/A vssd1 vssd1 vccd1 vccd1 _12372_/Y sky130_fd_sc_hd__clkinv_2
X_11323_ _11297_/A _11319_/X _11321_/Y _11322_/X vssd1 vssd1 vccd1 vccd1 _13906_/D
+ sky130_fd_sc_hd__o22a_1
X_14111_ _14250_/CLK _14111_/D vssd1 vssd1 vccd1 vccd1 _14111_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11254_ _11271_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11344_/B sky130_fd_sc_hd__nand2_1
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14042_ _14054_/CLK _14042_/D vssd1 vssd1 vccd1 vccd1 _14042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10205_ _10205_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10213_/A sky130_fd_sc_hd__xor2_1
X_11185_ _10761_/B _11184_/X _11140_/X vssd1 vssd1 vccd1 vccd1 _11185_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10136_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10136_/X sky130_fd_sc_hd__and2_1
XANTENNA_output142_A _11822_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10067_ _10067_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _10085_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08397__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12607__A0 _12932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__D _08547_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13826_ _13826_/CLK _13826_/D vssd1 vssd1 vccd1 vccd1 _13826_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_91_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13757_ _13820_/CLK _13757_/D _11947_/Y vssd1 vssd1 vccd1 vccd1 _13757_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13280__B1 _13245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10866__S _10871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ _10648_/A _10965_/X _10975_/B _10744_/X _10968_/X vssd1 vssd1 vccd1 vccd1
+ _11035_/A sky130_fd_sc_hd__a221oi_4
XFILLER_31_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12708_ _12709_/A vssd1 vssd1 vccd1 vccd1 _12708_/Y sky130_fd_sc_hd__inv_2
X_13688_ _13695_/A _13688_/B vssd1 vssd1 vccd1 vccd1 _13689_/A sky130_fd_sc_hd__and2_1
XFILLER_31_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ _12656_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__and2_1
XFILLER_15_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09378__D _13869_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08860__A _08944_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14309_ _14417_/CLK _14309_/D _13177_/Y vssd1 vssd1 vccd1 vccd1 _14309_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09850_ _10127_/A _10126_/A vssd1 vssd1 vccd1 vccd1 _09895_/B sky130_fd_sc_hd__xnor2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _08801_/A _08801_/B _08801_/C vssd1 vssd1 vccd1 vccd1 _08814_/B sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_29_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13905_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13099__A0 _12645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _14454_/Q _14278_/Q vssd1 vssd1 vccd1 vccd1 _06993_/Y sky130_fd_sc_hd__nand2_1
X_09781_ _09781_/A _10515_/B _09781_/C vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__and3_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _08731_/A _08731_/C _08764_/A vssd1 vssd1 vccd1 vccd1 _08735_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12846__A0 _12645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08663_ _08663_/A _08663_/B vssd1 vssd1 vccd1 vccd1 _08664_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07614_ _07614_/A vssd1 vssd1 vccd1 vccd1 _14077_/D sky130_fd_sc_hd__clkbuf_1
X_08594_ _09207_/C vssd1 vssd1 vccd1 vccd1 _09844_/B sky130_fd_sc_hd__buf_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07545_ _14256_/Q vssd1 vssd1 vccd1 vccd1 _07548_/S sky130_fd_sc_hd__buf_4
XFILLER_35_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11461__A _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07476_ _14079_/Q _07459_/X _07460_/X _13879_/Q _07471_/X vssd1 vssd1 vccd1 vccd1
+ _07476_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09490__A2 _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09215_ _09215_/A _09215_/B _09215_/C vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__nand3_2
XFILLER_72_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09866__A _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _09362_/A _09870_/A vssd1 vssd1 vccd1 vccd1 _09148_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14444__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09077_ _09015_/A _09014_/B _09014_/A vssd1 vssd1 vccd1 vccd1 _09079_/B sky130_fd_sc_hd__o21bai_2
Xclkbuf_leaf_68_io_wbs_clk clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14258_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07386__A _14095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08028_ _14017_/Q vssd1 vssd1 vccd1 vccd1 _09443_/A sky130_fd_sc_hd__buf_2
XANTENNA__11337__B1 _10851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10524__B _10524_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07005__A1 _14309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09979_ _10285_/B _10159_/A vssd1 vssd1 vccd1 vccd1 _09980_/B sky130_fd_sc_hd__xnor2_2
XFILLER_44_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12837__A0 _12633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12990_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12990_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11941_ _12223_/A vssd1 vssd1 vccd1 vccd1 _11971_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08010__A _13873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11872_/A vssd1 vssd1 vccd1 vccd1 _11872_/X sky130_fd_sc_hd__buf_2
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08945__A _10171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ input82/X _14428_/Q _13611_/S vssd1 vssd1 vccd1 vccd1 _13612_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10823_ _10832_/A _10832_/B vssd1 vssd1 vccd1 vccd1 _10828_/C sky130_fd_sc_hd__or2_1
XFILLER_38_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ input92/X _14408_/Q _13542_/S vssd1 vssd1 vccd1 vccd1 _13543_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11812__B2 _14236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10754_ _13934_/Q _10800_/B vssd1 vssd1 vccd1 vccd1 _10868_/B sky130_fd_sc_hd__and2_1
XFILLER_13_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13473_ _06881_/Y _13475_/S _11935_/A vssd1 vssd1 vccd1 vccd1 _13473_/Y sky130_fd_sc_hd__a21oi_1
X_10685_ _13946_/Q vssd1 vssd1 vccd1 vccd1 _11467_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12424_ _12429_/A _11988_/A _12440_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _12425_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08680__A _09044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12355_ _12379_/A vssd1 vssd1 vccd1 vccd1 _12360_/A sky130_fd_sc_hd__buf_4
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13811__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _11311_/B _11312_/A _11312_/B _11305_/Y vssd1 vssd1 vccd1 vccd1 _11309_/A
+ sky130_fd_sc_hd__a31o_1
X_12286_ _12286_/A vssd1 vssd1 vccd1 vccd1 _12291_/A sky130_fd_sc_hd__buf_2
XFILLER_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11237_ _11237_/A _11237_/B vssd1 vssd1 vccd1 vccd1 _11282_/B sky130_fd_sc_hd__xnor2_4
XFILLER_45_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14025_ _14275_/CLK _14025_/D vssd1 vssd1 vccd1 vccd1 _14025_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_106_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12930__A _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ _10648_/A _11164_/X _11167_/X vssd1 vssd1 vccd1 vccd1 _11262_/C sky130_fd_sc_hd__a21oi_2
XFILLER_45_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13961__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10119_ _10383_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _10120_/C sky130_fd_sc_hd__xnor2_1
X_11099_ _11080_/X _11099_/B _11099_/C vssd1 vssd1 vccd1 vccd1 _11099_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_64_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07180__A0 _14283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13809_ _13809_/CLK _13809_/D vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07330_ _07321_/X _07327_/X _07328_/X _07329_/X vssd1 vssd1 vccd1 vccd1 _07330_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07261_ _14165_/Q vssd1 vssd1 vccd1 vccd1 _07274_/A sky130_fd_sc_hd__clkbuf_2
X_09000_ _09000_/A _09000_/B vssd1 vssd1 vccd1 vccd1 _09000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07192_ _14280_/Q _07191_/X _07201_/S vssd1 vssd1 vccd1 vccd1 _07193_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09224__A2 _09223_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _10191_/A _09902_/B vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__xnor2_2
XFILLER_28_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07934__A _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _10436_/B vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__inv_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06887__A1_N _14392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__B2 _10528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_16_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_6_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09188_/B _09088_/A _09762_/Y _10528_/A vssd1 vssd1 vccd1 vccd1 _09764_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_74_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06976_ _06972_/X _14313_/Q _06976_/S vssd1 vssd1 vccd1 vccd1 _06977_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08715_ _09084_/D vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09695_ _09696_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09697_/A sky130_fd_sc_hd__nor2_2
XFILLER_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _08645_/A _08645_/C _08645_/B vssd1 vssd1 vccd1 vccd1 _08675_/C sky130_fd_sc_hd__a21oi_2
XANTENNA__07171__A0 _14286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ _08716_/B _08899_/A _08558_/B _08555_/X vssd1 vssd1 vccd1 vccd1 _08587_/A
+ sky130_fd_sc_hd__a31o_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07528_ _07528_/A _07528_/B _07520_/B vssd1 vssd1 vccd1 vccd1 _07528_/X sky130_fd_sc_hd__or3b_1
XFILLER_70_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07459_ _07459_/A vssd1 vssd1 vccd1 vccd1 _07459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10470_ _10485_/B _10470_/B vssd1 vssd1 vccd1 vccd1 _10473_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09129_ _09060_/B _09060_/C _09060_/A vssd1 vssd1 vccd1 vccd1 _09130_/C sky130_fd_sc_hd__a21bo_1
XFILLER_68_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12140_ _13819_/Q _12133_/X _12139_/X _12131_/X vssd1 vssd1 vccd1 vccd1 _13819_/D
+ sky130_fd_sc_hd__o211a_1
X_12071_ _13802_/Q _12059_/X _12060_/X _13818_/Q vssd1 vssd1 vccd1 vccd1 _12072_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _11058_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11117_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12973_ _12973_/A vssd1 vssd1 vccd1 vccd1 _12978_/A sky130_fd_sc_hd__buf_2
XFILLER_92_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11924_ _14200_/Q _14208_/Q _14216_/Q _14224_/Q _14230_/Q _14231_/Q vssd1 vssd1 vccd1
+ vccd1 _11924_/X sky130_fd_sc_hd__mux4_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07162__A0 _14288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11855_ _11855_/A vssd1 vssd1 vccd1 vccd1 _11864_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06907__B _14262_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10806_ _13936_/Q _10806_/B vssd1 vssd1 vccd1 vccd1 _10807_/B sky130_fd_sc_hd__or2_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11786_ _11786_/A vssd1 vssd1 vccd1 vccd1 _11786_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13525_ _13525_/A vssd1 vssd1 vccd1 vccd1 _13637_/B sky130_fd_sc_hd__inv_2
X_10737_ _10746_/A _11228_/A _10737_/S vssd1 vssd1 vccd1 vccd1 _10809_/B sky130_fd_sc_hd__mux2_1
XFILLER_9_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13456_ _13456_/A vssd1 vssd1 vccd1 vccd1 _14383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ _11108_/A _07804_/B _10663_/Y _11319_/A _11152_/S vssd1 vssd1 vccd1 vccd1
+ _13949_/D sky130_fd_sc_hd__o32ai_1
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12407_ _12409_/A vssd1 vssd1 vccd1 vccd1 _12407_/Y sky130_fd_sc_hd__inv_2
X_13387_ _13387_/A vssd1 vssd1 vccd1 vccd1 _14363_/D sky130_fd_sc_hd__clkbuf_1
X_10599_ _10614_/A _10588_/B _10598_/X _10562_/B vssd1 vssd1 vccd1 vccd1 _10599_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_103_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput107 _14066_/Q vssd1 vssd1 vccd1 vccd1 addr1[6] sky130_fd_sc_hd__buf_2
XFILLER_115_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput118 _11840_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[14] sky130_fd_sc_hd__buf_2
XFILLER_56_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _12341_/A vssd1 vssd1 vccd1 vccd1 _12338_/Y sky130_fd_sc_hd__inv_2
Xoutput129 _11857_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[24] sky130_fd_sc_hd__buf_2
XFILLER_47_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12660__A input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ _12273_/A vssd1 vssd1 vccd1 vccd1 _12269_/Y sky130_fd_sc_hd__inv_2
X_14008_ _14008_/CLK _14008_/D vssd1 vssd1 vccd1 vccd1 _14008_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_7_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_110_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08500_ _08543_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _08502_/B sky130_fd_sc_hd__and2_1
XFILLER_48_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09480_ _08623_/B _09818_/B _09875_/A _08623_/A vssd1 vssd1 vccd1 vccd1 _09481_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_110_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08431_ _09361_/C vssd1 vssd1 vccd1 vccd1 _08449_/C sky130_fd_sc_hd__buf_2
XFILLER_93_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08362_ _08362_/A _08362_/B vssd1 vssd1 vccd1 vccd1 _08363_/C sky130_fd_sc_hd__xnor2_1
X_07313_ _14165_/D _07541_/B _07313_/C vssd1 vssd1 vccd1 vccd1 _07374_/A sky130_fd_sc_hd__and3_1
XANTENNA__08653__B1 _09000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08293_ _08622_/A _09962_/B _08318_/A _08292_/B vssd1 vssd1 vccd1 vccd1 _08295_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07244_ _14265_/Q _07243_/X _07253_/S vssd1 vssd1 vccd1 vccd1 _07245_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07175_ _07175_/A vssd1 vssd1 vccd1 vccd1 _14285_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12570__A _12576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07664__A _14068_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09816_ _10122_/A _10214_/A _09914_/A vssd1 vssd1 vccd1 vccd1 _09829_/B sky130_fd_sc_hd__o21ba_1
XFILLER_41_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09747_ _10524_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _10530_/A sky130_fd_sc_hd__nand2_2
XFILLER_36_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06959_ _06956_/X _14315_/Q _06959_/S vssd1 vssd1 vccd1 vccd1 _06960_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08495__A _13862_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09678_ _09678_/A _09678_/B _09678_/C vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__and3_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08629_/A vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__buf_4
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _13844_/Q _11639_/Y _11652_/S vssd1 vssd1 vccd1 vccd1 _11641_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ _11543_/Y _11614_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__o21ai_4
XFILLER_74_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13310_ _14343_/Q _13289_/X _13309_/X _13301_/X vssd1 vssd1 vccd1 vccd1 _14343_/D
+ sky130_fd_sc_hd__o211a_1
X_10522_ _10644_/A _10522_/B _10522_/C vssd1 vssd1 vccd1 vccd1 _10522_/X sky130_fd_sc_hd__or3_1
X_14290_ _14322_/CLK _14290_/D _13155_/Y vssd1 vssd1 vccd1 vccd1 _14290_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_7_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13241_ _14441_/Q _13201_/X _13204_/X _14393_/Q vssd1 vssd1 vccd1 vccd1 _13241_/X
+ sky130_fd_sc_hd__a22o_1
X_10453_ _10453_/A _10453_/B vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__nand2_1
XFILLER_108_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08947__A1 _08944_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input66_A io_wbs_datwr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13172_ _13178_/A vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__buf_2
X_10384_ _10384_/A _10351_/B vssd1 vssd1 vccd1 vccd1 _10384_/X sky130_fd_sc_hd__or2b_1
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12123_ _12940_/A _12130_/B vssd1 vssd1 vccd1 vccd1 _12123_/X sky130_fd_sc_hd__or2_1
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07080__C1 _14363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12054_ _12065_/A _12054_/B vssd1 vssd1 vccd1 vccd1 _12055_/A sky130_fd_sc_hd__and2_1
XFILLER_81_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11005_ _11005_/A _11005_/B vssd1 vssd1 vccd1 vccd1 _11070_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12956_ _12960_/A vssd1 vssd1 vccd1 vccd1 _12956_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11907_ _13817_/Q _11872_/A _11905_/X _11906_/Y hold38/X vssd1 vssd1 vccd1 vccd1
+ _13757_/D sky130_fd_sc_hd__o221a_1
XFILLER_61_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _12930_/A _12896_/B vssd1 vssd1 vccd1 vccd1 _12887_/X sky130_fd_sc_hd__or2_1
XFILLER_61_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11838_ _14337_/Q _11833_/X _11834_/X _13796_/Q _11837_/X vssd1 vssd1 vccd1 vccd1
+ _11838_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11769_ _12181_/A vssd1 vssd1 vccd1 vccd1 _13035_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13508_ _12673_/X _14399_/Q _13511_/S vssd1 vssd1 vccd1 vccd1 _13509_/B sky130_fd_sc_hd__mux2_1
X_13439_ _13439_/A vssd1 vssd1 vccd1 vccd1 _14378_/D sky130_fd_sc_hd__clkbuf_1
X_08980_ _08980_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _08981_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07931_ _14023_/Q vssd1 vssd1 vccd1 vccd1 _09145_/A sky130_fd_sc_hd__buf_2
XFILLER_111_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09363__A1 _09145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__B2 _09145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07862_ _07919_/S _07862_/B vssd1 vssd1 vccd1 vccd1 _07863_/B sky130_fd_sc_hd__or2_1
XFILLER_29_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09601_ _09601_/A _09601_/B _09601_/C vssd1 vssd1 vccd1 vccd1 _09676_/B sky130_fd_sc_hd__nand3_2
XFILLER_56_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07793_ _10951_/A vssd1 vssd1 vccd1 vccd1 _10648_/A sky130_fd_sc_hd__buf_2
X_09532_ _09465_/A _09513_/B _09511_/X vssd1 vssd1 vccd1 vccd1 _09582_/A sky130_fd_sc_hd__a21oi_2
XFILLER_97_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _09462_/A _09462_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _09464_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08414_ _08905_/A vssd1 vssd1 vccd1 vccd1 _09044_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09394_ _09390_/X _09392_/Y _09393_/A _09393_/Y vssd1 vssd1 vccd1 vccd1 _09396_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_40_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08345_ _13866_/Q vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__buf_2
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08276_ _08276_/A _08276_/B vssd1 vssd1 vccd1 vccd1 _08277_/B sky130_fd_sc_hd__or2_1
XFILLER_20_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07227_ _14270_/Q _07226_/X _07236_/S vssd1 vssd1 vccd1 vccd1 _07228_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14185__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07158_ _14105_/Q _07140_/X _07143_/X vssd1 vssd1 vccd1 vccd1 _07158_/X sky130_fd_sc_hd__a21o_1
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07089_ _14266_/Q _07085_/X _07088_/X _14362_/Q vssd1 vssd1 vccd1 vccd1 _07089_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08937__B _08937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ _14159_/Q _12801_/X _12803_/X _14143_/Q _12809_/X vssd1 vssd1 vccd1 vccd1
+ _12810_/X sky130_fd_sc_hd__a221o_1
XFILLER_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13790_ _13809_/CLK _13790_/D vssd1 vssd1 vccd1 vccd1 _13790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12753_/A vssd1 vssd1 vccd1 vccd1 _12746_/A sky130_fd_sc_hd__buf_2
XFILLER_27_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12672_ _12672_/A vssd1 vssd1 vccd1 vccd1 _14050_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14411_/CLK _14411_/D vssd1 vssd1 vccd1 vccd1 _14411_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11623_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11623_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_8_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14342_ _14348_/CLK _14342_/D vssd1 vssd1 vccd1 vccd1 _14342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ _14042_/Q _13954_/Q vssd1 vssd1 vccd1 vccd1 _11554_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12194__B _12900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10505_ _10505_/A _10505_/B vssd1 vssd1 vccd1 vccd1 _10506_/B sky130_fd_sc_hd__xnor2_1
X_14273_ _14275_/CLK _14273_/D _13133_/Y vssd1 vssd1 vccd1 vccd1 _14273_/Q sky130_fd_sc_hd__dfrtp_4
X_11485_ _10009_/A _11455_/X _11483_/X _11484_/X vssd1 vssd1 vccd1 vccd1 _13870_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13224_ _14325_/Q _13196_/X _13223_/X _13053_/X vssd1 vssd1 vccd1 vccd1 _14325_/D
+ sky130_fd_sc_hd__o211a_1
X_10436_ _10463_/S _10436_/B vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_output172_A _14297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ _13159_/A vssd1 vssd1 vccd1 vccd1 _13155_/Y sky130_fd_sc_hd__inv_2
X_10367_ _10367_/A _10367_/B vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _12930_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12106_/X sky130_fd_sc_hd__or2_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13677__A0 _12673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13086_ _13089_/A _13086_/B vssd1 vssd1 vccd1 vccd1 _13087_/A sky130_fd_sc_hd__and2_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10298_/A _10298_/B vssd1 vssd1 vccd1 vccd1 _10324_/B sky130_fd_sc_hd__nor2_2
X_12037_ _12037_/A vssd1 vssd1 vccd1 vccd1 _13793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ _13988_/CLK _13988_/D _12419_/Y vssd1 vssd1 vccd1 vccd1 _13988_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_65_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14058__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12939_ hold7/A _12928_/X _12938_/X _12934_/X vssd1 vssd1 vccd1 vccd1 _14162_/D sky130_fd_sc_hd__o211a_1
XFILLER_94_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08130_ _08130_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08131_/B sky130_fd_sc_hd__nor2_2
XFILLER_30_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08061_ _08251_/A _09234_/B _09233_/C _09084_/A vssd1 vssd1 vccd1 vccd1 _08061_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_105_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07012_ _07090_/A vssd1 vssd1 vccd1 vccd1 _07012_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09694__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08963_ _08778_/X _08779_/Y _08857_/Y _08961_/X _08962_/Y vssd1 vssd1 vccd1 vccd1
+ _08963_/X sky130_fd_sc_hd__a221o_1
XFILLER_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10352__B _10420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07914_ _07914_/A _07836_/Y vssd1 vssd1 vccd1 vccd1 _07915_/B sky130_fd_sc_hd__or2b_1
XFILLER_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08894_ _09055_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _08895_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07942__A _13869_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07845_ _14031_/Q _13977_/Q vssd1 vssd1 vccd1 vccd1 _07892_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07776_ _13987_/Q vssd1 vssd1 vccd1 vccd1 _07806_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07153__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ _09515_/A _09528_/B vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__xnor2_2
XFILLER_25_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09446_ _09545_/C _08291_/C _09489_/A _09445_/D vssd1 vssd1 vccd1 vccd1 _09447_/C
+ sky130_fd_sc_hd__a22o_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09377_ _09377_/A _09302_/A vssd1 vssd1 vccd1 vccd1 _09388_/A sky130_fd_sc_hd__or2b_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08328_ _08325_/X _08326_/Y _08380_/A _08324_/Y vssd1 vssd1 vccd1 vccd1 _08391_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08259_ _09771_/B _08259_/B vssd1 vssd1 vccd1 vccd1 _08262_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11270_ _11350_/A _11350_/B _11351_/B vssd1 vssd1 vccd1 vccd1 _11347_/B sky130_fd_sc_hd__o21ai_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10221_ _10213_/C _10214_/Y _10219_/Y _10220_/Y vssd1 vssd1 vccd1 vccd1 _10221_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _10285_/B _10153_/B vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__xnor2_2
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10083_ _10083_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__xnor2_1
XFILLER_102_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13911_ _13915_/CLK _13911_/D _12321_/Y vssd1 vssd1 vccd1 vccd1 _13911_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input29_A dout1[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13842_ _14275_/CLK _13842_/D _12235_/Y vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfrtp_1
XFILLER_63_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13773_ _14465_/CLK _13773_/D vssd1 vssd1 vccd1 vccd1 _13773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10985_ _11207_/A _10993_/A _10993_/B vssd1 vssd1 vccd1 vccd1 _10990_/B sky130_fd_sc_hd__o21a_1
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12724_ _12727_/A vssd1 vssd1 vccd1 vccd1 _12724_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08683__A _08937_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12655_ _12654_/X _14047_/Q _12665_/S vssd1 vssd1 vccd1 vccd1 _12656_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10718__A _11240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06915__B _14288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11606_ _11606_/A _11606_/B vssd1 vssd1 vccd1 vccd1 _11606_/Y sky130_fd_sc_hd__xnor2_4
X_12586_ _12611_/S vssd1 vssd1 vccd1 vccd1 _12600_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14325_ _14396_/CLK _14325_/D vssd1 vssd1 vccd1 vccd1 _14325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11537_ _14056_/Q _13968_/Q vssd1 vssd1 vccd1 vccd1 _11587_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14256_ _14256_/CLK hold11/X _13110_/Y vssd1 vssd1 vccd1 vccd1 _14256_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06931__A _06970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _11464_/X _11302_/A _11465_/Y _11466_/Y _11467_/Y vssd1 vssd1 vccd1 vccd1
+ _11468_/X sky130_fd_sc_hd__a221o_1
XFILLER_48_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13207_ _13328_/A vssd1 vssd1 vccd1 vccd1 _13236_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__08369__A2 _13874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ _10435_/A _10435_/B vssd1 vssd1 vccd1 vccd1 _10421_/A sky130_fd_sc_hd__xor2_1
X_14187_ _14256_/CLK _14187_/D _12975_/Y vssd1 vssd1 vccd1 vccd1 _14187_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11399_ _13844_/Q _11403_/B vssd1 vssd1 vccd1 vccd1 _11399_/X sky130_fd_sc_hd__or2_1
XFILLER_48_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _13140_/A vssd1 vssd1 vccd1 vccd1 _13138_/Y sky130_fd_sc_hd__inv_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_19_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14107_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _12579_/X _14243_/Q _13076_/S vssd1 vssd1 vccd1 vccd1 _13070_/B sky130_fd_sc_hd__mux2_1
XFILLER_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07630_ _14125_/Q _14060_/Q vssd1 vssd1 vccd1 vccd1 _07685_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07561_ _07561_/A vssd1 vssd1 vccd1 vccd1 _14101_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09300_ _09210_/A _09209_/B _09209_/A vssd1 vssd1 vccd1 vccd1 _09302_/B sky130_fd_sc_hd__o21bai_1
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08593__A _08867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07492_ _14230_/Q _07534_/B vssd1 vssd1 vccd1 vccd1 _07492_/Y sky130_fd_sc_hd__nor2_1
X_09231_ _09198_/A _09198_/Y _09229_/X _09230_/Y vssd1 vssd1 vccd1 vccd1 _09276_/A
+ sky130_fd_sc_hd__a211oi_2
X_09162_ _09177_/A vssd1 vssd1 vccd1 vccd1 _09198_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13050__A1 _14236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08113_ _08113_/A vssd1 vssd1 vccd1 vccd1 _08389_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ _08573_/B _09887_/A _08494_/D _08012_/A vssd1 vssd1 vccd1 vccd1 _09094_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_io_wbs_clk clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14449_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08044_ _08078_/A vssd1 vssd1 vccd1 vccd1 _08295_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__07937__A _13869_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13353__A2 _13265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10082__B _10092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _10346_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _09996_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08946_ _08946_/A _10206_/A vssd1 vssd1 vccd1 vccd1 _08946_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11116__A1 _11014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11906__B _11906_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _08877_/A vssd1 vssd1 vccd1 vccd1 _08887_/A sky130_fd_sc_hd__inv_2
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08487__B _09493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ _14028_/Q _13974_/Q vssd1 vssd1 vccd1 vccd1 _07839_/B sky130_fd_sc_hd__or2_1
XFILLER_45_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07759_ _07759_/A vssd1 vssd1 vccd1 vccd1 _14062_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11922__A _14228_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10770_ _10770_/A vssd1 vssd1 vccd1 vccd1 _10770_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09429_ _09364_/B _09364_/C _09364_/A vssd1 vssd1 vccd1 vccd1 _09430_/C sky130_fd_sc_hd__a21bo_1
X_12440_ _12440_/A _12440_/B vssd1 vssd1 vccd1 vccd1 _12441_/A sky130_fd_sc_hd__and2_1
XANTENNA__08008__A _13874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12371_ _12372_/A vssd1 vssd1 vccd1 vccd1 _12371_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14110_ _14239_/CLK _14110_/D vssd1 vssd1 vccd1 vccd1 _14110_/Q sky130_fd_sc_hd__dfxtp_1
X_11322_ _11322_/A vssd1 vssd1 vccd1 vccd1 _11322_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14041_ _14041_/CLK _14041_/D vssd1 vssd1 vccd1 vccd1 _14041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11253_ _11253_/A _11253_/B vssd1 vssd1 vccd1 vccd1 _11271_/B sky130_fd_sc_hd__xor2_2
XFILLER_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10204_ _10204_/A _10204_/B _10204_/C vssd1 vssd1 vccd1 vccd1 _10204_/Y sky130_fd_sc_hd__nand3_1
XFILLER_84_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11184_ _11142_/B _11169_/X _11184_/S vssd1 vssd1 vccd1 vccd1 _11184_/X sky130_fd_sc_hd__mux2_1
X_10135_ _10307_/A _10135_/B vssd1 vssd1 vccd1 vccd1 _10162_/B sky130_fd_sc_hd__xnor2_2
XFILLER_76_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10066_ _10069_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output135_A _11803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13825_ _13825_/CLK _13825_/D vssd1 vssd1 vccd1 vccd1 _13825_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_21_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12607__A1 _14035_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12928__A _12928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11815__C1 _11814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13756_ _13825_/CLK _13756_/D _11946_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Q sky130_fd_sc_hd__dfrtp_1
X_10968_ _10722_/B _10953_/B _10967_/X _10730_/B vssd1 vssd1 vccd1 vccd1 _10968_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _12709_/A vssd1 vssd1 vccd1 vccd1 _12707_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11551__B _13952_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13687_ _12561_/X _14450_/Q _13687_/S vssd1 vssd1 vccd1 vccd1 _13688_/B sky130_fd_sc_hd__mux2_1
X_10899_ _10899_/A _10899_/B vssd1 vssd1 vccd1 vccd1 _10899_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12638_ _12579_/X _14043_/Q _12642_/S vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__mux2_1
XFILLER_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12569_ _12218_/X _14024_/Q _12583_/S vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08860__B _10215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14308_ _14453_/CLK _14308_/D _13176_/Y vssd1 vssd1 vccd1 vccd1 _14308_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14239_ _14239_/CLK _14239_/D vssd1 vssd1 vccd1 vccd1 _14239_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11346__B2 _07784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09972__A _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08820_/B _08820_/C _08820_/A vssd1 vssd1 vccd1 vccd1 _08801_/C sky130_fd_sc_hd__a21bo_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09780_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09781_/C sky130_fd_sc_hd__xor2_4
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _06992_/A vssd1 vssd1 vccd1 vccd1 _14311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10911__A _13926_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08731_/A _08764_/A _08731_/C vssd1 vssd1 vccd1 vccd1 _08735_/A sky130_fd_sc_hd__nand3_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08662_ _09053_/A _09053_/B _09482_/B _08982_/B vssd1 vssd1 vccd1 vccd1 _08663_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_96_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07613_ _14077_/Q input12/X _07615_/S vssd1 vssd1 vccd1 vccd1 _07614_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08593_ _08867_/A _08703_/B vssd1 vssd1 vccd1 vccd1 _08600_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07544_ _14179_/Q _07526_/X _07543_/Y _07519_/X vssd1 vssd1 vccd1 vccd1 _14171_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12074__A2 _12059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07475_ _07483_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07475_/X sky130_fd_sc_hd__or2_1
XFILLER_50_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09214_ _09158_/B _09158_/C _09158_/A vssd1 vssd1 vccd1 vccd1 _09215_/C sky130_fd_sc_hd__a21bo_1
X_09145_ _09145_/A _09145_/B _09884_/A _09145_/D vssd1 vssd1 vccd1 vccd1 _09148_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__08498__A2_N _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12573__A _12576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09076_ _09164_/A _09076_/B _09076_/C vssd1 vssd1 vccd1 vccd1 _09079_/A sky130_fd_sc_hd__or3_1
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08027_ _09545_/C vssd1 vssd1 vccd1 vccd1 _08716_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_116_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11337__A1 _10826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09978_ _09978_/A _09978_/B vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__nor2_4
X_08929_ _08939_/A _08939_/B vssd1 vssd1 vccd1 vccd1 _08940_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13763__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11940_ _11940_/A vssd1 vssd1 vccd1 vccd1 _11940_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _11871_/A vssd1 vssd1 vccd1 vccd1 _11871_/X sky130_fd_sc_hd__clkbuf_1
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13625_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10822_ _10834_/B _10835_/B _10834_/A vssd1 vssd1 vccd1 vccd1 _10832_/B sky130_fd_sc_hd__o21ba_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09122__A _09336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ _13592_/A vssd1 vssd1 vccd1 vccd1 _13556_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10753_ _10719_/A _11240_/A _10753_/S vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11812__A2 _11848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13472_ _13522_/S vssd1 vssd1 vccd1 vccd1 _13475_/S sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input96_A io_wbs_datwr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10684_ _10684_/A vssd1 vssd1 vccd1 vccd1 _13947_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14269__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ input33/X input44/X vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__nor2_2
XFILLER_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08680__B _10486_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12354_ _12385_/A vssd1 vssd1 vccd1 vccd1 _12379_/A sky130_fd_sc_hd__clkbuf_4
X_11305_ _11457_/A _11305_/B vssd1 vssd1 vccd1 vccd1 _11305_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12285_ _12285_/A vssd1 vssd1 vccd1 vccd1 _12285_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14024_ _14275_/CLK _14024_/D vssd1 vssd1 vccd1 vccd1 _14024_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09792__A _09792_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11236_ _11236_/A _11236_/B vssd1 vssd1 vccd1 vccd1 _11237_/B sky130_fd_sc_hd__nor2_2
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11167_ _10771_/Y _11165_/X _11166_/X _10744_/A vssd1 vssd1 vccd1 vccd1 _11167_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10118_ _10118_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10119_/B sky130_fd_sc_hd__xor2_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11098_ _10831_/X _11084_/X _11097_/Y _10675_/X _11082_/A vssd1 vssd1 vccd1 vccd1
+ _13925_/D sky130_fd_sc_hd__a32o_1
X_10049_ _10124_/B _10050_/B vssd1 vssd1 vccd1 vccd1 _10056_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09016__B _09084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__A1 _11014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13808_ _13809_/CLK _13808_/D vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfxtp_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13253__A1 _14363_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13739_ _13745_/A _13739_/B vssd1 vssd1 vccd1 vccd1 _13740_/A sky130_fd_sc_hd__and2_1
XFILLER_56_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07260_ _07260_/A vssd1 vssd1 vccd1 vccd1 _14260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07191_ _14096_/Q _07185_/X _07186_/X vssd1 vssd1 vccd1 vccd1 _07191_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_9_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14281_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12516__A0 _12515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09901_ _10435_/A _09901_/B vssd1 vssd1 vccd1 vccd1 _09938_/A sky130_fd_sc_hd__xor2_2
XFILLER_116_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09832_ _09801_/A _10048_/A _09801_/B vssd1 vssd1 vccd1 vccd1 _10436_/B sky130_fd_sc_hd__a21bo_2
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__A1 hold3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _10578_/A vssd1 vssd1 vccd1 vccd1 _10528_/A sky130_fd_sc_hd__clkinv_2
XFILLER_101_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06975_ _06973_/X _06974_/X _14377_/Q vssd1 vssd1 vccd1 vccd1 _06976_/S sky130_fd_sc_hd__o21a_1
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__B2 _14147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08714_ _09084_/C vssd1 vssd1 vccd1 vccd1 _08925_/C sky130_fd_sc_hd__buf_2
XFILLER_6_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08468__D _08703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09694_ _09694_/A _09731_/B vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07950__A _14021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ _08645_/A _08645_/B _08645_/C vssd1 vssd1 vccd1 vccd1 _08675_/B sky130_fd_sc_hd__and3_2
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07171__A1 _07169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12568__A _12611_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08576_ _08576_/A _08576_/B vssd1 vssd1 vccd1 vccd1 _08643_/A sky130_fd_sc_hd__xnor2_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07527_ _14175_/Q _07534_/A _14176_/Q vssd1 vssd1 vccd1 vccd1 _07528_/B sky130_fd_sc_hd__o21a_1
XANTENNA__10088__A _10126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07458_ _07458_/A _07458_/B vssd1 vssd1 vccd1 vccd1 _07458_/X sky130_fd_sc_hd__or2_1
XFILLER_109_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07389_ _14212_/Q _07373_/X _07375_/X _07388_/X vssd1 vssd1 vccd1 vccd1 _14212_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11411__S _11415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09128_ _09127_/A _09127_/C _09127_/B vssd1 vssd1 vccd1 vccd1 _09130_/B sky130_fd_sc_hd__o21ai_1
XFILLER_68_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10230__A1 _10271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09059_ _09508_/B _09218_/B _09875_/A _08445_/X vssd1 vssd1 vccd1 vccd1 _09060_/C
+ sky130_fd_sc_hd__a22o_2
X_12070_ _12070_/A vssd1 vssd1 vccd1 vccd1 _13801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11021_ _11021_/A _11021_/B vssd1 vssd1 vccd1 vccd1 _11058_/B sky130_fd_sc_hd__xnor2_1
XFILLER_103_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09117__A _10632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12972_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12972_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13483__A1 _12911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input11_A dout1[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _14229_/Q _14192_/Q vssd1 vssd1 vccd1 vccd1 _14168_/D sky130_fd_sc_hd__xnor2_2
XFILLER_57_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07162__A1 _07161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _14347_/Q _11808_/X _11823_/X _13806_/Q vssd1 vssd1 vccd1 vccd1 _11854_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__B2 _14392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _10868_/B _10874_/A _10868_/A vssd1 vssd1 vccd1 vccd1 _10869_/A sky130_fd_sc_hd__o21a_1
X_11785_ _11785_/A _11785_/B vssd1 vssd1 vccd1 vccd1 _11786_/A sky130_fd_sc_hd__or2_4
X_13524_ _13524_/A vssd1 vssd1 vccd1 vccd1 _14403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10736_ _10761_/C _10735_/X _10748_/A vssd1 vssd1 vccd1 vccd1 _10737_/S sky130_fd_sc_hd__o21ai_1
XFILLER_15_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13455_ _13461_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__and2_1
XFILLER_51_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10667_ _10916_/A vssd1 vssd1 vccd1 vccd1 _11152_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ _12409_/A vssd1 vssd1 vccd1 vccd1 _12406_/Y sky130_fd_sc_hd__inv_2
X_13386_ _13392_/A _13386_/B vssd1 vssd1 vccd1 vccd1 _13387_/A sky130_fd_sc_hd__and2_1
X_10598_ _10598_/A _10598_/B _10598_/C vssd1 vssd1 vccd1 vccd1 _10598_/X sky130_fd_sc_hd__and3_1
X_12337_ _12341_/A vssd1 vssd1 vccd1 vccd1 _12337_/Y sky130_fd_sc_hd__inv_2
Xoutput108 _14067_/Q vssd1 vssd1 vccd1 vccd1 addr1[7] sky130_fd_sc_hd__buf_2
XFILLER_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput119 _11842_/X vssd1 vssd1 vccd1 vccd1 io_wbs_datrd[15] sky130_fd_sc_hd__buf_2
XANTENNA__06976__A1 _14313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ _12286_/A vssd1 vssd1 vccd1 vccd1 _12273_/A sky130_fd_sc_hd__clkbuf_2
X_14007_ _14441_/CLK _14007_/D vssd1 vssd1 vccd1 vccd1 _14007_/Q sky130_fd_sc_hd__dfxtp_2
X_11219_ _13905_/Q vssd1 vssd1 vccd1 vccd1 _11294_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12199_ _12213_/A _13042_/B vssd1 vssd1 vccd1 vccd1 _12205_/B sky130_fd_sc_hd__nor2_1
XFILLER_96_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13474__A1 _12209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07153__A1 _07144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08430_ _09869_/A vssd1 vssd1 vccd1 vccd1 _09361_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_17_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08361_ _09434_/A _09445_/B vssd1 vssd1 vccd1 vccd1 _08362_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07312_ _07312_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07541_/B sky130_fd_sc_hd__nand2_1
X_08292_ _08292_/A _08292_/B vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08653__B2 _08983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07243_ _14081_/Q _13881_/Q _07252_/S vssd1 vssd1 vccd1 vccd1 _07243_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07174_ _14285_/Q _07173_/X _07183_/S vssd1 vssd1 vccd1 vccd1 _07175_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07945__A _14021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07156__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _10271_/B _09913_/B vssd1 vssd1 vccd1 vccd1 _09914_/A sky130_fd_sc_hd__nor2_1
XANTENNA_input3_A dout1[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10090__B _10090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09746_ _09751_/C _08407_/B _08407_/C vssd1 vssd1 vccd1 vccd1 _09747_/B sky130_fd_sc_hd__o21ai_1
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06958_ _06934_/X _06957_/X _14379_/Q vssd1 vssd1 vccd1 vccd1 _06959_/S sky130_fd_sc_hd__o21a_1
XFILLER_74_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09677_ _09678_/A _09678_/B _09678_/C vssd1 vssd1 vccd1 vccd1 _09677_/Y sky130_fd_sc_hd__a21oi_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _14394_/Q _13781_/Q vssd1 vssd1 vccd1 vccd1 _06889_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07144__A1 _14107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08628_ _09434_/A _10081_/A _08575_/B _08573_/X vssd1 vssd1 vccd1 vccd1 _08636_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08559_/A _08559_/B vssd1 vssd1 vccd1 vccd1 _08561_/A sky130_fd_sc_hd__xnor2_1
XFILLER_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13621__S _13628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11570_ _14050_/Q _13962_/Q vssd1 vssd1 vccd1 vccd1 _11613_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10521_ _10520_/A _10520_/B _10520_/C vssd1 vssd1 vccd1 vccd1 _10522_/C sky130_fd_sc_hd__a21oi_1
XFILLER_109_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _13265_/A vssd1 vssd1 vccd1 vccd1 _13240_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10452_ _10493_/A _10452_/B vssd1 vssd1 vccd1 vccd1 _10453_/B sky130_fd_sc_hd__or2_1
XANTENNA__08016__A _13875_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ _13171_/A vssd1 vssd1 vccd1 vccd1 _13171_/Y sky130_fd_sc_hd__inv_2
X_10383_ _10383_/A _10396_/A vssd1 vssd1 vccd1 vccd1 _10386_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__14307__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12122_ input71/X vssd1 vssd1 vccd1 vccd1 _12940_/A sky130_fd_sc_hd__buf_6
XANTENNA__07855__A _14036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input59_A io_wbs_adr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12053_ _13797_/Q _12038_/X _12039_/X _13813_/Q vssd1 vssd1 vccd1 vccd1 _12054_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11004_ _11228_/A _11008_/A _11008_/B vssd1 vssd1 vccd1 vccd1 _11005_/B sky130_fd_sc_hd__o21ai_1
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13592__A _13592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12955_ _12973_/A vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__buf_2
XFILLER_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07135__A1 _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06918__B _06942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11906_ _13757_/Q _11906_/B vssd1 vssd1 vccd1 vccd1 _11906_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12001__A _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12886_ _12898_/B vssd1 vssd1 vccd1 vccd1 _12896_/B sky130_fd_sc_hd__clkbuf_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11837_ _14002_/Q _11797_/A _11830_/X _14121_/Q vssd1 vssd1 vccd1 vccd1 _11837_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10690__A1 _11533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12936__A _12936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11768_ _11768_/A _12762_/C vssd1 vssd1 vccd1 vccd1 _12181_/A sky130_fd_sc_hd__nor2_1
XFILLER_105_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06934__A _06973_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12431__A2 _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09310__A _09508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13507_ _13507_/A vssd1 vssd1 vccd1 vccd1 _14398_/D sky130_fd_sc_hd__clkbuf_1
X_10719_ _10719_/A vssd1 vssd1 vccd1 vccd1 _10746_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11699_ _13756_/Q _11902_/B vssd1 vssd1 vccd1 vccd1 _11906_/B sky130_fd_sc_hd__or2_2
X_13438_ _13444_/A _13438_/B vssd1 vssd1 vccd1 vccd1 _13439_/A sky130_fd_sc_hd__and2_1
XANTENNA__08938__A2 _08941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ _13375_/A _13369_/B vssd1 vssd1 vccd1 vccd1 _13370_/A sky130_fd_sc_hd__and2_1
XFILLER_115_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ _10547_/A vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__buf_4
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07861_ _14039_/Q _07861_/B vssd1 vssd1 vccd1 vccd1 _07862_/B sky130_fd_sc_hd__xnor2_1
XFILLER_111_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09600_ _09560_/A _09560_/C _09560_/B vssd1 vssd1 vccd1 vccd1 _09601_/C sky130_fd_sc_hd__a21bo_1
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07792_ _10758_/A vssd1 vssd1 vccd1 vccd1 _10951_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__13824__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08596__A _13866_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09531_ _09629_/A _09581_/B vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07126__A1 _14289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09462_ _09462_/A _09462_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _09464_/A sky130_fd_sc_hd__nand3_1
XFILLER_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08413_ _08941_/A vssd1 vssd1 vccd1 vccd1 _08905_/A sky130_fd_sc_hd__buf_2
X_09393_ _09393_/A _09393_/B _09393_/C vssd1 vssd1 vccd1 vccd1 _09393_/Y sky130_fd_sc_hd__nand3_1
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08344_ _09425_/A _09848_/A _08313_/A _08312_/D vssd1 vssd1 vccd1 vccd1 _08353_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08275_ _08276_/A _08276_/B vssd1 vssd1 vccd1 vccd1 _08277_/A sky130_fd_sc_hd__nand2_1
X_07226_ _14086_/Q _13886_/Q _07235_/S vssd1 vssd1 vccd1 vccd1 _07226_/X sky130_fd_sc_hd__mux2_2
XANTENNA_clkbuf_leaf_28_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_106_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07157_ _07157_/A vssd1 vssd1 vccd1 vccd1 _14290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07088_ _14410_/Q _07086_/Y _07087_/X vssd1 vssd1 vccd1 vccd1 _07088_/X sky130_fd_sc_hd__a21o_1
XFILLER_65_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08937__C _08937_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _09729_/A _09729_/B _09729_/C vssd1 vssd1 vccd1 vccd1 _09729_/X sky130_fd_sc_hd__or3_2
XFILLER_41_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ _12740_/A vssd1 vssd1 vccd1 vccd1 _12740_/Y sky130_fd_sc_hd__inv_2
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12671_ _12678_/A _12671_/B vssd1 vssd1 vccd1 vccd1 _12672_/A sky130_fd_sc_hd__and2_1
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14410_/CLK _14410_/D vssd1 vssd1 vccd1 vccd1 _14410_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11622_ _11544_/Y _11622_/B vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__and2b_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14341_ _14348_/CLK _14341_/D vssd1 vssd1 vccd1 vccd1 _14341_/Q sky130_fd_sc_hd__dfxtp_1
X_11553_ _11650_/B _11651_/B _11650_/A vssd1 vssd1 vccd1 vccd1 _11647_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__10276__A _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10504_ _09999_/Y _10395_/A _10000_/Y vssd1 vssd1 vccd1 vccd1 _10505_/B sky130_fd_sc_hd__a21oi_4
X_14272_ _14275_/CLK _14272_/D _13132_/Y vssd1 vssd1 vccd1 vccd1 _14272_/Q sky130_fd_sc_hd__dfrtp_4
X_11484_ _11002_/B _11460_/X _11475_/X _11294_/A _11461_/X vssd1 vssd1 vccd1 vccd1
+ _11484_/X sky130_fd_sc_hd__o221a_1
XFILLER_6_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13374__A0 _12641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13223_ hold33/A _13215_/X _13220_/X _13222_/X vssd1 vssd1 vccd1 vccd1 _13223_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ _10435_/A _10435_/B vssd1 vssd1 vccd1 vccd1 _10438_/B sky130_fd_sc_hd__nor2_1
XFILLER_100_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11924__A1 _14208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ _13178_/A vssd1 vssd1 vccd1 vccd1 _13159_/A sky130_fd_sc_hd__clkbuf_4
X_10366_ _10366_/A _10317_/B vssd1 vssd1 vccd1 vccd1 _10369_/B sky130_fd_sc_hd__or2b_1
XFILLER_88_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output165_A _14320_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12105_ input67/X vssd1 vssd1 vccd1 vccd1 _12930_/A sky130_fd_sc_hd__buf_4
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13084_/X hold34/A _13096_/S vssd1 vssd1 vccd1 vccd1 _13086_/B sky130_fd_sc_hd__mux2_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10297_ _10297_/A _10297_/B _10297_/C vssd1 vssd1 vccd1 vccd1 _10298_/B sky130_fd_sc_hd__and3_1
X_12036_ _12044_/A _12036_/B vssd1 vssd1 vccd1 vccd1 _12037_/A sky130_fd_sc_hd__and2_1
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_30_io_wbs_clk_A clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13997__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__B _13954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A1 _14296_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13987_ _13987_/CLK _13987_/D _12415_/Y vssd1 vssd1 vccd1 vccd1 _13987_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12938_ _12938_/A _12940_/B vssd1 vssd1 vccd1 vccd1 _12938_/X sky130_fd_sc_hd__or2_1
XFILLER_46_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _14136_/Q _12857_/X _12868_/X _12866_/X vssd1 vssd1 vccd1 vccd1 _14136_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08863__B _09241_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10186__A _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_48_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13825_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__07292__A0 _14241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08060_ _09796_/A vssd1 vssd1 vccd1 vccd1 _09233_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_31_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12168__A1 _13828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13365__A0 _13084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07011_ _14276_/Q _07007_/X _07010_/X _14372_/Q vssd1 vssd1 vccd1 vccd1 _07011_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08962_ _08962_/A _08962_/B vssd1 vssd1 vccd1 vccd1 _08962_/Y sky130_fd_sc_hd__nor2_1
XFILLER_102_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07913_ _07913_/A vssd1 vssd1 vccd1 vccd1 _13973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08893_ _08893_/A vssd1 vssd1 vccd1 vccd1 _08941_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_57_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07844_ _07896_/A _07897_/A _07843_/Y vssd1 vssd1 vccd1 vccd1 _07893_/A sky130_fd_sc_hd__o21a_1
XFILLER_111_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07775_ _13988_/Q vssd1 vssd1 vccd1 vccd1 _10655_/A sky130_fd_sc_hd__clkbuf_2
X_09514_ _09514_/A _09514_/B vssd1 vssd1 vccd1 vccd1 _09528_/B sky130_fd_sc_hd__xnor2_2
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09445_ _09545_/C _09445_/B _09489_/A _09445_/D vssd1 vssd1 vccd1 vccd1 _09489_/B
+ sky130_fd_sc_hd__nand4_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12576__A _12576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _09376_/A _09376_/B _09376_/C vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__nand3_1
XFILLER_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08712__A2_N _09942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08327_ _08380_/A _08324_/Y _08325_/X _08326_/Y vssd1 vssd1 vccd1 vccd1 _08391_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_32_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08258_ _08258_/A _08258_/B vssd1 vssd1 vccd1 vccd1 _08259_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07209_ _14091_/Q _13891_/Q _07218_/S vssd1 vssd1 vccd1 vccd1 _07209_/X sky130_fd_sc_hd__mux2_2
X_08189_ _09673_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08192_/B sky130_fd_sc_hd__xnor2_1
X_10220_ _10220_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10220_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13200__A _13206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ _10151_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _10151_/X sky130_fd_sc_hd__xor2_1
XFILLER_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10082_ _10092_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10083_/B sky130_fd_sc_hd__xnor2_1
XFILLER_43_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13910_ _13950_/CLK _13910_/D _12320_/Y vssd1 vssd1 vccd1 vccd1 _13910_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09125__A _09349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ _14028_/CLK _13841_/D _12233_/Y vssd1 vssd1 vccd1 vccd1 _13841_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13772_ _13825_/CLK _13772_/D _11965_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Q sky130_fd_sc_hd__dfrtp_2
X_10984_ _10999_/B _11000_/A _10997_/A _11207_/A vssd1 vssd1 vccd1 vccd1 _10993_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_74_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12723_ _12727_/A vssd1 vssd1 vccd1 vccd1 _12723_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12486__A _12486_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12654_ input95/X vssd1 vssd1 vccd1 vccd1 _12654_/X sky130_fd_sc_hd__buf_4
XFILLER_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _11541_/Y _11605_/B vssd1 vssd1 vccd1 vccd1 _11606_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12585_ _12585_/A vssd1 vssd1 vccd1 vccd1 _14028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14324_ _14396_/CLK _14324_/D vssd1 vssd1 vccd1 vccd1 _14324_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11536_ _11536_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09795__A _13871_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14255_ _14256_/CLK hold15/X _13109_/Y vssd1 vssd1 vccd1 vccd1 _14255_/Q sky130_fd_sc_hd__dfrtp_1
X_11467_ _11467_/A _11533_/S vssd1 vssd1 vccd1 vccd1 _11467_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13206_ _13206_/A _13359_/A vssd1 vssd1 vccd1 vccd1 _13328_/A sky130_fd_sc_hd__nand2_4
XANTENNA__13110__A _13115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10418_ _10418_/A _10564_/C vssd1 vssd1 vccd1 vccd1 _10418_/X sky130_fd_sc_hd__or2_1
X_14186_ _14256_/CLK _14186_/D _12974_/Y vssd1 vssd1 vccd1 vccd1 _14186_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11549__B _13954_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11398_ _13881_/Q _11392_/X _11396_/X _11397_/X vssd1 vssd1 vccd1 vccd1 _13881_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13137_ _13140_/A vssd1 vssd1 vccd1 vccd1 _13137_/Y sky130_fd_sc_hd__inv_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10349_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10360_/A sky130_fd_sc_hd__nor2_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09318__A2 _08091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ _13068_/A vssd1 vssd1 vccd1 vccd1 _14242_/D sky130_fd_sc_hd__clkbuf_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12019_ _12019_/A vssd1 vssd1 vccd1 vccd1 _13788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07560_ _14101_/Q input18/X _07560_/S vssd1 vssd1 vccd1 vccd1 _07561_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07491_ _07491_/A vssd1 vssd1 vccd1 vccd1 _07534_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08593__B _08703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09230_ _09277_/A _09277_/C _09277_/B vssd1 vssd1 vccd1 vccd1 _09230_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13586__A0 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09161_ _09161_/A _09161_/B _09161_/C vssd1 vssd1 vccd1 vccd1 _09177_/A sky130_fd_sc_hd__nand3_1
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08112_ _09514_/A _08116_/B _08110_/X vssd1 vssd1 vccd1 vccd1 _08113_/A sky130_fd_sc_hd__o21bai_4
X_09092_ _09153_/A _09153_/B _09092_/C _09092_/D vssd1 vssd1 vccd1 vccd1 _09094_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08043_ _08043_/A _09596_/A vssd1 vssd1 vccd1 vccd1 _08078_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10644__A _10644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13020__A _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09994_ _09994_/A _09994_/B vssd1 vssd1 vccd1 vccd1 _09995_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07953__A _09793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ _10171_/A vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__buf_2
XANTENNA__11116__A2 _11110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08876_ _08880_/A _08880_/B _08875_/X vssd1 vssd1 vccd1 vccd1 _08877_/A sky130_fd_sc_hd__o21ai_1
XFILLER_111_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07827_ _14028_/Q _13974_/Q vssd1 vssd1 vccd1 vccd1 _07840_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12077__B1 _12021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ _14062_/Q _07757_/X _07761_/S vssd1 vssd1 vccd1 vccd1 _07759_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07689_ _14133_/Q _07763_/A _07686_/Y _07687_/Y _07688_/Y vssd1 vssd1 vccd1 vccd1
+ _07689_/X sky130_fd_sc_hd__o311a_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09428_ _09427_/A _09427_/C _09427_/B vssd1 vssd1 vccd1 vccd1 _09430_/B sky130_fd_sc_hd__o21ai_1
X_09359_ _09626_/B _09359_/B vssd1 vssd1 vccd1 vccd1 _09360_/B sky130_fd_sc_hd__xor2_2
XFILLER_40_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07256__A0 _14261_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12370_ _12372_/A vssd1 vssd1 vccd1 vccd1 _12370_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11321_ _11321_/A _11321_/B vssd1 vssd1 vccd1 vccd1 _11321_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_10_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ _14041_/CLK _14040_/D vssd1 vssd1 vccd1 vccd1 _14040_/Q sky130_fd_sc_hd__dfxtp_1
X_11252_ _11252_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11253_/B sky130_fd_sc_hd__or2_1
XFILLER_69_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10203_ _10205_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10204_/C sky130_fd_sc_hd__or2b_1
XFILLER_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ _11244_/B _11245_/A vssd1 vssd1 vccd1 vccd1 _11240_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10134_ _10122_/Y _10123_/Y _10124_/Y vssd1 vssd1 vccd1 vccd1 _10307_/A sky130_fd_sc_hd__a21o_1
XANTENNA_input41_A io_wbs_adr[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09781__C _09781_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__A0 _12664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10065_ _10065_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__and2_1
XFILLER_47_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12068__B1 _12060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13824_ _13825_/CLK _13824_/D vssd1 vssd1 vccd1 vccd1 _13824_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_47_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08694__A _09349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967_ _13899_/Q _13900_/Q _10967_/S vssd1 vssd1 vccd1 vccd1 _10967_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13755_ _13826_/CLK _13755_/D _11945_/Y vssd1 vssd1 vccd1 vccd1 _13755_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _12709_/A vssd1 vssd1 vccd1 vccd1 _12706_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13686_ _13686_/A vssd1 vssd1 vccd1 vccd1 _14449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10898_ _10898_/A vssd1 vssd1 vccd1 vccd1 _13930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12637_ _12637_/A vssd1 vssd1 vccd1 vccd1 _12656_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12944__A _13010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09238__B1_N _09127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07247__A0 _14264_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12568_ _12611_/S vssd1 vssd1 vccd1 vccd1 _12583_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_102_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11519_ _11054_/A _11513_/X _11499_/X _11273_/A _11514_/X vssd1 vssd1 vccd1 vccd1
+ _11519_/X sky130_fd_sc_hd__o221a_1
X_14307_ _14417_/CLK _14307_/D _13175_/Y vssd1 vssd1 vccd1 vccd1 _14307_/Q sky130_fd_sc_hd__dfrtp_4
X_12499_ _14003_/Q _12481_/X _12497_/X _12498_/X vssd1 vssd1 vccd1 vccd1 _14003_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11279__B _11279_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14238_ _14239_/CLK _14238_/D vssd1 vssd1 vccd1 vccd1 _14238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14169_ _14283_/CLK _14169_/D _12950_/Y vssd1 vssd1 vccd1 vccd1 _14169_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _06987_/X _14311_/Q _06991_/S vssd1 vssd1 vccd1 vccd1 _06992_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _08566_/B _08566_/C _08566_/A vssd1 vssd1 vccd1 vccd1 _08731_/C sky130_fd_sc_hd__a21o_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08661_ _08468_/B _09482_/B _09434_/B _08925_/A vssd1 vssd1 vccd1 vccd1 _08663_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_96_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07612_ _07612_/A vssd1 vssd1 vccd1 vccd1 _14078_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08592_ _08592_/A _08592_/B vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__nand2_1
XFILLER_54_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07543_ _14171_/Q _07543_/B vssd1 vssd1 vccd1 vccd1 _07543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13271__A2 _13306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07486__B1 _07460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _14195_/Q _14197_/Q _07482_/S vssd1 vssd1 vccd1 vccd1 _07475_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13559__A0 _12664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08109__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ _09212_/A _09212_/C _09212_/B vssd1 vssd1 vccd1 vccd1 _09215_/B sky130_fd_sc_hd__a21o_1
XFILLER_10_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09144_ _09144_/A _09144_/B _09144_/C vssd1 vssd1 vccd1 vccd1 _09144_/Y sky130_fd_sc_hd__nand3_1
XFILLER_108_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09075_ _08580_/B _09811_/B _08629_/A _09493_/A vssd1 vssd1 vccd1 vccd1 _09076_/C
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__07159__S _07165_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ _09297_/A vssd1 vssd1 vccd1 vccd1 _09545_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_104_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ _10090_/A _09930_/B _10039_/A vssd1 vssd1 vccd1 vccd1 _09978_/B sky130_fd_sc_hd__a21oi_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08928_ _08928_/A _08928_/B vssd1 vssd1 vccd1 vccd1 _08939_/B sky130_fd_sc_hd__or2_1
XFILLER_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08859_ _08859_/A _08859_/B vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__xnor2_1
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07713__A1 hold7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13624__S _13628_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11933__A _13153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ _14355_/Q _11870_/B vssd1 vssd1 vccd1 vccd1 _11871_/A sky130_fd_sc_hd__and2_1
XFILLER_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10821_ _10716_/B _10727_/C _10716_/A vssd1 vssd1 vccd1 vccd1 _10834_/A sky130_fd_sc_hd__a21oi_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13540_ _13540_/A vssd1 vssd1 vccd1 vccd1 _14407_/D sky130_fd_sc_hd__clkbuf_1
X_10752_ _10730_/A _10744_/X _10748_/X vssd1 vssd1 vccd1 vccd1 _10753_/S sky130_fd_sc_hd__a21bo_1
XFILLER_38_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _13497_/A vssd1 vssd1 vccd1 vccd1 _13522_/S sky130_fd_sc_hd__buf_2
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ _10826_/A _11110_/A _10730_/A vssd1 vssd1 vccd1 vccd1 _10684_/A sky130_fd_sc_hd__mux2_1
XANTENNA__07229__A0 _14085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11025__A1 _11244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ _12460_/A vssd1 vssd1 vccd1 vccd1 _12422_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07858__A _14038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input89_A io_wbs_datwr[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08977__B1 _09482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12353_ _12353_/A vssd1 vssd1 vccd1 vccd1 _12353_/Y sky130_fd_sc_hd__inv_2
X_11304_ _11315_/B _11315_/C _11315_/A vssd1 vssd1 vccd1 vccd1 _11312_/B sky130_fd_sc_hd__a21o_1
XFILLER_107_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12284_ _12285_/A vssd1 vssd1 vccd1 vccd1 _12284_/Y sky130_fd_sc_hd__inv_2
X_14023_ _14304_/CLK _14023_/D vssd1 vssd1 vccd1 vccd1 _14023_/Q sky130_fd_sc_hd__dfxtp_2
X_11235_ _13901_/Q vssd1 vssd1 vccd1 vccd1 _11282_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07401__A0 _14208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ _13916_/Q _13917_/Q _13918_/Q _13919_/Q _10960_/S _10662_/A vssd1 vssd1 vccd1
+ vccd1 _11166_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10117_ _10079_/A _10078_/B _10076_/Y vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__a21oi_1
XFILLER_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11097_ _11083_/X _11097_/B _11097_/C vssd1 vssd1 vccd1 vccd1 _11097_/Y sky130_fd_sc_hd__nand3b_1
XFILLER_49_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10048_ _10048_/A _10048_/B vssd1 vssd1 vccd1 vccd1 _10351_/B sky130_fd_sc_hd__xor2_4
XFILLER_82_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07704__A1 _07548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13807_ _13809_/CLK _13807_/D vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13253__A2 _13215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11999_ _11999_/A vssd1 vssd1 vccd1 vccd1 _13783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13738_ input87/X _14465_/Q _13738_/S vssd1 vssd1 vccd1 vccd1 _13739_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13669_ _13669_/A vssd1 vssd1 vccd1 vccd1 _14444_/D sky130_fd_sc_hd__clkbuf_1
X_07190_ _07190_/A vssd1 vssd1 vccd1 vccd1 _14281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12516__A1 _08683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09900_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09990_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10010__A2_N _10127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08196__A1 _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _10435_/B _09829_/B _09830_/X vssd1 vssd1 vccd1 vccd1 _09921_/A sky130_fd_sc_hd__o21ai_2
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ _14425_/Q _06981_/B _14457_/Q vssd1 vssd1 vccd1 vccd1 _06974_/X sky130_fd_sc_hd__and3b_1
X_09762_ _09762_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09762_/Y sky130_fd_sc_hd__nor2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__A2 _12772_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08713_/A _08713_/B vssd1 vssd1 vccd1 vccd1 _08742_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09693_ _08389_/A _09685_/B _09684_/A vssd1 vssd1 vccd1 vccd1 _09731_/B sky130_fd_sc_hd__a21oi_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12849__A _13072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11753__A _11753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ _08997_/A _08997_/B vssd1 vssd1 vccd1 vccd1 _08645_/C sky130_fd_sc_hd__or2_1
XFILLER_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09223__A _09223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08575_ _08573_/X _08575_/B vssd1 vssd1 vccd1 vccd1 _08576_/B sky130_fd_sc_hd__and2b_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07526_ _07543_/B vssd1 vssd1 vccd1 vccd1 _07526_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07457_ _14198_/Q _14200_/Q _07469_/S vssd1 vssd1 vccd1 vccd1 _07458_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09877__B _10067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07388_ _07376_/X _07386_/X _07387_/X _07379_/X vssd1 vssd1 vccd1 vccd1 _07388_/X
+ sky130_fd_sc_hd__a22o_1
X_09127_ _09127_/A _09127_/B _09127_/C vssd1 vssd1 vccd1 vccd1 _09130_/A sky130_fd_sc_hd__or3_1
XFILLER_68_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09058_ _09234_/A _09058_/B vssd1 vssd1 vccd1 vccd1 _09060_/B sky130_fd_sc_hd__and2_1
XFILLER_117_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13704__A0 input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08009_ _09545_/D vssd1 vssd1 vccd1 vccd1 _08208_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_117_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11928__A input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11020_ _11020_/A _11020_/B vssd1 vssd1 vccd1 vccd1 _11021_/B sky130_fd_sc_hd__or2_1
XFILLER_1_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08302__A _09336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09117__B _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12971_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12971_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11663__A _11920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ _14228_/Q _14225_/Q vssd1 vssd1 vccd1 vccd1 _14167_/D sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_35_io_wbs_clk_A clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _14346_/Q _11847_/X _11848_/X _13805_/Q vssd1 vssd1 vccd1 vccd1 _11853_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__A2 _13201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _10863_/B _10804_/B vssd1 vssd1 vccd1 vccd1 _10868_/A sky130_fd_sc_hd__nor2_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ _14324_/Q _13194_/A _12192_/A _13833_/Q _11783_/X vssd1 vssd1 vccd1 vccd1
+ _11785_/B sky130_fd_sc_hd__a221o_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _13539_/A _13523_/B vssd1 vssd1 vccd1 vccd1 _13524_/A sky130_fd_sc_hd__and2_1
XFILLER_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10735_ _11181_/A vssd1 vssd1 vccd1 vccd1 _10735_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10666_ _10950_/S vssd1 vssd1 vccd1 vccd1 _10916_/A sky130_fd_sc_hd__inv_2
X_13454_ input85/X _14383_/Q _13460_/S vssd1 vssd1 vccd1 vccd1 _13455_/B sky130_fd_sc_hd__mux2_1
XFILLER_90_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12405_ _12409_/A vssd1 vssd1 vccd1 vccd1 _12405_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13385_ _12654_/X _14363_/Q _13391_/S vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__mux2_1
X_10597_ _10597_/A _10597_/B _10597_/C vssd1 vssd1 vccd1 vccd1 _10597_/X sky130_fd_sc_hd__or3_1
XFILLER_12_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12336_ _12348_/A vssd1 vssd1 vccd1 vccd1 _12341_/A sky130_fd_sc_hd__buf_2
Xoutput109 _14068_/Q vssd1 vssd1 vccd1 vccd1 addr1[8] sky130_fd_sc_hd__buf_2
XFILLER_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13529__S _13542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ _12267_/A vssd1 vssd1 vccd1 vccd1 _12267_/Y sky130_fd_sc_hd__inv_2
X_11218_ _11297_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11317_/B sky130_fd_sc_hd__and2_1
X_14006_ _14442_/CLK _14006_/D vssd1 vssd1 vccd1 vccd1 _14006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12198_ _13079_/A vssd1 vssd1 vccd1 vccd1 _13042_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_68_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11149_ _11181_/A _11149_/B vssd1 vssd1 vccd1 vccd1 _11149_/X sky130_fd_sc_hd__or2_1
XFILLER_1_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11485__A1 _10009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12682__A0 _12681_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09043__A _09999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13226__A2 _13216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08360_ _08360_/A _08360_/B vssd1 vssd1 vccd1 vccd1 _08362_/A sky130_fd_sc_hd__nor2_1
XFILLER_108_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07311_ _07373_/A vssd1 vssd1 vccd1 vccd1 _07311_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08291_ _08573_/A _08547_/A _08291_/C _09233_/C vssd1 vssd1 vccd1 vccd1 _08292_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__08653__A2 _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07242_ _07242_/A vssd1 vssd1 vccd1 vccd1 _14266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07173_ _14101_/Q _07167_/X _07168_/X vssd1 vssd1 vccd1 vccd1 _07173_/X sky130_fd_sc_hd__a21o_2
XFILLER_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07613__A0 _14077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11467__B _11533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09218__A _09491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09814_ _10036_/B _10123_/A vssd1 vssd1 vccd1 vccd1 _09913_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07961__A _09818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09745_ _10541_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09745_/X sky130_fd_sc_hd__or2_1
X_06957_ _14427_/Q _06981_/B _14459_/Q vssd1 vssd1 vccd1 vccd1 _06957_/X sky130_fd_sc_hd__and3b_1
XFILLER_41_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12579__A input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__A1 _11079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _14393_/Q _11659_/A _06858_/Y _14392_/Q vssd1 vssd1 vccd1 vccd1 _06891_/B
+ sky130_fd_sc_hd__a22o_1
X_09676_ _09676_/A _09676_/B _09676_/C vssd1 vssd1 vccd1 vccd1 _09676_/Y sky130_fd_sc_hd__nand3_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _09010_/A _08627_/B vssd1 vssd1 vccd1 vccd1 _08997_/A sky130_fd_sc_hd__xnor2_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08558_ _08555_/X _08558_/B vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__and2b_1
XFILLER_74_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07509_ hold20/X _14183_/Q _07517_/S vssd1 vssd1 vccd1 vccd1 _07510_/A sky130_fd_sc_hd__mux2_1
X_08489_ _09145_/D vssd1 vssd1 vccd1 vccd1 _09084_/C sky130_fd_sc_hd__buf_2
XFILLER_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13203__A _13206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ _10520_/A _10520_/B _10520_/C vssd1 vssd1 vccd1 vccd1 _10522_/B sky130_fd_sc_hd__and3_1
XFILLER_11_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10451_ _10478_/A _10451_/B vssd1 vssd1 vccd1 vccd1 _10455_/C sky130_fd_sc_hd__nand2_1
XFILLER_108_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07604__A0 _14081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ _13171_/A vssd1 vssd1 vccd1 vccd1 _13170_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10382_ _10397_/B _10382_/B vssd1 vssd1 vccd1 vccd1 _10396_/A sky130_fd_sc_hd__xor2_1
XFILLER_109_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12121_ _13812_/Q _12117_/X _12120_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _13812_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07080__A1 _14267_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ _12052_/A vssd1 vssd1 vccd1 vccd1 _13796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08032__A _09443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _11011_/B _11012_/A _11236_/A vssd1 vssd1 vccd1 vccd1 _11008_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12954_ _12954_/A vssd1 vssd1 vccd1 vccd1 _14170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11905_ _13757_/Q _11906_/B vssd1 vssd1 vccd1 vccd1 _11905_/X sky130_fd_sc_hd__and2_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12885_/A vssd1 vssd1 vccd1 vccd1 _12885_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09798__A _09800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _14336_/Q _11833_/X _11834_/X _13795_/Q _11835_/X vssd1 vssd1 vccd1 vccd1
+ _11836_/X sky130_fd_sc_hd__a221o_2
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11767_ input59/X _11767_/B vssd1 vssd1 vccd1 vccd1 _12762_/C sky130_fd_sc_hd__nand2_2
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _13518_/A _13506_/B vssd1 vssd1 vccd1 vccd1 _13507_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_38_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14452_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09310__B _09508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ _11240_/A _10768_/B vssd1 vssd1 vccd1 vccd1 _10719_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11698_ _13755_/Q _13754_/Q _11897_/B vssd1 vssd1 vccd1 vccd1 _11902_/B sky130_fd_sc_hd__or3_1
XANTENNA__08207__A _09762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13437_ input80/X _14378_/Q _13443_/S vssd1 vssd1 vccd1 vccd1 _13438_/B sky130_fd_sc_hd__mux2_1
X_10649_ _10715_/A vssd1 vssd1 vccd1 vccd1 _10650_/A sky130_fd_sc_hd__buf_2
XFILLER_61_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13368_ _12633_/X _14358_/Q _13374_/S vssd1 vssd1 vccd1 vccd1 _13369_/B sky130_fd_sc_hd__mux2_1
X_12319_ _12322_/A vssd1 vssd1 vccd1 vccd1 _12319_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13299_ _13299_/A vssd1 vssd1 vccd1 vccd1 _13299_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10191__B _10191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _14038_/Q _13984_/Q _07859_/Y vssd1 vssd1 vccd1 vccd1 _07861_/B sky130_fd_sc_hd__a21o_1
XFILLER_3_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold12_A hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07791_ _13950_/Q vssd1 vssd1 vccd1 vccd1 _10758_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12655__A0 _12654_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ _09694_/A _09580_/B vssd1 vssd1 vccd1 vccd1 _09581_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11458__A1 _11533_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _09351_/B _09351_/C _09351_/A vssd1 vssd1 vccd1 vccd1 _09462_/C sky130_fd_sc_hd__o21bai_1
Xclkbuf_leaf_77_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14065_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06885__A1 _14395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08412_ _08412_/A vssd1 vssd1 vccd1 vccd1 _08412_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09392_ _09423_/A _09423_/C _09423_/B vssd1 vssd1 vccd1 vccd1 _09392_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08343_ _08343_/A _08343_/B _08343_/C vssd1 vssd1 vccd1 vccd1 _08407_/B sky130_fd_sc_hd__nor3_1
XANTENNA__13023__A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _08274_/A _08274_/B vssd1 vssd1 vccd1 vccd1 _08276_/B sky130_fd_sc_hd__or2_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08117__A _09590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07225_ _07225_/A vssd1 vssd1 vccd1 vccd1 _14271_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_5_0_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12862__A _12906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ _14290_/Q _07155_/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07157_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06860__A _14396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07087_ _07087_/A vssd1 vssd1 vccd1 vccd1 _07087_/X sky130_fd_sc_hd__buf_4
XFILLER_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07989_ _13874_/Q vssd1 vssd1 vccd1 vccd1 _09821_/B sky130_fd_sc_hd__buf_2
XFILLER_86_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ _09729_/A _09729_/B _09729_/C vssd1 vssd1 vccd1 vccd1 _09728_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_90_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09659_ _09263_/X _09415_/Y _09416_/Y _09417_/X vssd1 vssd1 vccd1 vccd1 _10604_/A
+ sky130_fd_sc_hd__a211o_4
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11941__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12668_/X _14050_/Q _12685_/S vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__mux2_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11621_/A vssd1 vssd1 vccd1 vccd1 _13849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14340_ _14400_/CLK _14340_/D vssd1 vssd1 vccd1 vccd1 _14340_/Q sky130_fd_sc_hd__dfxtp_1
X_11552_ _14041_/Q _13953_/Q vssd1 vssd1 vccd1 vccd1 _11650_/A sky130_fd_sc_hd__and2_1
XFILLER_13_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10503_ _10492_/A _10492_/B _10503_/S vssd1 vssd1 vccd1 vccd1 _10505_/A sky130_fd_sc_hd__mux2_1
X_11483_ _11478_/A _11482_/X _11472_/X vssd1 vssd1 vccd1 vccd1 _11483_/X sky130_fd_sc_hd__a21o_1
X_14271_ _14275_/CLK _14271_/D _13131_/Y vssd1 vssd1 vccd1 vccd1 _14271_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_100_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13374__A1 _14360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input71_A io_wbs_datwr[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13222_ _13299_/A vssd1 vssd1 vccd1 vccd1 _13222_/X sky130_fd_sc_hd__clkbuf_2
X_10434_ _10478_/A _10452_/B vssd1 vssd1 vccd1 vccd1 _10453_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13153_ _13153_/A vssd1 vssd1 vccd1 vccd1 _13178_/A sky130_fd_sc_hd__clkbuf_4
X_10365_ _10378_/A _10377_/A vssd1 vssd1 vccd1 vccd1 _10572_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12104_ hold36/A _12095_/X _12103_/X _11931_/X vssd1 vssd1 vccd1 vccd1 _13808_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ input77/X vssd1 vssd1 vccd1 vccd1 _13084_/X sky130_fd_sc_hd__buf_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10297_/A _10297_/B _10297_/C vssd1 vssd1 vccd1 vccd1 _10298_/A sky130_fd_sc_hd__a21oi_1
XANTENNA_output158_A _14313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12035_ _13793_/Q _12020_/X _12021_/X hold40/A vssd1 vssd1 vccd1 vccd1 _12036_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13108__A _13115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13986_ _13986_/CLK _13986_/D _12414_/Y vssd1 vssd1 vccd1 vccd1 _13986_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12937_ hold10/A _12928_/X _12936_/X _12934_/X vssd1 vssd1 vccd1 vccd1 _14161_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13542__S _13542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06867__B2 _14397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12868_ _12911_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__or2_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08863__C _09906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11819_ _13789_/Q _11793_/X _11818_/X vssd1 vssd1 vccd1 vccd1 _11819_/X sky130_fd_sc_hd__a21o_2
XFILLER_18_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12799_ _14115_/Q _12782_/X _12797_/X _12798_/X _12216_/X vssd1 vssd1 vccd1 vccd1
+ _14115_/D sky130_fd_sc_hd__o221a_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11997__S _12000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07292__A1 _14228_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ _14420_/Q _07008_/Y _07009_/X vssd1 vssd1 vccd1 vccd1 _07010_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13365__A1 hold33/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07044__A1 _14304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ _08914_/X _08958_/X _08959_/Y _08960_/Y vssd1 vssd1 vccd1 vccd1 _08961_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11128__B1 _11319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07912_ _07911_/Y _13973_/Q _07912_/S vssd1 vssd1 vccd1 vccd1 _07913_/A sky130_fd_sc_hd__mux2_1
X_08892_ _08892_/A _08892_/B vssd1 vssd1 vccd1 vccd1 _08895_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07843_ _14030_/Q _13976_/Q vssd1 vssd1 vccd1 vccd1 _07843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13018__A _13022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07774_ _11615_/A vssd1 vssd1 vccd1 vccd1 _11585_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09513_ _09511_/X _09513_/B vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__and2b_1
XFILLER_25_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11761__A input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09543_/B _09796_/A _09123_/C _09543_/A vssd1 vssd1 vccd1 vccd1 _09445_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _09291_/B _09291_/C _09291_/A vssd1 vssd1 vccd1 vccd1 _09376_/C sky130_fd_sc_hd__a21bo_1
X_08326_ _08325_/A _08325_/B _08325_/C vssd1 vssd1 vccd1 vccd1 _08326_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__11603__A1 _11602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14447__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08257_ _08257_/A _08257_/B _08257_/C vssd1 vssd1 vccd1 vccd1 _08258_/B sky130_fd_sc_hd__nand3_1
XFILLER_71_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07208_ _07208_/A vssd1 vssd1 vccd1 vccd1 _14276_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08188_ _09685_/A _08121_/B _08120_/A vssd1 vssd1 vccd1 vccd1 _08239_/B sky130_fd_sc_hd__a21oi_1
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13200__B _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07139_ _12205_/A _13838_/Q vssd1 vssd1 vccd1 vccd1 _07185_/A sky130_fd_sc_hd__or2_2
X_10150_ _10636_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _10645_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10081_ _10081_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__xnor2_1
XFILLER_47_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12828__D_N _13200_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08948__C _10206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13840_ _14028_/CLK _13840_/D _12232_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ _13820_/CLK _13771_/D _11964_/Y vssd1 vssd1 vccd1 vccd1 _13771_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10983_ _10652_/A _10934_/X _10920_/X vssd1 vssd1 vccd1 vccd1 _10997_/A sky130_fd_sc_hd__o21ai_1
XFILLER_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12722_ _12722_/A vssd1 vssd1 vccd1 vccd1 _12727_/A sky130_fd_sc_hd__buf_2
XANTENNA__11842__A1 _14339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12653_ _12653_/A vssd1 vssd1 vccd1 vccd1 _14046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11604_ _11604_/A vssd1 vssd1 vccd1 vccd1 _13853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08980__A _08980_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12584_ _12594_/A _12584_/B vssd1 vssd1 vccd1 vccd1 _12585_/A sky130_fd_sc_hd__and2_1
XFILLER_54_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14323_ _14411_/CLK _14323_/D _13193_/Y vssd1 vssd1 vccd1 vccd1 _14323_/Q sky130_fd_sc_hd__dfrtp_4
X_11535_ _11535_/A vssd1 vssd1 vccd1 vccd1 _13859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14254_ _14256_/CLK _14254_/D _13108_/Y vssd1 vssd1 vccd1 vccd1 _14254_/Q sky130_fd_sc_hd__dfstp_1
X_11466_ _11466_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11466_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13205_ _14436_/Q _13201_/X _13204_/X _14388_/Q vssd1 vssd1 vccd1 vccd1 _13205_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07026__A1 _14274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10417_ _10417_/A _10417_/B vssd1 vssd1 vccd1 vccd1 _10564_/C sky130_fd_sc_hd__nand2_1
X_14185_ _14256_/CLK _14185_/D _12972_/Y vssd1 vssd1 vccd1 vccd1 _14185_/Q sky130_fd_sc_hd__dfrtp_1
X_11397_ _13845_/Q _11403_/B vssd1 vssd1 vccd1 vccd1 _11397_/X sky130_fd_sc_hd__or2_1
XFILLER_48_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13136_ _13140_/A vssd1 vssd1 vccd1 vccd1 _13136_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _10341_/A _10341_/B _10347_/X vssd1 vssd1 vccd1 vccd1 _10362_/A sky130_fd_sc_hd__a21o_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13070_/A _13067_/B vssd1 vssd1 vccd1 vccd1 _13068_/A sky130_fd_sc_hd__and2_1
X_10279_ _10279_/A _10279_/B vssd1 vssd1 vccd1 vccd1 _10281_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12018_ _12026_/A _12018_/B vssd1 vssd1 vccd1 vccd1 _12019_/A sky130_fd_sc_hd__and2_1
XFILLER_39_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13969_ _13988_/CLK _13969_/D _12394_/Y vssd1 vssd1 vccd1 vccd1 _13969_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07490_ _14231_/Q _07307_/A _07489_/X _14191_/Q vssd1 vssd1 vccd1 vccd1 _14191_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ _09097_/B _09097_/C _09097_/A vssd1 vssd1 vccd1 vccd1 _09161_/C sky130_fd_sc_hd__a21bo_1
XFILLER_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08111_ _08098_/X _09535_/B _08110_/X vssd1 vssd1 vccd1 vccd1 _08116_/B sky130_fd_sc_hd__a21o_2
X_09091_ _09482_/A _09091_/B vssd1 vssd1 vccd1 vccd1 _09095_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13301__A _13343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08042_ _09491_/A _09508_/C vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__nand2_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10644__B _10644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09993_ _09993_/A _09993_/B vssd1 vssd1 vccd1 vccd1 _09994_/B sky130_fd_sc_hd__and2_1
XFILLER_115_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _08941_/C _08944_/B _08944_/C _08944_/D vssd1 vssd1 vccd1 vccd1 _08944_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_85_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08875_ _08875_/A _08908_/A vssd1 vssd1 vccd1 vccd1 _08875_/X sky130_fd_sc_hd__or2b_1
XFILLER_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08487__D _09941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ _14029_/Q _13975_/Q vssd1 vssd1 vccd1 vccd1 _07900_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12077__B2 _13820_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ _07687_/B _14151_/Q _07757_/S vssd1 vssd1 vccd1 vccd1 _07757_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07688_ _07688_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _07688_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07180__S _07183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09427_ _09427_/A _09427_/B _09427_/C vssd1 vssd1 vccd1 vccd1 _09430_/A sky130_fd_sc_hd__or3_1
XFILLER_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13837__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09358_ _09626_/A _09626_/C vssd1 vssd1 vccd1 vccd1 _09359_/B sky130_fd_sc_hd__and2_1
X_08309_ _13868_/Q vssd1 vssd1 vccd1 vccd1 _09296_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_60_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09289_ _09289_/A _09289_/B vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__xor2_2
X_11320_ _11320_/A _11325_/A vssd1 vssd1 vccd1 vccd1 _11321_/B sky130_fd_sc_hd__or2_1
XFILLER_107_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08305__A _14022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ _13897_/Q vssd1 vssd1 vccd1 vccd1 _11271_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ _10209_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10205_/B sky130_fd_sc_hd__xor2_1
X_11182_ _10975_/A _11166_/X _11180_/X _10918_/A _11181_/X vssd1 vssd1 vccd1 vccd1
+ _11245_/A sky130_fd_sc_hd__o221a_1
XANTENNA__10563__A1 _07924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10133_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10162_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11666__A hold5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13501__A1 _14397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _10064_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__xor2_1
XANTENNA_input34_A io_wbs_adr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_0_io_wbs_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_88_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07192__A0 _14280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13823_ _13826_/CLK _13823_/D vssd1 vssd1 vccd1 vccd1 _13823_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_78_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13754_ _13825_/CLK _13754_/D _11944_/Y vssd1 vssd1 vccd1 vccd1 _13754_/Q sky130_fd_sc_hd__dfrtp_1
X_10966_ _13901_/Q _13902_/Q _13903_/Q _13904_/Q _10670_/B _11186_/S vssd1 vssd1 vccd1
+ vccd1 _10975_/B sky130_fd_sc_hd__mux4_2
X_12705_ _12709_/A vssd1 vssd1 vccd1 vccd1 _12705_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13685_ _13695_/A _13685_/B vssd1 vssd1 vccd1 vccd1 _13686_/A sky130_fd_sc_hd__and2_1
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10897_ _13930_/Q _10896_/Y _10897_/S vssd1 vssd1 vccd1 vccd1 _10898_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12636_ _12636_/A vssd1 vssd1 vccd1 vccd1 _14042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12567_ _13062_/A _12567_/B vssd1 vssd1 vccd1 vccd1 _12611_/S sky130_fd_sc_hd__or2_2
XANTENNA__06942__B _06942_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14306_ _14417_/CLK _14306_/D _13174_/Y vssd1 vssd1 vccd1 vccd1 _14306_/Q sky130_fd_sc_hd__dfrtp_4
X_11518_ _11511_/A _11517_/Y _11464_/X vssd1 vssd1 vccd1 vccd1 _11518_/X sky130_fd_sc_hd__a21o_1
X_12498_ _12817_/A vssd1 vssd1 vccd1 vccd1 _12498_/X sky130_fd_sc_hd__buf_2
XFILLER_8_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_42_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_14237_ _14239_/CLK _14237_/D vssd1 vssd1 vccd1 vccd1 _14237_/Q sky130_fd_sc_hd__dfxtp_1
X_11449_ _11465_/B _11447_/Y _11474_/A vssd1 vssd1 vccd1 vccd1 _11451_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08747__A1 _09234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09944__B1 _10173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14168_ _14283_/CLK _14168_/D _12949_/Y vssd1 vssd1 vccd1 vccd1 _14168_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11576__A _14053_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13121_/A vssd1 vssd1 vccd1 vccd1 _13119_/Y sky130_fd_sc_hd__inv_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _06973_/X _06989_/X hold33/X vssd1 vssd1 vccd1 vccd1 _06991_/S sky130_fd_sc_hd__o21a_1
X_14099_ _14104_/CLK _14099_/D _12749_/Y vssd1 vssd1 vccd1 vccd1 _14099_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07707__C1 _14256_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08660_ _09818_/A vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__07183__A0 _14282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07611_ _14078_/Q input23/X _07615_/S vssd1 vssd1 vccd1 vccd1 _07612_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08591_ _08591_/A _08561_/A vssd1 vssd1 vccd1 vccd1 _08681_/A sky130_fd_sc_hd__or2b_1
XFILLER_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07542_ _14180_/Q _07526_/X _07541_/X _14192_/D vssd1 vssd1 vccd1 vccd1 _14172_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11806__B2 _14235_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07486__A1 _14076_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07473_ _07452_/X _07470_/X _07472_/X _07462_/X _14197_/Q vssd1 vssd1 vccd1 vccd1
+ _14197_/D sky130_fd_sc_hd__a32o_1
XFILLER_90_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08109__B _08791_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09212_ _09212_/A _09212_/B _09212_/C vssd1 vssd1 vccd1 vccd1 _09215_/A sky130_fd_sc_hd__nand3_2
X_09143_ _09140_/X _09141_/Y _09065_/B _09067_/B vssd1 vssd1 vccd1 vccd1 _09180_/B
+ sky130_fd_sc_hd__o211ai_2
X_09074_ _09297_/A _09074_/B vssd1 vssd1 vccd1 vccd1 _09076_/B sky130_fd_sc_hd__nand2_1
XFILLER_108_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08025_ _14015_/Q vssd1 vssd1 vccd1 vccd1 _09297_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12870__A _12913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11486__A _11510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09976_ _10122_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _10285_/B sky130_fd_sc_hd__xnor2_4
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08927_ _08936_/A _09943_/B _08783_/A _08891_/A vssd1 vssd1 vccd1 vccd1 _08928_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_44_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08858_ _08858_/A _08858_/B vssd1 vssd1 vccd1 vccd1 _08859_/B sky130_fd_sc_hd__or2_1
XFILLER_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07174__A0 _14285_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07809_ _07784_/X _11510_/A _07808_/X vssd1 vssd1 vccd1 vccd1 _13987_/D sky130_fd_sc_hd__a21oi_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08789_ _08789_/A _09884_/A vssd1 vssd1 vccd1 vccd1 _08821_/B sky130_fd_sc_hd__and2_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13206__A _13206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10820_ _13940_/Q _10818_/B _10819_/X vssd1 vssd1 vccd1 vccd1 _10835_/B sky130_fd_sc_hd__a21oi_2
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07204__A _07258_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12470__A1 _14031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ _13935_/Q _10803_/B vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__and2_1
XFILLER_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13640__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _13470_/A _13525_/A vssd1 vssd1 vccd1 vccd1 _13497_/A sky130_fd_sc_hd__or2_1
XFILLER_9_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10682_ _10757_/B vssd1 vssd1 vccd1 vccd1 _10730_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14015__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12421_ _12481_/A vssd1 vssd1 vccd1 vccd1 _12460_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12352_ _12353_/A vssd1 vssd1 vccd1 vccd1 _12352_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08977__B2 _08925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08035__A _14016_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ _11312_/A _11303_/B vssd1 vssd1 vccd1 vccd1 _11315_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12283_ _12285_/A vssd1 vssd1 vccd1 vccd1 _12283_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14022_ _14417_/CLK _14022_/D vssd1 vssd1 vccd1 vccd1 _14022_/Q sky130_fd_sc_hd__dfxtp_2
X_11234_ _11285_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11330_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11165_ _13912_/Q _13913_/Q _13914_/Q _13915_/Q _10960_/S _10662_/A vssd1 vssd1 vccd1
+ vccd1 _11165_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10116_ _10116_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_output140_A _11816_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11096_ _11094_/Y _11095_/X _11092_/A _10701_/X vssd1 vssd1 vccd1 vccd1 _13926_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_49_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09154__A1 _08573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09154__B2 _08012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10047_ _10384_/A vssd1 vssd1 vccd1 vccd1 _10053_/A sky130_fd_sc_hd__inv_2
XANTENNA__07165__A0 _14287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06912__B1 _14358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13806_ _14400_/CLK _13806_/D vssd1 vssd1 vccd1 vccd1 _13806_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13116__A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_opt_1_0_io_wbs_clk_A clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12020__A _12059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ _12008_/A _11998_/B vssd1 vssd1 vccd1 vccd1 _11999_/A sky130_fd_sc_hd__and2_1
XFILLER_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13737_ _13737_/A vssd1 vssd1 vccd1 vccd1 _14464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10949_ _11044_/B vssd1 vssd1 vccd1 vccd1 _11134_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12461__A1 _08983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13668_ _13678_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13669_/A sky130_fd_sc_hd__and2_1
XFILLER_31_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12619_ _12635_/A _12619_/B vssd1 vssd1 vccd1 vccd1 _12620_/A sky130_fd_sc_hd__and2_1
X_13599_ _13599_/A vssd1 vssd1 vccd1 vccd1 _14424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__A _11322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10527__B2 _10526_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12921__C1 _12920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08196__A2 _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _10435_/A _09901_/B vssd1 vssd1 vccd1 vccd1 _09830_/X sky130_fd_sc_hd__or2_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _09771_/B _08259_/B _08258_/A vssd1 vssd1 vccd1 vccd1 _09770_/A sky130_fd_sc_hd__o21ai_1
XFILLER_101_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06973_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _09000_/A _09942_/A _08484_/A _08479_/Y vssd1 vssd1 vccd1 vccd1 _08713_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07008__B _14276_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ _09692_/A _09692_/B _09692_/C vssd1 vssd1 vccd1 vccd1 _09692_/Y sky130_fd_sc_hd__nor3_2
XFILLER_67_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08643_ _08643_/A _08643_/B vssd1 vssd1 vccd1 vccd1 _08645_/B sky130_fd_sc_hd__and2_1
XFILLER_26_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ _08547_/A _08824_/C _08547_/D _08573_/A vssd1 vssd1 vccd1 vccd1 _08575_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07525_ _14185_/Q _07534_/B _07519_/X _07524_/X vssd1 vssd1 vccd1 vccd1 _14177_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12452__A1 _14027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10463__A0 _10436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ _07452_/X _07454_/X _07455_/X _07435_/X _14200_/Q vssd1 vssd1 vccd1 vccd1
+ _14200_/D sky130_fd_sc_hd__a32o_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07387_ _14211_/Q _14213_/Q _07387_/S vssd1 vssd1 vccd1 vccd1 _07387_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09126_ _09508_/B _09818_/A _09218_/B _08445_/X vssd1 vssd1 vccd1 vccd1 _09127_/C
+ sky130_fd_sc_hd__a22oi_4
XFILLER_108_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09057_ _09233_/A _09233_/B _09218_/B _09848_/B vssd1 vssd1 vccd1 vccd1 _09060_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_2_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08008_ _13874_/Q vssd1 vssd1 vccd1 vccd1 _09545_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_116_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09959_ _09959_/A _09959_/B vssd1 vssd1 vccd1 vccd1 _09959_/Y sky130_fd_sc_hd__nor2_1
XFILLER_103_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11944__A _11947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12970_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11663__B _11663_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _13822_/Q _11716_/X _11920_/X vssd1 vssd1 vccd1 vccd1 _13762_/D sky130_fd_sc_hd__a21o_1
XFILLER_66_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09414__A _09414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11852_ _14345_/Q _11847_/X _11848_/X _13804_/Q vssd1 vssd1 vccd1 vccd1 _11852_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10279__B _10279_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10803_ _13935_/Q _10803_/B vssd1 vssd1 vccd1 vccd1 _10804_/B sky130_fd_sc_hd__nor2_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13640__A0 _12827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12443__A1 _08683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _13783_/Q _11823_/A _12773_/A _14108_/Q vssd1 vssd1 vccd1 vccd1 _11783_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13522_ _12688_/X _14403_/Q _13522_/S vssd1 vssd1 vccd1 vccd1 _13523_/B sky130_fd_sc_hd__mux2_1
X_10734_ _10936_/A vssd1 vssd1 vccd1 vccd1 _11181_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_28_io_wbs_clk clkbuf_3_3_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13949_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13453_ _13453_/A vssd1 vssd1 vccd1 vccd1 _14382_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665_ _10902_/S vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__buf_4
XFILLER_16_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12404_ _12410_/A vssd1 vssd1 vccd1 vccd1 _12409_/A sky130_fd_sc_hd__buf_2
X_13384_ _13384_/A vssd1 vssd1 vccd1 vccd1 _14362_/D sky130_fd_sc_hd__clkbuf_1
X_10596_ _10596_/A _10596_/B _10596_/C vssd1 vssd1 vccd1 vccd1 _10597_/C sky130_fd_sc_hd__and3_1
XFILLER_86_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12335_ _12335_/A vssd1 vssd1 vccd1 vccd1 _12335_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12266_ _12267_/A vssd1 vssd1 vccd1 vccd1 _12266_/Y sky130_fd_sc_hd__inv_2
X_14005_ _14442_/CLK _14005_/D vssd1 vssd1 vccd1 vccd1 _14005_/Q sky130_fd_sc_hd__dfxtp_1
X_11217_ _11217_/A _11217_/B vssd1 vssd1 vccd1 vccd1 _11297_/B sky130_fd_sc_hd__xnor2_2
X_12197_ _13197_/B vssd1 vssd1 vccd1 vccd1 _13079_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_110_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11148_ _13919_/Q _13920_/Q _13921_/Q _13922_/Q _11169_/S _07798_/A vssd1 vssd1 vccd1
+ vccd1 _11149_/B sky130_fd_sc_hd__mux4_1
XFILLER_62_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11079_ _11079_/A _11079_/B vssd1 vssd1 vccd1 vccd1 _11080_/B sky130_fd_sc_hd__or2_1
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07689__A1 _14133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12682__A1 _14053_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_io_wbs_clk clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14442_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13631__A0 input89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07310_ _07462_/A vssd1 vssd1 vccd1 vccd1 _07373_/A sky130_fd_sc_hd__buf_2
X_08290_ _08126_/A _09445_/B _09793_/A _08128_/A vssd1 vssd1 vccd1 vccd1 _08292_/A
+ sky130_fd_sc_hd__a22oi_1
X_07241_ _14266_/Q _07239_/X _07253_/S vssd1 vssd1 vccd1 vccd1 _07242_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07172_ _07172_/A vssd1 vssd1 vccd1 vccd1 _14286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13698__A0 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08403__A _08403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09218__B _09218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09813_ _10045_/A vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__buf_2
XFILLER_28_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09744_ _10540_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09745_/B sky130_fd_sc_hd__or2_2
XFILLER_86_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06956_ _14283_/Q _06929_/X _06955_/X _14379_/Q vssd1 vssd1 vccd1 vccd1 _06956_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09234__A _09234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09675_ _09675_/A vssd1 vssd1 vccd1 vccd1 _09675_/Y sky130_fd_sc_hd__inv_2
X_06887_ _14392_/Q _06858_/Y _11679_/A _14391_/Q vssd1 vssd1 vccd1 vccd1 _06891_/A
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08626_ _08626_/A _08626_/B vssd1 vssd1 vccd1 vccd1 _08627_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11881__C1 _11874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _08555_/B _09906_/A _08863_/D _09001_/A vssd1 vssd1 vccd1 vccd1 _08558_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07508_ _07521_/D vssd1 vssd1 vccd1 vccd1 _07517_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_11_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08488_ _09865_/B vssd1 vssd1 vccd1 vccd1 _09085_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07439_ _07458_/A _07439_/B vssd1 vssd1 vccd1 vccd1 _07439_/X sky130_fd_sc_hd__or2_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10450_ _10450_/A _10450_/B vssd1 vssd1 vccd1 vccd1 _10457_/A sky130_fd_sc_hd__or2_1
XFILLER_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09109_ _09106_/Y _09107_/X _09025_/C _09025_/Y vssd1 vssd1 vccd1 vccd1 _09110_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__07065__C1 _14356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _10381_/A _10358_/A vssd1 vssd1 vccd1 vccd1 _10391_/C sky130_fd_sc_hd__or2b_1
X_12120_ _12938_/A _12130_/B vssd1 vssd1 vccd1 vccd1 _12120_/X sky130_fd_sc_hd__or2_1
XANTENNA__10562__B _10562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12051_ _12065_/A _12051_/B vssd1 vssd1 vccd1 vccd1 _12052_/A sky130_fd_sc_hd__and2_1
XFILLER_85_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11002_ _11073_/B _11002_/B vssd1 vssd1 vccd1 vccd1 _11102_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07907__A2 _07921_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12953_ _14170_/Q _13111_/B _13358_/B vssd1 vssd1 vccd1 vccd1 _12954_/A sky130_fd_sc_hd__and3b_1
X_11904_ hold17/X _11872_/X _11903_/Y _11874_/X vssd1 vssd1 vccd1 vccd1 _13756_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06879__C1 _14365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12884_ _14142_/Q _12872_/X _12883_/X _12879_/X vssd1 vssd1 vccd1 vccd1 _14142_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08983__A _08983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _14001_/Q _11797_/A _11830_/X _14120_/Q vssd1 vssd1 vccd1 vccd1 _11835_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11766_ _12951_/A _11766_/B vssd1 vssd1 vccd1 vccd1 _11768_/A sky130_fd_sc_hd__nand2_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _12668_/X _14398_/Q _13511_/S vssd1 vssd1 vccd1 vccd1 _13506_/B sky130_fd_sc_hd__mux2_1
X_10717_ _10727_/B _10727_/C vssd1 vssd1 vccd1 vccd1 _10768_/B sky130_fd_sc_hd__nand2_1
X_11697_ _13753_/Q _11893_/B vssd1 vssd1 vccd1 vccd1 _11897_/B sky130_fd_sc_hd__or2_1
XANTENNA__08207__B _09999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13436_ _13436_/A vssd1 vssd1 vccd1 vccd1 _14377_/D sky130_fd_sc_hd__clkbuf_1
X_10648_ _10648_/A vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__buf_2
XFILLER_42_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12952__B _12952_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13367_ _13367_/A vssd1 vssd1 vccd1 vccd1 _14357_/D sky130_fd_sc_hd__clkbuf_1
X_10579_ _10644_/A _10572_/Y _10578_/X vssd1 vssd1 vccd1 vccd1 _10579_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09319__A _09319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12318_ _12322_/A vssd1 vssd1 vccd1 vccd1 _12318_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _14373_/Q _13215_/A _13294_/X _14453_/Q vssd1 vssd1 vccd1 vccd1 _13298_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08223__A _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12249_ _12251_/A vssd1 vssd1 vccd1 vccd1 _12249_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07790_ _10875_/S vssd1 vssd1 vccd1 vccd1 _11119_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09460_ _09459_/B _09459_/C _08098_/X vssd1 vssd1 vccd1 vccd1 _09462_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__08893__A _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ _10524_/A _10523_/B vssd1 vssd1 vccd1 vccd1 _08412_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09391_ _09391_/A vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08342_ _08343_/A _08343_/B _08343_/C vssd1 vssd1 vccd1 vccd1 _09751_/C sky130_fd_sc_hd__o21a_1
X_08273_ _08273_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _08276_/A sky130_fd_sc_hd__xnor2_1
X_07224_ _14271_/Q _07222_/X _07236_/S vssd1 vssd1 vccd1 vccd1 _07225_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11759__A input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _14106_/Q _07140_/X _07143_/X vssd1 vssd1 vccd1 vccd1 _07155_/X sky130_fd_sc_hd__a21o_4
XANTENNA__07598__A0 _14084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14473__185 vssd1 vssd1 vccd1 vccd1 _14473__185/HI io_oeb[5] sky130_fd_sc_hd__conb_1
XFILLER_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07086_ _14442_/Q _14266_/Q vssd1 vssd1 vccd1 vccd1 _07086_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08133__A _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07972__A _13873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07988_ _09434_/A vssd1 vssd1 vccd1 vccd1 _08571_/A sky130_fd_sc_hd__buf_2
XANTENNA__07183__S _07183_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09727_ _09727_/A _09727_/B _09727_/C vssd1 vssd1 vccd1 vccd1 _09727_/Y sky130_fd_sc_hd__nor3_2
X_06939_ _14461_/Q _14285_/Q vssd1 vssd1 vccd1 vccd1 _06939_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_3_7_0_io_wbs_clk clkbuf_3_7_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_io_wbs_clk/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_55_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09658_ _09657_/X _09273_/A _09267_/B vssd1 vssd1 vccd1 vccd1 _10613_/B sky130_fd_sc_hd__a21oi_4
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _08681_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08610_/B sky130_fd_sc_hd__xnor2_1
XFILLER_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09589_ _09549_/A _09549_/B _09588_/X vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__a21o_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13214__A _13328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ hold9/A _11619_/Y _11632_/S vssd1 vssd1 vccd1 vccd1 _11621_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ _14040_/Q _13952_/Q vssd1 vssd1 vccd1 vccd1 _11651_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10502_ _10503_/S _10497_/B _10496_/A vssd1 vssd1 vccd1 vccd1 _10506_/A sky130_fd_sc_hd__a21oi_1
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14270_ _14275_/CLK _14270_/D _13130_/Y vssd1 vssd1 vccd1 vccd1 _14270_/Q sky130_fd_sc_hd__dfrtp_4
X_11482_ _11482_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11482_/X sky130_fd_sc_hd__or2_1
XFILLER_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13221_ _13341_/A vssd1 vssd1 vccd1 vccd1 _13299_/A sky130_fd_sc_hd__clkbuf_2
X_10433_ _10449_/B _10433_/B vssd1 vssd1 vccd1 vccd1 _10452_/B sky130_fd_sc_hd__and2_1
XFILLER_87_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input64_A io_wbs_adr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ _13152_/A vssd1 vssd1 vccd1 vccd1 _13152_/Y sky130_fd_sc_hd__inv_2
X_10364_ _10364_/A _10364_/B _10364_/C vssd1 vssd1 vccd1 vccd1 _10377_/A sky130_fd_sc_hd__nand3_1
XFILLER_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_47_io_wbs_clk_A clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_3_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12103_ _12926_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12103_/X sky130_fd_sc_hd__or2_1
XFILLER_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13083_ _13083_/A vssd1 vssd1 vccd1 vccd1 _14246_/D sky130_fd_sc_hd__clkbuf_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10295_ _10367_/A vssd1 vssd1 vccd1 vccd1 _10407_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08978__A _08978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ _12034_/A vssd1 vssd1 vccd1 vccd1 _13792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13985_ _13986_/CLK _13985_/D _12413_/Y vssd1 vssd1 vccd1 vccd1 _13985_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12936_ _12936_/A _12940_/B vssd1 vssd1 vccd1 vccd1 _12936_/X sky130_fd_sc_hd__or2_1
XANTENNA__07106__B _07134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _14135_/Q _12857_/X _12864_/X _12866_/X vssd1 vssd1 vccd1 vccd1 _14135_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11818_ _14330_/Q _11833_/A _11770_/X _14238_/Q _11817_/X vssd1 vssd1 vccd1 vccd1
+ _11818_/X sky130_fd_sc_hd__a221o_1
XFILLER_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12798_ _14140_/Q _12776_/A _12791_/X vssd1 vssd1 vccd1 vccd1 _12798_/X sky130_fd_sc_hd__a21o_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11749_ _14255_/Q vssd1 vssd1 vccd1 vccd1 _11749_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13419_ input74/X _14373_/Q _13425_/S vssd1 vssd1 vccd1 vccd1 _13420_/B sky130_fd_sc_hd__mux2_1
X_14399_ _14400_/CLK _14399_/D vssd1 vssd1 vccd1 vccd1 _14399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08960_ _08960_/A _08960_/B vssd1 vssd1 vccd1 vccd1 _08960_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11128__A1 _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08888__A _08978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07911_ _07911_/A _07911_/B vssd1 vssd1 vccd1 vccd1 _07911_/Y sky130_fd_sc_hd__nor2_1
X_08891_ _08891_/A _08936_/A _09942_/A _08925_/C vssd1 vssd1 vccd1 vccd1 _08892_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07842_ _07900_/B _07901_/B _07900_/A vssd1 vssd1 vccd1 vccd1 _07897_/A sky130_fd_sc_hd__o21ba_1
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12203__A _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07773_ _11655_/B vssd1 vssd1 vccd1 vccd1 _11615_/A sky130_fd_sc_hd__inv_2
X_09512_ _09511_/B _09511_/C _09511_/A vssd1 vssd1 vccd1 vccd1 _09513_/B sky130_fd_sc_hd__a21o_1
XFILLER_65_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07504__A0 hold29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11761__B _11774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ _09443_/A _09493_/B _09493_/D _09818_/A vssd1 vssd1 vccd1 vccd1 _09489_/A
+ sky130_fd_sc_hd__nand4_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09374_ _09373_/A _09373_/C _09373_/B vssd1 vssd1 vccd1 vccd1 _09376_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08325_ _08325_/A _08325_/B _08325_/C vssd1 vssd1 vccd1 vccd1 _08325_/X sky130_fd_sc_hd__and3_1
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08256_ _08257_/B _08257_/C _08257_/A vssd1 vssd1 vccd1 vccd1 _08258_/A sky130_fd_sc_hd__a21o_1
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07207_ _14276_/Q _07205_/X _07219_/S vssd1 vssd1 vccd1 vccd1 _07208_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13356__A2 _13265_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ _09694_/A vssd1 vssd1 vccd1 vccd1 _09673_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10393__A _10393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07138_ _13839_/Q vssd1 vssd1 vccd1 vccd1 _12205_/A sky130_fd_sc_hd__clkbuf_2
X_07069_ _07065_/X _14301_/Q _07069_/S vssd1 vssd1 vccd1 vccd1 _07070_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10080_ _10080_/A vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__buf_2
XANTENNA__13766__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12113__A _13609_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13643__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13770_ _13825_/CLK _13770_/D _11963_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08299__A1 _08113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ _10651_/A _10965_/X _10920_/X vssd1 vssd1 vccd1 vccd1 _11000_/A sky130_fd_sc_hd__o21ai_2
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12721_ _12721_/A vssd1 vssd1 vccd1 vccd1 _12721_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12652_ _12656_/A _12652_/B vssd1 vssd1 vccd1 vccd1 _12653_/A sky130_fd_sc_hd__and2_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11603_ _13853_/Q _11602_/Y _11611_/S vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12583_ _12913_/A _14028_/Q _12583_/S vssd1 vssd1 vccd1 vccd1 _12584_/B sky130_fd_sc_hd__mux2_1
XFILLER_15_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08980__B _08980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14322_ _14322_/CLK _14322_/D _13192_/Y vssd1 vssd1 vccd1 vccd1 _14322_/Q sky130_fd_sc_hd__dfrtp_4
X_11534_ _10206_/A _11533_/X _11534_/S vssd1 vssd1 vccd1 vccd1 _11535_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14253_ _14259_/CLK _14253_/D vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_2
XFILLER_99_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11465_ _11474_/A _11465_/B vssd1 vssd1 vccd1 vccd1 _11465_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12555__A0 _12936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13204_ _13245_/A vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__clkbuf_2
X_10416_ _10416_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10417_/B sky130_fd_sc_hd__or2_1
X_14184_ _14256_/CLK _14184_/D _12971_/Y vssd1 vssd1 vccd1 vccd1 _14184_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_output170_A _14295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11396_ _11396_/A vssd1 vssd1 vccd1 vccd1 _11396_/X sky130_fd_sc_hd__clkbuf_2
X_13135_ _13147_/A vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__buf_2
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10347_ _10347_/A _10347_/B vssd1 vssd1 vccd1 vccd1 _10347_/X sky130_fd_sc_hd__and2_1
XFILLER_97_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _12633_/X hold23/A _13076_/S vssd1 vssd1 vccd1 vccd1 _13067_/B sky130_fd_sc_hd__mux2_1
X_10278_ _10278_/A _10278_/B vssd1 vssd1 vccd1 vccd1 _10288_/A sky130_fd_sc_hd__xor2_1
X_12017_ _13788_/Q _12000_/X _12003_/X _13828_/Q vssd1 vssd1 vccd1 vccd1 _12018_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13968_ _13988_/CLK _13968_/D _12393_/Y vssd1 vssd1 vccd1 vccd1 _13968_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12919_ _12919_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _12919_/X sky130_fd_sc_hd__or2_1
X_13899_ _13905_/CLK _13899_/D _12307_/Y vssd1 vssd1 vccd1 vccd1 _13899_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08110_ _08435_/A _09535_/A vssd1 vssd1 vccd1 vccd1 _08110_/X sky130_fd_sc_hd__and2_1
XFILLER_119_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09090_ _09090_/A _09090_/B _09090_/C vssd1 vssd1 vccd1 vccd1 _09097_/A sky130_fd_sc_hd__nand3_1
XFILLER_30_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08041_ _14015_/Q vssd1 vssd1 vccd1 vccd1 _09491_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11349__B2 _10669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10644__C _10644_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09992_ _09993_/A _09993_/B vssd1 vssd1 vccd1 vccd1 _09994_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08943_ _08937_/B _08937_/C _10171_/A _08946_/A vssd1 vssd1 vccd1 vccd1 _08944_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13029__A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ _08908_/A _08875_/A vssd1 vssd1 vccd1 vccd1 _08880_/B sky130_fd_sc_hd__xor2_1
XFILLER_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07825_ _14030_/Q _13976_/Q vssd1 vssd1 vccd1 vccd1 _07896_/A sky130_fd_sc_hd__nor2_1
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12868__A _12911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07756_ _14063_/Q _07720_/X _07754_/X _07755_/Y vssd1 vssd1 vccd1 vccd1 _14063_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_72_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12077__A2 _12000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14414__CLK _14449_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07687_ _07687_/A _07687_/B vssd1 vssd1 vccd1 vccd1 _07687_/Y sky130_fd_sc_hd__nand2_1
X_09426_ _09472_/B _09844_/B _09807_/A _09361_/A vssd1 vssd1 vccd1 vccd1 _09427_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09357_ _09455_/A _09356_/C _09537_/A vssd1 vssd1 vccd1 vccd1 _09626_/C sky130_fd_sc_hd__a21o_1
XANTENNA__07332__B_N _07323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _09424_/A _09361_/B _09803_/B _09473_/B vssd1 vssd1 vccd1 vccd1 _08313_/A
+ sky130_fd_sc_hd__nand4_2
X_09288_ _08794_/B _09286_/X _09287_/X vssd1 vssd1 vccd1 vccd1 _09289_/B sky130_fd_sc_hd__a21bo_1
X_08239_ _09777_/B _08239_/B vssd1 vssd1 vccd1 vccd1 _08239_/X sky130_fd_sc_hd__or2_1
XFILLER_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12537__A0 _12922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _11273_/A _11273_/B vssd1 vssd1 vccd1 vccd1 _11341_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10201_ _10209_/A _10202_/B vssd1 vssd1 vccd1 vccd1 _10204_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11947__A _11947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07413__C1 _07521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ _11181_/A _11181_/B vssd1 vssd1 vccd1 vccd1 _11181_/X sky130_fd_sc_hd__or2_1
XFILLER_106_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10132_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10136_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11666__B _14259_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10063_ _10112_/B _10063_/B vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__xnor2_1
XFILLER_87_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input27_A dout1[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13822_ _13825_/CLK _13822_/D vssd1 vssd1 vccd1 vccd1 _13822_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12068__A2 _12059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14094__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__A _09152_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13753_ _13826_/CLK _13753_/D _11943_/Y vssd1 vssd1 vccd1 vccd1 _13753_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10965_ _10914_/X _10964_/X _11152_/S vssd1 vssd1 vccd1 vccd1 _10965_/X sky130_fd_sc_hd__mux2_2
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ _12722_/A vssd1 vssd1 vccd1 vccd1 _12709_/A sky130_fd_sc_hd__buf_2
XFILLER_91_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ _12681_/X _14449_/Q _13687_/S vssd1 vssd1 vccd1 vccd1 _13685_/B sky130_fd_sc_hd__mux2_1
X_10896_ _10906_/A _10889_/C _10894_/X _10895_/Y vssd1 vssd1 vccd1 vccd1 _10896_/Y
+ sky130_fd_sc_hd__o31ai_1
X_12635_ _12635_/A _12635_/B vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__and2_1
XFILLER_19_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12566_ _12942_/A _12520_/S _12565_/Y vssd1 vssd1 vccd1 vccd1 _14023_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07400__A _07464_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ _11517_/A _11517_/B vssd1 vssd1 vccd1 vccd1 _11517_/Y sky130_fd_sc_hd__nand2_1
X_14305_ _14417_/CLK _14305_/D _13173_/Y vssd1 vssd1 vccd1 vccd1 _14305_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _14038_/Q _12485_/X _12496_/X _12473_/A vssd1 vssd1 vccd1 vccd1 _12497_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14236_ _14239_/CLK _14236_/D vssd1 vssd1 vccd1 vccd1 _14236_/Q sky130_fd_sc_hd__dfxtp_2
X_11448_ _11467_/A vssd1 vssd1 vccd1 vccd1 _11474_/A sky130_fd_sc_hd__clkinv_2
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08747__A2 _09887_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14167_ _14283_/CLK _14167_/D _12948_/Y vssd1 vssd1 vccd1 vccd1 _14167_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11379_ _11392_/A vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__clkbuf_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07546__S _07548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13118_ _13121_/A vssd1 vssd1 vccd1 vccd1 _13118_/Y sky130_fd_sc_hd__inv_2
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14102_/CLK _14098_/D _12748_/Y vssd1 vssd1 vccd1 vccd1 _14098_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ hold21/A _13036_/S _13042_/Y hold20/A _13032_/A vssd1 vssd1 vccd1 vccd1 _13049_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07610_ _07610_/A vssd1 vssd1 vccd1 vccd1 _14079_/D sky130_fd_sc_hd__clkbuf_1
X_08590_ _08590_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _08682_/A sky130_fd_sc_hd__and2_1
XFILLER_54_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13256__B2 _14396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07541_ _07541_/A _07541_/B _07541_/C vssd1 vssd1 vccd1 vccd1 _07541_/X sky130_fd_sc_hd__or3_1
XFILLER_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09997__A _10393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07486__A2 _11746_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ _14080_/Q _07459_/X _07460_/X _13880_/Q _07471_/X vssd1 vssd1 vccd1 vccd1
+ _07472_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09211_ _09205_/A _09205_/B _09205_/C vssd1 vssd1 vccd1 vccd1 _09212_/C sky130_fd_sc_hd__a21o_1
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08109__C _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09142_ _09065_/B _09067_/B _09140_/X _09141_/Y vssd1 vssd1 vccd1 vccd1 _09194_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07310__A _07462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ _09543_/A _09217_/B _09843_/A _09881_/B vssd1 vssd1 vccd1 vccd1 _09164_/A
+ sky130_fd_sc_hd__and4_2
XANTENNA__06884__A1_N _14395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08024_ _08024_/A _08024_/B _08024_/C vssd1 vssd1 vccd1 vccd1 _08325_/B sky130_fd_sc_hd__nand3_1
XFILLER_116_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11767__A input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09975_ _10123_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__xor2_2
X_08926_ _09055_/A _08944_/D vssd1 vssd1 vccd1 vccd1 _08939_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08857_ _08962_/A _08962_/B _08856_/X vssd1 vssd1 vccd1 vccd1 _08857_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07174__A1 _07173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07808_ _11119_/A _10705_/B _07807_/Y _07779_/A vssd1 vssd1 vccd1 vccd1 _07808_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08788_ _08787_/A _08787_/C _08787_/B vssd1 vssd1 vccd1 vccd1 _08799_/C sky130_fd_sc_hd__o21ai_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13206__B _13359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07739_ _14068_/Q _07720_/X _07737_/X _07738_/Y vssd1 vssd1 vccd1 vccd1 _14068_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10750_ _11236_/A _10746_/A _10750_/S vssd1 vssd1 vccd1 vccd1 _10803_/B sky130_fd_sc_hd__mux2_1
XFILLER_77_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09871__B1 _10092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13892_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_09409_ _09335_/A _09335_/B _09408_/X vssd1 vssd1 vccd1 vccd1 _09411_/B sky130_fd_sc_hd__o21ai_2
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ _11155_/S vssd1 vssd1 vccd1 vccd1 _10757_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _12440_/A _13209_/A _13194_/C vssd1 vssd1 vccd1 vccd1 _12481_/A sky130_fd_sc_hd__and3_1
XANTENNA__10565__B _10565_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ _12353_/A vssd1 vssd1 vccd1 vccd1 _12351_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08977__A2 _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11302_ _11302_/A _11302_/B vssd1 vssd1 vccd1 vccd1 _11303_/B sky130_fd_sc_hd__or2_1
XFILLER_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _12285_/A vssd1 vssd1 vccd1 vccd1 _12282_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14021_ _14304_/CLK _14021_/D vssd1 vssd1 vccd1 vccd1 _14021_/Q sky130_fd_sc_hd__dfxtp_2
X_11233_ _11233_/A _11233_/B vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__xor2_4
XFILLER_20_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11733__B2 _13826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ _11181_/B _11163_/X _11164_/S vssd1 vssd1 vccd1 vccd1 _11164_/X sky130_fd_sc_hd__mux2_2
XFILLER_96_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10115_ _10245_/B _10115_/B vssd1 vssd1 vccd1 vccd1 _10116_/B sky130_fd_sc_hd__xnor2_2
Xclkbuf_1_0_1_io_wbs_clk clkbuf_1_0_1_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_io_wbs_clk/A
+ sky130_fd_sc_hd__clkbuf_2
X_11095_ _11083_/A _11084_/X _11093_/Y _11125_/A vssd1 vssd1 vccd1 vccd1 _11095_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_1_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10046_ _10271_/A _10044_/X _10045_/X vssd1 vssd1 vccd1 vccd1 _10384_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07165__A1 _07164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_io_wbs_clk clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14450_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12301__A _12304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06912__A1 _06894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13805_ _14348_/CLK _13805_/D vssd1 vssd1 vccd1 vccd1 _13805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11997_ _11991_/X _13783_/Q _12000_/A vssd1 vssd1 vccd1 vccd1 _11998_/B sky130_fd_sc_hd__mux2_1
XFILLER_95_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10948_ _10758_/A _10943_/X _10932_/X _10743_/A _10947_/X vssd1 vssd1 vccd1 vccd1
+ _11044_/B sky130_fd_sc_hd__a221oi_2
X_13736_ _13745_/A _13736_/B vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__and2_1
XFILLER_44_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ _12660_/X _14444_/Q _13670_/S vssd1 vssd1 vccd1 vccd1 _13668_/B sky130_fd_sc_hd__mux2_1
X_10879_ _10798_/Y _10879_/B _10879_/C vssd1 vssd1 vccd1 vccd1 _10879_/X sky130_fd_sc_hd__and3b_1
XFILLER_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12618_ _12940_/A _14038_/Q _12621_/S vssd1 vssd1 vccd1 vccd1 _12619_/B sky130_fd_sc_hd__mux2_1
X_13598_ _13607_/A _13598_/B vssd1 vssd1 vccd1 vccd1 _13599_/A sky130_fd_sc_hd__and2_1
XFILLER_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12549_ _12549_/A vssd1 vssd1 vccd1 vccd1 _14018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14219_ _14284_/CLK _14219_/D _13015_/Y vssd1 vssd1 vccd1 vccd1 _14219_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10527__A2 _07924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _09777_/A _08272_/B _08271_/A vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__o21a_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _14281_/Q _06968_/X _06971_/X _14377_/Q vssd1 vssd1 vccd1 vccd1 _06972_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08896__A _08896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13827__CLK _14335_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _09905_/A vssd1 vssd1 vccd1 vccd1 _09942_/A sky130_fd_sc_hd__buf_4
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11488__B1 _10686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09691_ _09687_/Y _09688_/X _09607_/B _09675_/Y vssd1 vssd1 vccd1 vccd1 _09692_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07156__A1 _07155_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08642_ _08997_/A _08997_/B vssd1 vssd1 vccd1 vccd1 _08645_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13307__A _13328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12211__A _12211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08573_ _08573_/A _08573_/B _08824_/C _09084_/D vssd1 vssd1 vccd1 vccd1 _08573_/X
+ sky130_fd_sc_hd__and4_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09223__C _09223_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13741__S _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07524_ _14177_/Q _07520_/B _07528_/A _07523_/X vssd1 vssd1 vccd1 vccd1 _07524_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07024__B _14274_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07455_ _14083_/Q _07432_/X _07433_/X _13883_/Q _07444_/X vssd1 vssd1 vccd1 vccd1
+ _07455_/X sky130_fd_sc_hd__a221o_1
XFILLER_74_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07959__B _08251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07386_ _14095_/Q _07363_/X vssd1 vssd1 vccd1 vccd1 _07386_/X sky130_fd_sc_hd__or2b_1
XFILLER_109_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09125_ _09349_/A _09553_/D vssd1 vssd1 vccd1 vccd1 _09127_/B sky130_fd_sc_hd__nand2_2
XFILLER_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12881__A _12924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09056_ _09056_/A _09056_/B vssd1 vssd1 vccd1 vccd1 _09065_/A sky130_fd_sc_hd__xnor2_1
XFILLER_117_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08007_ _08623_/B vssd1 vssd1 vccd1 vccd1 _08126_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09958_ _10346_/A _09997_/B _09957_/X vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__a21boi_2
X_08909_ _08915_/A _08915_/B vssd1 vssd1 vccd1 vccd1 _08916_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11479__B1 _10686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A1 _13951_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _10050_/B _10059_/A vssd1 vssd1 vccd1 vccd1 _10129_/B sky130_fd_sc_hd__nor2_2
XANTENNA__10274__C_N _10272_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13217__A _13637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11920_ _11920_/A _13762_/Q _11920_/C vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__and3_1
XANTENNA__09414__B _09660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _14344_/Q _11847_/X _11848_/X _13803_/Q vssd1 vssd1 vccd1 vccd1 _11851_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11960__A _11971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10802_ _10873_/B _10873_/C _10873_/A vssd1 vssd1 vccd1 vccd1 _10874_/A sky130_fd_sc_hd__o21a_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _12193_/A _12762_/B _12762_/C vssd1 vssd1 vccd1 vccd1 _12773_/A sky130_fd_sc_hd__nor3_4
XFILLER_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ _10951_/A _11158_/S vssd1 vssd1 vccd1 vccd1 _10936_/A sky130_fd_sc_hd__or2b_2
X_13521_ _13592_/A vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__buf_2
X_13452_ _13461_/A _13452_/B vssd1 vssd1 vccd1 vccd1 _13453_/A sky130_fd_sc_hd__and2_1
XANTENNA_input94_A io_wbs_datwr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10664_ _11452_/A _10664_/B vssd1 vssd1 vccd1 vccd1 _10902_/S sky130_fd_sc_hd__nor2_2
XANTENNA__08046__A _09482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12403_ _12403_/A vssd1 vssd1 vccd1 vccd1 _12403_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13383_ _13392_/A _13383_/B vssd1 vssd1 vccd1 vccd1 _13384_/A sky130_fd_sc_hd__and2_1
X_10595_ _13959_/Q _10545_/X _10594_/X vssd1 vssd1 vccd1 vccd1 _13959_/D sky130_fd_sc_hd__o21a_1
XFILLER_12_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12334_ _12335_/A vssd1 vssd1 vccd1 vccd1 _12334_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12265_ _12267_/A vssd1 vssd1 vccd1 vccd1 _12265_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14004_ _14442_/CLK _14004_/D vssd1 vssd1 vccd1 vccd1 _14004_/Q sky130_fd_sc_hd__dfxtp_1
X_11216_ _11216_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11217_/B sky130_fd_sc_hd__nand2_1
X_12196_ input33/X input44/X _12196_/C vssd1 vssd1 vccd1 vccd1 _13197_/B sky130_fd_sc_hd__or3_4
XFILLER_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11147_ _10713_/A _11146_/X _11140_/X vssd1 vssd1 vccd1 vccd1 _11147_/X sky130_fd_sc_hd__o21a_1
XFILLER_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11078_ _11102_/B _11105_/B _11102_/A vssd1 vssd1 vccd1 vccd1 _11099_/C sky130_fd_sc_hd__o21ai_1
XFILLER_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10029_ _10244_/A _10244_/B _10028_/X vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__a21oi_2
XFILLER_36_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06897__B1 _14365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_54_io_wbs_clk_A clkbuf_3_6_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_60_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13719_ _13729_/A _13719_/B vssd1 vssd1 vccd1 vccd1 _13720_/A sky130_fd_sc_hd__and2_1
XFILLER_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07240_ _07240_/A vssd1 vssd1 vccd1 vccd1 _07253_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07171_ _14286_/Q _07169_/X _07183_/S vssd1 vssd1 vccd1 vccd1 _07172_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08574__B1 _08547_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ _09842_/A _09875_/B _09811_/X vssd1 vssd1 vccd1 vccd1 _10045_/A sky130_fd_sc_hd__a21oi_4
XFILLER_119_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06955_ _14427_/Q _06954_/Y _06931_/X vssd1 vssd1 vccd1 vccd1 _06955_/X sky130_fd_sc_hd__a21o_1
X_09743_ _09739_/C _09737_/X _09704_/X _09706_/Y vssd1 vssd1 vccd1 vccd1 _09744_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_100_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07129__A1 _14293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09674_ _09777_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09674_/X sky130_fd_sc_hd__or2_1
X_06886_ _13778_/Q vssd1 vssd1 vccd1 vccd1 _11679_/A sky130_fd_sc_hd__inv_2
XFILLER_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _08623_/X _08625_/B vssd1 vssd1 vccd1 vccd1 _08626_/B sky130_fd_sc_hd__and2b_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__A _12919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08556_ _08748_/B vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__buf_4
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07507_ _07507_/A vssd1 vssd1 vccd1 vccd1 _14184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08487_ _09443_/A _09493_/B _09199_/D _09941_/A vssd1 vssd1 vccd1 vccd1 _08560_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07438_ _14202_/Q _14204_/Q _07442_/S vssd1 vssd1 vccd1 vccd1 _07439_/B sky130_fd_sc_hd__mux2_1
XFILLER_74_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07369_ _14098_/Q _07363_/X vssd1 vssd1 vccd1 vccd1 _07369_/X sky130_fd_sc_hd__or2b_1
X_09108_ _09025_/C _09025_/Y _09106_/Y _09107_/X vssd1 vssd1 vccd1 vccd1 _09118_/A
+ sky130_fd_sc_hd__a211o_1
X_10380_ _10380_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__or2_1
X_09039_ _08780_/X _08963_/X _10631_/A _09037_/X _09038_/Y vssd1 vssd1 vccd1 vccd1
+ _10644_/B sky130_fd_sc_hd__a2111o_4
XFILLER_108_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11020__A _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ _13796_/Q _12038_/X _12039_/X _13812_/Q vssd1 vssd1 vccd1 vccd1 _12051_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11001_ _13922_/Q vssd1 vssd1 vccd1 vccd1 _11002_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__08032__C _08097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09425__A _09425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08868__A1 _08896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ _13197_/A _12952_/B vssd1 vssd1 vccd1 vccd1 _13358_/B sky130_fd_sc_hd__nor2_4
XANTENNA__08868__B2 _08983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14224_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11903_ _11906_/B _11903_/B vssd1 vssd1 vccd1 vccd1 _11903_/Y sky130_fd_sc_hd__nand2_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12926_/A _12883_/B vssd1 vssd1 vccd1 vccd1 _12883_/X sky130_fd_sc_hd__or2_1
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08983__B _08983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _11848_/A vssd1 vssd1 vccd1 vccd1 _11834_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ input60/X vssd1 vssd1 vccd1 vccd1 _12951_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _13504_/A vssd1 vssd1 vccd1 vccd1 _13518_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10716_ _10716_/A _10716_/B _10727_/C vssd1 vssd1 vccd1 vccd1 _10834_/B sky130_fd_sc_hd__and3_1
X_11696_ _13752_/Q _13751_/Q _11888_/B vssd1 vssd1 vccd1 vccd1 _11893_/B sky130_fd_sc_hd__or3_1
XFILLER_9_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13435_ _13444_/A _13435_/B vssd1 vssd1 vccd1 vccd1 _13436_/A sky130_fd_sc_hd__and2_1
X_10647_ _13952_/Q _10550_/X _10644_/X _10646_/X vssd1 vssd1 vccd1 vccd1 _13952_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10426__A_N _10399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13366_ _13375_/A _13366_/B vssd1 vssd1 vccd1 vccd1 _13367_/A sky130_fd_sc_hd__and2_1
XFILLER_6_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10578_ _10578_/A _10578_/B _10578_/C vssd1 vssd1 vccd1 vccd1 _10578_/X sky130_fd_sc_hd__or3_1
XFILLER_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12317_ _12317_/A vssd1 vssd1 vccd1 vccd1 _12322_/A sky130_fd_sc_hd__clkbuf_4
X_13297_ _14340_/Q _13289_/X _13296_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _14340_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12248_ _12251_/A vssd1 vssd1 vccd1 vccd1 _12248_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12179_ _13343_/A _12179_/B _12179_/C vssd1 vssd1 vccd1 vccd1 _12180_/A sky130_fd_sc_hd__and3_1
XFILLER_25_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14178__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08410_ _09751_/B _09751_/C _09751_/A vssd1 vssd1 vccd1 vccd1 _10523_/B sky130_fd_sc_hd__o21ai_1
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09390_ _09391_/A _09423_/B _09423_/C vssd1 vssd1 vccd1 vccd1 _09390_/X sky130_fd_sc_hd__and3_1
XFILLER_52_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08341_ _09751_/B _08341_/B vssd1 vssd1 vccd1 vccd1 _08343_/C sky130_fd_sc_hd__nor2_1
XFILLER_51_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11105__A _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08272_ _09777_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11091__A1 _11142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11091__B2 _10826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13368__A0 _12633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07223_ _07240_/A vssd1 vssd1 vccd1 vccd1 _07236_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13320__A _13341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ _07154_/A vssd1 vssd1 vccd1 vccd1 _14291_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_69_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08414__A _08905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07085_ _07085_/A vssd1 vssd1 vccd1 vccd1 _07085_/X sky130_fd_sc_hd__buf_4
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input1_A dout1[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07987_ _09553_/C vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06938_ _06938_/A vssd1 vssd1 vccd1 vccd1 _14318_/D sky130_fd_sc_hd__clkbuf_1
X_09726_ _09717_/X _09724_/A _09718_/A vssd1 vssd1 vccd1 vccd1 _09741_/A sky130_fd_sc_hd__a21o_1
XFILLER_68_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10657__A1 _10826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06869_ _06869_/A _06869_/B _06869_/C _06868_/X vssd1 vssd1 vccd1 vccd1 _06875_/C
+ sky130_fd_sc_hd__or4b_1
XANTENNA__11854__B1 _11823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _09187_/X _09190_/Y _09262_/X _09264_/Y vssd1 vssd1 vccd1 vccd1 _09657_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _08608_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08609_/B sky130_fd_sc_hd__xnor2_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13056__C1 _13053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09588_ _09548_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__and2b_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08539_ _08966_/A _08658_/B _08615_/B _08538_/A vssd1 vssd1 vccd1 vccd1 _08692_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11550_ _14041_/Q _13953_/Q vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__nor2_1
XFILLER_11_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ _10520_/C vssd1 vssd1 vccd1 vccd1 _10501_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ _08658_/B _11455_/X _11479_/Y _11480_/X vssd1 vssd1 vccd1 vccd1 _13871_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13220_ _14405_/Q _13216_/X _13219_/X vssd1 vssd1 vccd1 vccd1 _13220_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13230__A _13526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10432_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10433_/B sky130_fd_sc_hd__or2_1
XFILLER_104_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13151_ _13152_/A vssd1 vssd1 vccd1 vccd1 _13151_/Y sky130_fd_sc_hd__inv_2
X_10363_ _10364_/A _10364_/B _10364_/C vssd1 vssd1 vccd1 vccd1 _10378_/A sky130_fd_sc_hd__a21o_1
XFILLER_100_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12102_ input97/X vssd1 vssd1 vccd1 vccd1 _12926_/A sky130_fd_sc_hd__clkbuf_8
X_13082_ _13089_/A _13082_/B vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__and2_1
XANTENNA_input57_A io_wbs_adr[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _10297_/A _10297_/B _10297_/C vssd1 vssd1 vccd1 vccd1 _10374_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08978__B _08978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12033_ _12044_/A _12033_/B vssd1 vssd1 vccd1 vccd1 _12034_/A sky130_fd_sc_hd__and2_1
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07210__A0 _14275_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13984_ _13986_/CLK _13984_/D _12412_/Y vssd1 vssd1 vccd1 vccd1 _13984_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12935_ hold1/A _12928_/X _12932_/X _12934_/X vssd1 vssd1 vccd1 vccd1 _14160_/D sky130_fd_sc_hd__o211a_1
XFILLER_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _12920_/A vssd1 vssd1 vccd1 vccd1 _12866_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11817_ _13995_/Q _11809_/A _11800_/X _14114_/Q vssd1 vssd1 vccd1 vccd1 _11817_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _14156_/Q _12783_/X _12774_/A _14132_/Q vssd1 vssd1 vccd1 vccd1 _12797_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11745_/Y _14254_/Q _14255_/Q hold16/X vssd1 vssd1 vccd1 vccd1 _14254_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09018__A1 _09088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14467_ _14467_/CLK _14467_/D vssd1 vssd1 vccd1 vccd1 _14467_/Q sky130_fd_sc_hd__dfxtp_1
X_11679_ _11679_/A _11679_/B vssd1 vssd1 vccd1 vccd1 _11680_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06961__B _14282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13418_ _13418_/A vssd1 vssd1 vccd1 vccd1 _14372_/D sky130_fd_sc_hd__clkbuf_1
X_14398_ _14440_/CLK _14398_/D vssd1 vssd1 vccd1 vccd1 _14398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13349_ _14433_/Q _13216_/X _13348_/X _13341_/X vssd1 vssd1 vccd1 vccd1 _13349_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13522__A0 _12688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07910_ _07909_/A _07909_/B _07909_/C vssd1 vssd1 vccd1 vccd1 _07911_/B sky130_fd_sc_hd__a21oi_1
X_08890_ _08936_/A _10081_/A _09943_/B _08891_/A vssd1 vssd1 vccd1 vccd1 _08892_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__07201__A0 _14277_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07841_ _14029_/Q _13975_/Q vssd1 vssd1 vccd1 vccd1 _07900_/A sky130_fd_sc_hd__and2_1
XFILLER_57_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07772_ _13987_/Q _13986_/Q _13988_/Q vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__or3b_4
XFILLER_37_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09511_ _09511_/A _09511_/B _09511_/C vssd1 vssd1 vccd1 vccd1 _09511_/X sky130_fd_sc_hd__and3_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11534__S _11534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13315__A _13315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ _09553_/C _09848_/B _09369_/X _09286_/X _09804_/A vssd1 vssd1 vccd1 vccd1
+ _09447_/A sky130_fd_sc_hd__a32o_1
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13589__A0 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09373_ _09373_/A _09373_/B _09373_/C vssd1 vssd1 vccd1 vccd1 _09376_/A sky130_fd_sc_hd__nand3_1
XFILLER_21_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08128__B _08128_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08324_ _08380_/A _08380_/B _08380_/C vssd1 vssd1 vccd1 vccd1 _08324_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__07032__B _14273_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08255_ _09769_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _08257_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ _07240_/A vssd1 vssd1 vccd1 vccd1 _07219_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_119_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08186_ _09584_/A vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_118_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07137_ _07137_/A vssd1 vssd1 vccd1 vccd1 _14292_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07983__A _13872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _07051_/X _07067_/X _14356_/Q vssd1 vssd1 vccd1 vccd1 _07069_/S sky130_fd_sc_hd__o21a_1
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11827__B1 _11823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09709_ _09692_/A _09692_/C _09692_/B vssd1 vssd1 vccd1 vccd1 _09709_/X sky130_fd_sc_hd__o21a_1
X_10981_ _11011_/B _11012_/A _11008_/A _11005_/A vssd1 vssd1 vccd1 vccd1 _10999_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_74_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12720_ _12721_/A vssd1 vssd1 vccd1 vccd1 _12720_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ _12650_/X _14046_/Q _12665_/S vssd1 vssd1 vccd1 vccd1 _12652_/B sky130_fd_sc_hd__mux2_1
XFILLER_90_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07259__A0 _14260_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ _11602_/A _11602_/B vssd1 vssd1 vccd1 vccd1 _11602_/Y sky130_fd_sc_hd__xnor2_4
X_12582_ _12582_/A vssd1 vssd1 vccd1 vccd1 _14027_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321_ _14411_/CLK _14321_/D _13191_/Y vssd1 vssd1 vccd1 vccd1 _14321_/Q sky130_fd_sc_hd__dfrtp_4
X_11533_ _11134_/A _11355_/A _11533_/S vssd1 vssd1 vccd1 vccd1 _11533_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11464_ _11474_/A vssd1 vssd1 vccd1 vccd1 _11464_/X sky130_fd_sc_hd__clkbuf_2
X_14252_ _14259_/CLK _14252_/D vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12555__A1 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13203_ _13206_/A _13203_/B _13203_/C vssd1 vssd1 vccd1 vccd1 _13245_/A sky130_fd_sc_hd__and3_4
X_10415_ _10416_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10417_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14183_ _14256_/CLK _14183_/D _12970_/Y vssd1 vssd1 vccd1 vccd1 _14183_/Q sky130_fd_sc_hd__dfrtp_1
X_11395_ _13882_/Q _11392_/X _11383_/X _11394_/X vssd1 vssd1 vccd1 vccd1 _13882_/D
+ sky130_fd_sc_hd__a22o_1
X_13134_ _13134_/A vssd1 vssd1 vccd1 vccd1 _13134_/Y sky130_fd_sc_hd__inv_2
X_10346_ _10346_/A _10367_/B vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__nand2_1
XANTENNA_output163_A _14318_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13065_/A vssd1 vssd1 vccd1 vccd1 _14241_/D sky130_fd_sc_hd__clkbuf_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10277_ _10302_/A _10486_/S _10277_/S vssd1 vssd1 vccd1 vccd1 _10278_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12304__A _12304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _12016_/A vssd1 vssd1 vccd1 vccd1 _13787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13967_ _13988_/CLK _13967_/D _12391_/Y vssd1 vssd1 vccd1 vccd1 _13967_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12918_ _14154_/Q _12915_/X _12917_/X _12907_/X vssd1 vssd1 vccd1 vccd1 _14154_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13898_ _13905_/CLK _13898_/D _12306_/Y vssd1 vssd1 vccd1 vccd1 _13898_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _13072_/A vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12794__A1 _14155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14366__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08040_ _08716_/B _08043_/A _08039_/A vssd1 vssd1 vccd1 vccd1 _08146_/A sky130_fd_sc_hd__a21oi_4
XFILLER_31_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11349__A2 _10845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09991_ _09921_/A _09921_/B _09990_/X vssd1 vssd1 vccd1 vccd1 _09993_/B sky130_fd_sc_hd__a21oi_1
XFILLER_118_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ _08949_/B _08950_/B _08949_/A vssd1 vssd1 vccd1 vccd1 _08942_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08873_ _08830_/A _08829_/A _08829_/B vssd1 vssd1 vccd1 vccd1 _08875_/A sky130_fd_sc_hd__o21ba_1
XFILLER_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13744__S _13744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07824_ _14031_/Q _13977_/Q vssd1 vssd1 vccd1 vccd1 _07824_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07755_ _07676_/X _07723_/X _07724_/X vssd1 vssd1 vccd1 vccd1 _07755_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10669__A _10826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06866__B _13778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _07688_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _07686_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09425_ _09425_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09427_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _09465_/A _09455_/A _09356_/C vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__nand3_1
XFILLER_100_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08307_ _09165_/C vssd1 vssd1 vccd1 vccd1 _09473_/B sky130_fd_sc_hd__clkbuf_2
X_09287_ _09286_/B _09881_/A _09207_/C _09286_/A vssd1 vssd1 vccd1 vccd1 _09287_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08238_ _09712_/A vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__buf_2
XFILLER_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12537__A1 _08842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08169_ _08245_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08170_/C sky130_fd_sc_hd__xnor2_1
XFILLER_107_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10200_ _10200_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10202_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ _10765_/B _11163_/X _11140_/X vssd1 vssd1 vccd1 vccd1 _11180_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08602__A _09055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10851__B _10851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ _10157_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10136_/A sky130_fd_sc_hd__and2_1
XANTENNA__10563__A3 _10561_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10062_ _10070_/A _10060_/X _10061_/X vssd1 vssd1 vccd1 vccd1 _10063_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_47_io_wbs_clk clkbuf_3_5_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13820_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13821_ _14348_/CLK _13821_/D vssd1 vssd1 vccd1 vccd1 _13821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11174__S _11175_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13752_ _13826_/CLK _13752_/D _11940_/Y vssd1 vssd1 vccd1 vccd1 _13752_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ _13905_/Q _13906_/Q _13907_/Q _13908_/Q _10960_/S _10662_/A vssd1 vssd1 vccd1
+ vccd1 _10964_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08049__A _08146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12703_ _12703_/A vssd1 vssd1 vccd1 vccd1 _12703_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ _13683_/A vssd1 vssd1 vccd1 vccd1 _14448_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10895_ _13972_/Q _10895_/B vssd1 vssd1 vccd1 vccd1 _10895_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12634_ _12633_/X _14042_/Q _12642_/S vssd1 vssd1 vccd1 vccd1 _12635_/B sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_59_io_wbs_clk_A clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12565_ _10614_/A _12520_/S _11935_/A vssd1 vssd1 vccd1 vccd1 _12565_/Y sky130_fd_sc_hd__a21oi_1
X_14304_ _14304_/CLK _14304_/D _13171_/Y vssd1 vssd1 vccd1 vccd1 _14304_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11516_ _08918_/B _11510_/X _11512_/X _11515_/X vssd1 vssd1 vccd1 vccd1 _13864_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ _09762_/A _12486_/X _12476_/A _14054_/Q vssd1 vssd1 vccd1 vccd1 _12496_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13725__A0 input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14235_ _14239_/CLK _14235_/D vssd1 vssd1 vccd1 vccd1 _14235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11447_ _11447_/A vssd1 vssd1 vccd1 vccd1 _11447_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09944__A2 _10191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ _14283_/CLK _14166_/D _12947_/Y vssd1 vssd1 vccd1 vccd1 _14166_/Q sky130_fd_sc_hd__dfrtp_4
X_11378_ hold35/A _11363_/X _11370_/X _11377_/X vssd1 vssd1 vccd1 vccd1 _13888_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08512__A _13863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13121_/A vssd1 vssd1 vccd1 vccd1 _13117_/Y sky130_fd_sc_hd__inv_2
X_10329_ _09968_/A _10302_/B _10328_/Y vssd1 vssd1 vccd1 vccd1 _10341_/A sky130_fd_sc_hd__o21ai_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14097_ _14102_/CLK _14097_/D _12746_/Y vssd1 vssd1 vccd1 vccd1 _14097_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13048_ _14235_/Q _13041_/X _13047_/X _13039_/X vssd1 vssd1 vccd1 vccd1 _14235_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07707__A1 _14148_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07540_ _14172_/Q _14171_/Q vssd1 vssd1 vccd1 vccd1 _07541_/C sky130_fd_sc_hd__and2_1
XFILLER_46_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07471_ _07471_/A vssd1 vssd1 vccd1 vccd1 _07471_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_90_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09210_ _09210_/A _09210_/B vssd1 vssd1 vccd1 vccd1 _09212_/B sky130_fd_sc_hd__xnor2_4
XFILLER_72_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12767__A1 hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13756__CLK _13825_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09141_ _09140_/A _09140_/C _09140_/B vssd1 vssd1 vccd1 vccd1 _09141_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12209__A _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ _09072_/A _09072_/B vssd1 vssd1 vccd1 vccd1 _09081_/A sky130_fd_sc_hd__nand2_1
X_08023_ _08024_/B _08024_/C _08024_/A vssd1 vssd1 vccd1 vccd1 _08325_/A sky130_fd_sc_hd__a21o_1
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08422__A _09457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_61_io_wbs_clk_A clkbuf_3_7_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_115_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _10274_/B _09974_/B vssd1 vssd1 vccd1 vccd1 _09980_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08925_ _08925_/A _08936_/A _08925_/C _10057_/A vssd1 vssd1 vccd1 vccd1 _08928_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_103_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12879__A _12920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08856_ _08856_/A _08856_/B _08856_/C vssd1 vssd1 vccd1 vccd1 _08856_/X sky130_fd_sc_hd__and3_1
XFILLER_111_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06877__A _06970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08371__A1 _08842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07807_ _14007_/Q _10690_/S vssd1 vssd1 vccd1 vccd1 _07807_/Y sky130_fd_sc_hd__nor2_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08787_ _08787_/A _08787_/B _08787_/C vssd1 vssd1 vccd1 vccd1 _08799_/A sky130_fd_sc_hd__or3_1
XFILLER_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _07665_/Y _07723_/X _07724_/X vssd1 vssd1 vccd1 vccd1 _07738_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11007__B _11007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07669_ _07669_/A _07640_/Y vssd1 vssd1 vccd1 vccd1 _07670_/B sky130_fd_sc_hd__or2b_1
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09408_ _09690_/A _09408_/B vssd1 vssd1 vccd1 vccd1 _09408_/X sky130_fd_sc_hd__or2_1
X_10680_ _10967_/S vssd1 vssd1 vccd1 vccd1 _11155_/S sky130_fd_sc_hd__buf_2
XFILLER_90_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09339_ _09274_/B _09274_/Y _09337_/Y _09338_/X vssd1 vssd1 vccd1 vccd1 _09339_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12119__A _12147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11430__A1 _11010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ _12353_/A vssd1 vssd1 vccd1 vccd1 _12350_/Y sky130_fd_sc_hd__inv_2
X_11301_ _11317_/B _11317_/C _11317_/A vssd1 vssd1 vccd1 vccd1 _11315_/C sky130_fd_sc_hd__o21ai_1
X_12281_ _12285_/A vssd1 vssd1 vccd1 vccd1 _12281_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _11240_/B _11241_/A _11237_/A _11236_/A vssd1 vssd1 vccd1 vccd1 _11233_/B
+ sky130_fd_sc_hd__a31o_1
X_14020_ _14020_/CLK _14020_/D vssd1 vssd1 vccd1 vccd1 _14020_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ _13924_/Q _13925_/Q _10912_/A _13927_/Q _10679_/A _10721_/C vssd1 vssd1 vccd1
+ vccd1 _11163_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _10114_/A _10114_/B vssd1 vssd1 vccd1 vccd1 _10115_/B sky130_fd_sc_hd__nor2_1
X_11094_ _11083_/A _11084_/X _11093_/Y vssd1 vssd1 vccd1 vccd1 _11094_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10045_ _10045_/A _10122_/A vssd1 vssd1 vccd1 vccd1 _10045_/X sky130_fd_sc_hd__or2_1
XFILLER_102_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13804_ _14348_/CLK _13804_/D vssd1 vssd1 vccd1 vccd1 _13804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11996_ _12059_/A vssd1 vssd1 vccd1 vccd1 _12000_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_91_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13735_ input86/X _14464_/Q _13738_/S vssd1 vssd1 vccd1 vccd1 _13736_/B sky130_fd_sc_hd__mux2_1
X_10947_ _10953_/A _10944_/X _10945_/X _10946_/X _10771_/Y vssd1 vssd1 vccd1 vccd1
+ _10947_/X sky130_fd_sc_hd__o2111a_1
XFILLER_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13666_ _13666_/A vssd1 vssd1 vccd1 vccd1 _14443_/D sky130_fd_sc_hd__clkbuf_1
X_10878_ _10878_/A vssd1 vssd1 vccd1 vccd1 _13934_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12617_ _12637_/A vssd1 vssd1 vccd1 vccd1 _12635_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13597_ input78/X _14424_/Q _13611_/S vssd1 vssd1 vccd1 vccd1 _13598_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12548_ _12551_/A _12548_/B vssd1 vssd1 vccd1 vccd1 _12549_/A sky130_fd_sc_hd__and2_1
XANTENNA__13559__S _13559_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12479_ _12817_/A vssd1 vssd1 vccd1 vccd1 _12479_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14218_ _14284_/CLK _14218_/D _13014_/Y vssd1 vssd1 vccd1 vccd1 _14218_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_1_0_io_wbs_clk clkbuf_2_1_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_io_wbs_clk/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14404__CLK _14440_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12921__A1 _14155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A2 _11872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14149_ _14149_/CLK _14149_/D vssd1 vssd1 vccd1 vccd1 _14149_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09057__B _09233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _14425_/Q _06969_/Y _06970_/X vssd1 vssd1 vccd1 vccd1 _06971_/X sky130_fd_sc_hd__a21o_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08896__B _10171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ _08532_/A _08531_/B _08531_/C vssd1 vssd1 vccd1 vccd1 _08719_/C sky130_fd_sc_hd__a21o_1
XFILLER_6_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12685__A0 _12940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09690_ _09690_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09692_/B sky130_fd_sc_hd__xnor2_1
XFILLER_67_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09550__B1 _09818_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09073__A _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08641_ _08641_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08997_/B sky130_fd_sc_hd__nor2_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12211__B input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11108__A _11108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08572_ _13859_/Q vssd1 vssd1 vccd1 vccd1 _09084_/D sky130_fd_sc_hd__clkbuf_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07523_ _14185_/Q _14178_/Q _07520_/Y vssd1 vssd1 vccd1 vccd1 _07523_/X sky130_fd_sc_hd__o21a_1
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07454_ _07458_/A _07454_/B vssd1 vssd1 vccd1 vccd1 _07454_/X sky130_fd_sc_hd__or2_1
XFILLER_23_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07959__C _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__A _13866_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07321__A _07376_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07385_ _14213_/Q _07373_/X _07375_/X _07384_/X vssd1 vssd1 vccd1 vccd1 _14213_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09124_ _13871_/Q vssd1 vssd1 vccd1 vccd1 _09553_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_109_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07092__A1 _07090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09055_ _09055_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09056_/B sky130_fd_sc_hd__nand2_1
X_08006_ _14019_/Q vssd1 vssd1 vccd1 vccd1 _08623_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_81_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09957_ _09957_/A _09956_/A vssd1 vssd1 vccd1 vccd1 _09957_/X sky130_fd_sc_hd__or2b_1
XFILLER_89_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08908_ _08908_/A _08908_/B vssd1 vssd1 vccd1 vccd1 _08915_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09888_ _10050_/B _10059_/A vssd1 vssd1 vccd1 vccd1 _10157_/A sky130_fd_sc_hd__xor2_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08344__A1 _09425_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08839_ _08839_/A _08839_/B vssd1 vssd1 vccd1 vccd1 _08859_/A sky130_fd_sc_hd__nand2_1
XFILLER_79_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11018__A _11061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _14343_/Q _11847_/X _11848_/X _13802_/Q vssd1 vssd1 vccd1 vccd1 _11850_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _10868_/B _10801_/B vssd1 vssd1 vccd1 vccd1 _10873_/A sky130_fd_sc_hd__nor2_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _11768_/A _11780_/X _11767_/B vssd1 vssd1 vccd1 vccd1 _11823_/A sky130_fd_sc_hd__a21bo_2
XFILLER_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13520_ _13609_/A vssd1 vssd1 vccd1 vccd1 _13592_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10732_ _13938_/Q _10812_/B vssd1 vssd1 vccd1 vccd1 _10846_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13451_ input84/X _14382_/Q _13460_/S vssd1 vssd1 vccd1 vccd1 _13452_/B sky130_fd_sc_hd__mux2_1
X_10663_ _10777_/B _10670_/B _11164_/S vssd1 vssd1 vccd1 vccd1 _10663_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_90_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07607__A0 _14080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12402_ _12403_/A vssd1 vssd1 vccd1 vccd1 _12402_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12600__A0 _12926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input87_A io_wbs_datwr[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13382_ _12650_/X _14362_/Q _13391_/S vssd1 vssd1 vccd1 vccd1 _13383_/B sky130_fd_sc_hd__mux2_1
X_10594_ _10565_/B _10589_/Y _10593_/Y _09788_/X vssd1 vssd1 vccd1 vccd1 _10594_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_103_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07083__A1 _14299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ _12335_/A vssd1 vssd1 vccd1 vccd1 _12333_/Y sky130_fd_sc_hd__inv_2
X_12264_ _12267_/A vssd1 vssd1 vccd1 vccd1 _12264_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08062__A _13873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14003_ _14442_/CLK _14003_/D vssd1 vssd1 vccd1 vccd1 _14003_/Q sky130_fd_sc_hd__dfxtp_1
X_11215_ _13906_/Q vssd1 vssd1 vccd1 vccd1 _11297_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12195_ input55/X input58/X vssd1 vssd1 vccd1 vccd1 _12196_/C sky130_fd_sc_hd__or2b_1
X_11146_ _13923_/Q _13924_/Q _13925_/Q _13926_/Q _11169_/S _07798_/A vssd1 vssd1 vccd1
+ vccd1 _11146_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11077_ _11099_/B _11077_/B vssd1 vssd1 vccd1 vccd1 _11102_/A sky130_fd_sc_hd__and2_1
XFILLER_48_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07406__A _07460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _10027_/B _10028_/B vssd1 vssd1 vccd1 vccd1 _10028_/X sky130_fd_sc_hd__and2b_1
XFILLER_49_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06897__A1 _06894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11870__B _11870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11979_ _12233_/A vssd1 vssd1 vccd1 vccd1 _11979_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09835__A1 _08291_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__A _11020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13143__A _13146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ input81/X _14459_/Q _13721_/S vssd1 vssd1 vccd1 vccd1 _13719_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08237__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07779__C _10585_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13649_ _13649_/A vssd1 vssd1 vccd1 vccd1 _14438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07170_ _07259_/S vssd1 vssd1 vccd1 vccd1 _07183_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_9_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10007__A _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09811_ _09811_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09811_/X sky130_fd_sc_hd__and2_1
XFILLER_8_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ _09742_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _10541_/A sky130_fd_sc_hd__or2_2
X_06954_ _14459_/Q _14283_/Q vssd1 vssd1 vccd1 vccd1 _06954_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09673_ _09673_/A _09673_/B vssd1 vssd1 vccd1 vccd1 _09690_/B sky130_fd_sc_hd__xnor2_1
X_06885_ _14395_/Q _06855_/Y _06865_/Y _14389_/Q _06884_/X vssd1 vssd1 vccd1 vccd1
+ _06885_/X sky130_fd_sc_hd__a221o_1
XFILLER_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08623_/B _09085_/B _09084_/C _08623_/A vssd1 vssd1 vccd1 vccd1 _08625_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06888__A1 _14393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06888__B2 _14392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09531__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08555_ _09001_/A _08555_/B _09870_/A _08863_/D vssd1 vssd1 vccd1 vccd1 _08555_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06874__B _14269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13053__A _13254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ hold25/X _14184_/Q _07506_/S vssd1 vssd1 vccd1 vccd1 _07507_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08486_ _13860_/Q vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07051__A _07090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07437_ _07464_/A vssd1 vssd1 vccd1 vccd1 _07458_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12892__A _12920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__A _14018_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07368_ _14216_/Q _07347_/X _07348_/X _07367_/X vssd1 vssd1 vccd1 vccd1 _14216_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07065__A1 _14260_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09107_ _09119_/B _09106_/B _09106_/C _09106_/D vssd1 vssd1 vccd1 vccd1 _09107_/X
+ sky130_fd_sc_hd__o22a_1
X_07299_ _07298_/Y _14192_/D _07307_/A vssd1 vssd1 vccd1 vccd1 _14226_/D sky130_fd_sc_hd__o21bai_1
X_09038_ _09038_/A _09038_/B vssd1 vssd1 vccd1 vccd1 _09038_/Y sky130_fd_sc_hd__nor2_1
XFILLER_117_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11000_ _11000_/A _11000_/B vssd1 vssd1 vccd1 vccd1 _11073_/B sky130_fd_sc_hd__xnor2_1
XFILLER_105_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13228__A _13254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09425__B _09811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12951_ _12951_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _13197_/A sky130_fd_sc_hd__or2_4
XFILLER_92_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08868__A2 _08925_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11971__A _11971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11902_ _13756_/Q _11902_/B vssd1 vssd1 vccd1 vccd1 _11903_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06879__A1 _14269_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _14141_/Q _12872_/X _12881_/X _12879_/X vssd1 vssd1 vccd1 vccd1 _14141_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_34_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _11833_/A vssd1 vssd1 vccd1 vccd1 _11833_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11624__A1 _11623_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _12440_/A vssd1 vssd1 vccd1 vccd1 _11809_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08057__A _13871_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13503_ _13503_/A vssd1 vssd1 vccd1 vccd1 _14397_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10715_/A _10761_/B _10761_/C vssd1 vssd1 vccd1 vccd1 _10727_/C sky130_fd_sc_hd__or3_2
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11695_ _13750_/Q _11883_/B vssd1 vssd1 vccd1 vccd1 _11888_/B sky130_fd_sc_hd__or2_2
X_13434_ input79/X _14377_/Q _13443_/S vssd1 vssd1 vccd1 vccd1 _13435_/B sky130_fd_sc_hd__mux2_1
X_10646_ _10565_/B _10636_/B _10645_/Y _09788_/A vssd1 vssd1 vccd1 vccd1 _10646_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_10_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13365_ _13084_/X hold33/A _13374_/S vssd1 vssd1 vccd1 vccd1 _13366_/B sky130_fd_sc_hd__mux2_1
X_10577_ _10576_/B _10576_/C _10576_/A vssd1 vssd1 vccd1 vccd1 _10578_/C sky130_fd_sc_hd__a21oi_1
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12316_ _12316_/A vssd1 vssd1 vccd1 vccd1 _12316_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13296_ _14420_/Q _13284_/X _13295_/X _13258_/X vssd1 vssd1 vccd1 vccd1 _13296_/X
+ sky130_fd_sc_hd__a211o_1
X_12247_ _12251_/A vssd1 vssd1 vccd1 vccd1 _12247_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12178_ _11990_/B _12092_/Y _11920_/A vssd1 vssd1 vccd1 vccd1 _12179_/C sky130_fd_sc_hd__a21o_1
XFILLER_25_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11129_ _11129_/A _11129_/B vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09808__A1 _08794_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ _08194_/X _08338_/Y _08336_/A _08337_/Y vssd1 vssd1 vccd1 vccd1 _08341_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_33_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08271_ _08271_/A _08271_/B vssd1 vssd1 vccd1 vccd1 _08272_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13368__A1 _14358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07222_ _14087_/Q _13887_/Q _07235_/S vssd1 vssd1 vccd1 vccd1 _07222_/X sky130_fd_sc_hd__mux2_2
XFILLER_118_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07153_ _14291_/Q _07144_/X _07165_/S vssd1 vssd1 vccd1 vccd1 _07154_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08795__B2 _08828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ _07084_/A vssd1 vssd1 vccd1 vccd1 _14299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11146__A3 _13926_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__B input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07986_ _14018_/Q vssd1 vssd1 vccd1 vccd1 _09553_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07770__A2 _07185_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07046__A _07085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09725_ _10557_/A _10557_/B _10557_/C _09718_/X _10566_/B vssd1 vssd1 vccd1 vccd1
+ _09725_/X sky130_fd_sc_hd__a311o_2
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06937_ _06933_/X _14318_/Q _06937_/S vssd1 vssd1 vccd1 vccd1 _06938_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12887__A _12930_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11791__A _11791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09656_ _10644_/B _09117_/Y _09421_/Y _10632_/A _09662_/A vssd1 vssd1 vccd1 vccd1
+ _10557_/A sky130_fd_sc_hd__a2111o_1
XANTENNA__10657__A2 _10705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06868_ _14398_/Q _06864_/Y _06865_/Y _14397_/Q vssd1 vssd1 vccd1 vccd1 _06868_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08607_ _08607_/A _08607_/B vssd1 vssd1 vccd1 vccd1 _08669_/B sky130_fd_sc_hd__xor2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09587_ _09514_/A _09537_/B _08110_/X vssd1 vssd1 vccd1 vccd1 _09591_/A sky130_fd_sc_hd__o21ba_1
XFILLER_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08615_/B sky130_fd_sc_hd__nor2_1
XFILLER_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08308__C _09803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08469_ _08469_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08470_/B sky130_fd_sc_hd__nor2_1
X_10500_ _10508_/A _10507_/B vssd1 vssd1 vccd1 vccd1 _10520_/C sky130_fd_sc_hd__and2b_1
X_11480_ _11076_/A _11460_/X _11475_/X _11297_/A _11461_/X vssd1 vssd1 vccd1 vccd1
+ _11480_/X sky130_fd_sc_hd__o221a_1
XFILLER_52_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10431_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10449_/B sky130_fd_sc_hd__nand2_1
XFILLER_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13150_ _13152_/A vssd1 vssd1 vccd1 vccd1 _13150_/Y sky130_fd_sc_hd__inv_2
X_10362_ _10362_/A _10414_/S vssd1 vssd1 vccd1 vccd1 _10364_/C sky130_fd_sc_hd__xnor2_1
XFILLER_87_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12101_ hold24/A _12095_/X _12100_/X _11931_/X vssd1 vssd1 vccd1 vccd1 _13807_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13657__S _13670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11966__A _13153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13081_ _12827_/X hold27/A _13096_/S vssd1 vssd1 vccd1 vccd1 _13082_/B sky130_fd_sc_hd__mux2_1
X_10293_ _10293_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10297_/C sky130_fd_sc_hd__xnor2_1
XFILLER_88_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12032_ _13792_/Q _12020_/X _12021_/X hold36/A vssd1 vssd1 vccd1 vccd1 _12033_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08978__C _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07210__A1 _07209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13983_ _13987_/CLK _13983_/D _12411_/Y vssd1 vssd1 vccd1 vccd1 _13983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12934_ _13254_/A vssd1 vssd1 vccd1 vccd1 _12934_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _12933_/A vssd1 vssd1 vccd1 vccd1 _12920_/A sky130_fd_sc_hd__buf_2
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _13788_/Q _11793_/X _11815_/X vssd1 vssd1 vccd1 vccd1 _11816_/X sky130_fd_sc_hd__a21o_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _14114_/Q _12782_/X _12794_/X _12795_/X _12216_/X vssd1 vssd1 vccd1 vccd1
+ _14114_/D sky130_fd_sc_hd__o221a_1
XFILLER_15_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _12205_/A _07146_/B _14259_/Q _11746_/X vssd1 vssd1 vccd1 vccd1 hold16/A
+ sky130_fd_sc_hd__o31a_2
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14466_ _14467_/CLK _14466_/D vssd1 vssd1 vccd1 vccd1 _14466_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08515__A _09234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09018__A2 _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11678_ _13777_/Q _13776_/Q _11682_/B _13778_/Q vssd1 vssd1 vccd1 vccd1 _11680_/B
+ sky130_fd_sc_hd__a31o_1
X_13417_ _13426_/A _13417_/B vssd1 vssd1 vccd1 vccd1 _13418_/A sky130_fd_sc_hd__and2_1
X_10629_ _13954_/Q _10628_/X _10629_/S vssd1 vssd1 vccd1 vccd1 _10630_/A sky130_fd_sc_hd__mux2_1
X_14397_ _14440_/CLK _14397_/D vssd1 vssd1 vccd1 vccd1 _14397_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12022__B2 _13829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13348_ _14385_/Q _13236_/A _13336_/X _14465_/Q vssd1 vssd1 vccd1 vccd1 _13348_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10584__B2 _10547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13279_ _14336_/Q _13265_/X _13277_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _14336_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_64_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08250__A _09762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__A1 _09969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_66_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_29_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07840_ _07840_/A _07840_/B vssd1 vssd1 vccd1 vccd1 _07901_/B sky130_fd_sc_hd__and2_1
XFILLER_96_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07771_ _11362_/A _07921_/C vssd1 vssd1 vccd1 vccd1 _07779_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09510_ _08098_/X _09510_/B _09510_/C vssd1 vssd1 vccd1 vccd1 _09511_/C sky130_fd_sc_hd__nand3b_1
XFILLER_83_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09441_ _09441_/A _09385_/A vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__or2b_1
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10020__A _10092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ _09367_/A _09367_/B _09367_/C vssd1 vssd1 vccd1 vccd1 _09373_/C sky130_fd_sc_hd__a21o_1
XFILLER_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08323_ _08323_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08380_/C sky130_fd_sc_hd__xor2_2
XANTENNA__08128__C _10000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__B1 _08703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08254_ _09755_/A _09755_/B vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08425__A _13864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07205_ _14092_/Q _13892_/Q _07218_/S vssd1 vssd1 vccd1 vccd1 _07205_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08185_ _08937_/B _08093_/A _08091_/A vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__a21oi_4
X_07136_ _07133_/X _14292_/Q _07136_/S vssd1 vssd1 vccd1 vccd1 _07137_/A sky130_fd_sc_hd__mux2_1
XFILLER_106_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11786__A _11786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ _14404_/Q _07098_/B _14436_/Q vssd1 vssd1 vccd1 vccd1 _07067_/X sky130_fd_sc_hd__and3b_1
XANTENNA__07440__A1 _14086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_io_wbs_clk clkbuf_3_4_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14417_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_82_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07969_ _07969_/A _07969_/B vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__xnor2_1
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09708_ _09708_/A _09708_/B _09708_/C vssd1 vssd1 vccd1 vccd1 _09708_/Y sky130_fd_sc_hd__nand3_1
XFILLER_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _10651_/A _10958_/X _10920_/A vssd1 vssd1 vccd1 vccd1 _11005_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12410__A _12410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09655_/B sky130_fd_sc_hd__xnor2_2
XFILLER_83_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12650_ input94/X vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__buf_4
XFILLER_15_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14018__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11601_ _11601_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11602_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12581_ _12594_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__and2_1
XFILLER_12_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14320_ _14322_/CLK _14320_/D _13190_/Y vssd1 vssd1 vccd1 vccd1 _14320_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11532_ _08937_/C _11510_/X _11530_/X _11531_/X vssd1 vssd1 vccd1 vccd1 _13860_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14251_ _14259_/CLK _14251_/D vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12004__B2 _13824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11463_ _09188_/B _11455_/X _11462_/X vssd1 vssd1 vccd1 vccd1 _13874_/D sky130_fd_sc_hd__a21o_1
XFILLER_99_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13202_ _13202_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _13203_/C sky130_fd_sc_hd__nand2_1
XFILLER_87_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10414_ _10478_/A _10362_/A _10414_/S vssd1 vssd1 vccd1 vccd1 _10416_/B sky130_fd_sc_hd__mux2_1
X_14182_ _14256_/CLK _14182_/D _12969_/Y vssd1 vssd1 vccd1 vccd1 _14182_/Q sky130_fd_sc_hd__dfrtp_1
X_11394_ hold19/X _11403_/B vssd1 vssd1 vccd1 vccd1 _11394_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_76_io_wbs_clk clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14075_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_13133_ _13134_/A vssd1 vssd1 vccd1 vccd1 _13133_/Y sky130_fd_sc_hd__inv_2
X_10345_ _10345_/A _10345_/B vssd1 vssd1 vccd1 vccd1 _10367_/B sky130_fd_sc_hd__xor2_1
XFILLER_87_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09166__A _09297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _13070_/A _13064_/B vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__and2_1
XFILLER_78_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10276_ _10487_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10277_/S sky130_fd_sc_hd__nor2_1
XANTENNA_output156_A _14311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12015_ _12026_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _12016_/A sky130_fd_sc_hd__and2_1
XFILLER_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07195__A0 _14279_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13966_ _14031_/CLK _13966_/D _12390_/Y vssd1 vssd1 vccd1 vccd1 _13966_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12917_ _12917_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _12917_/X sky130_fd_sc_hd__or2_1
XANTENNA__12491__A1 _14036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ _13897_/CLK _13897_/D _12304_/Y vssd1 vssd1 vccd1 vccd1 _13897_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12848_ _12848_/A vssd1 vssd1 vccd1 vccd1 _14130_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13440__A0 input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ _14151_/Q _12772_/X _12774_/X _14127_/Q vssd1 vssd1 vccd1 vccd1 _12779_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14449_ _14449_/CLK _14449_/D vssd1 vssd1 vccd1 vccd1 _14449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09990_ _09920_/B _09990_/B vssd1 vssd1 vccd1 vccd1 _09990_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09076__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08941_ _08941_/A _08941_/B _08941_/C vssd1 vssd1 vccd1 vccd1 _08949_/A sky130_fd_sc_hd__nand3_1
XFILLER_103_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _08872_/A _08872_/B _08872_/C vssd1 vssd1 vccd1 vccd1 _08908_/A sky130_fd_sc_hd__and3_1
XFILLER_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07823_ _14032_/Q _13978_/Q vssd1 vssd1 vccd1 vccd1 _07847_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09804__A _09804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07754_ _14152_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07754_/X sky130_fd_sc_hd__and2_1
XANTENNA__12230__A _12517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07324__A _14107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12482__A1 _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07685_ _07685_/A _07685_/B vssd1 vssd1 vccd1 vccd1 _07688_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09424_ _09424_/A _09424_/B _09881_/B _09806_/A vssd1 vssd1 vccd1 vccd1 _09427_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_53_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13431__A0 input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09355_ _09354_/A _09354_/B _09354_/C vssd1 vssd1 vccd1 vccd1 _09356_/C sky130_fd_sc_hd__a21o_1
X_08306_ _13867_/Q vssd1 vssd1 vccd1 vccd1 _09165_/C sky130_fd_sc_hd__clkbuf_2
X_09286_ _09286_/A _09286_/B _09881_/A vssd1 vssd1 vccd1 vccd1 _09286_/X sky130_fd_sc_hd__and3_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ _09634_/A vssd1 vssd1 vccd1 vccd1 _09712_/A sky130_fd_sc_hd__buf_2
XFILLER_101_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08168_ _08168_/A _08168_/B vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__nor2_1
XFILLER_4_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07119_ _14291_/Q _07085_/X _07118_/X _14387_/Q vssd1 vssd1 vccd1 vccd1 _07119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08099_ _14014_/Q vssd1 vssd1 vccd1 vccd1 _08750_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10130_ _10283_/A _10135_/B _10129_/Y vssd1 vssd1 vccd1 vccd1 _10166_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__13498__A0 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10061_ _10061_/A _10069_/A vssd1 vssd1 vccd1 vccd1 _10061_/X sky130_fd_sc_hd__and2_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07177__A0 _14284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13820_ _13820_/CLK _13820_/D vssd1 vssd1 vccd1 vccd1 _13820_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13236__A _13236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13751_ _13826_/CLK _13751_/D _11939_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Q sky130_fd_sc_hd__dfrtp_1
X_10963_ _11134_/B _10963_/B _10963_/C _11039_/A vssd1 vssd1 vccd1 vccd1 _10970_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__13670__A0 _12664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13670__S _13670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12702_ _12703_/A vssd1 vssd1 vccd1 vccd1 _12702_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13682_ _13695_/A _13682_/B vssd1 vssd1 vccd1 vccd1 _13683_/A sky130_fd_sc_hd__and2_1
XFILLER_44_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10894_ _10894_/A _10894_/B _10894_/C vssd1 vssd1 vccd1 vccd1 _10894_/X sky130_fd_sc_hd__and3_1
XFILLER_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12633_ input88/X vssd1 vssd1 vccd1 vccd1 _12633_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12225__A1 _12906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13422__A0 input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ _12564_/A vssd1 vssd1 vccd1 vccd1 _14022_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14303_ _14367_/CLK _14303_/D _13170_/Y vssd1 vssd1 vccd1 vccd1 _14303_/Q sky130_fd_sc_hd__dfrtp_4
X_11515_ _11056_/A _11513_/X _11499_/X _11276_/A _11514_/X vssd1 vssd1 vccd1 vccd1
+ _11515_/X sky130_fd_sc_hd__o221a_1
XFILLER_8_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12495_ _14002_/Q _12481_/X _12494_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _14002_/D
+ sky130_fd_sc_hd__o211a_1
X_14234_ _14239_/CLK _14234_/D vssd1 vssd1 vccd1 vccd1 _14234_/Q sky130_fd_sc_hd__dfxtp_1
X_11446_ _11457_/A _10912_/A _11446_/S vssd1 vssd1 vccd1 vccd1 _11447_/A sky130_fd_sc_hd__mux2_1
X_14165_ _14283_/CLK _14165_/D _12946_/Y vssd1 vssd1 vccd1 vccd1 _14165_/Q sky130_fd_sc_hd__dfrtp_2
X_11377_ _13852_/Q _11377_/B vssd1 vssd1 vccd1 vccd1 _11377_/X sky130_fd_sc_hd__or2_1
XFILLER_4_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13116_ _13116_/A vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__buf_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _10421_/B _10328_/B vssd1 vssd1 vccd1 vccd1 _10328_/Y sky130_fd_sc_hd__nand2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14096_ _14104_/CLK _14096_/D _12745_/Y vssd1 vssd1 vccd1 vccd1 _14096_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _14243_/Q _13036_/S _13042_/Y hold32/A _13032_/A vssd1 vssd1 vccd1 vccd1
+ _13047_/X sky130_fd_sc_hd__a221o_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10259_ _10259_/A _10259_/B vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13146__A _13146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13949_ _13949_/CLK _13949_/D _12369_/Y vssd1 vssd1 vccd1 vccd1 _13949_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07470_ _07483_/A _07470_/B vssd1 vssd1 vccd1 vccd1 _07470_/X sky130_fd_sc_hd__or2_1
XFILLER_22_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13413__A0 _12688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _09140_/A _09140_/B _09140_/C vssd1 vssd1 vccd1 vccd1 _09140_/X sky130_fd_sc_hd__and3_1
XANTENNA__09093__B1 _08494_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09071_ _09071_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09071_/X sky130_fd_sc_hd__or2_1
X_08022_ _08054_/A _08054_/B vssd1 vssd1 vccd1 vccd1 _08024_/A sky130_fd_sc_hd__xnor2_1
XFILLER_116_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08703__A _09134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09973_ _10151_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__and2_1
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08924_ _08924_/A _08924_/B vssd1 vssd1 vccd1 vccd1 _08924_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07159__A0 _14289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08855_ _08818_/A _08816_/Y _08814_/X _08815_/X vssd1 vssd1 vccd1 vccd1 _08856_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08371__A2 _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ _10655_/A _07806_/B _11452_/B vssd1 vssd1 vccd1 vccd1 _10690_/S sky130_fd_sc_hd__or3_2
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08786_ _08785_/A _08785_/B _08785_/C vssd1 vssd1 vccd1 vccd1 _08801_/B sky130_fd_sc_hd__a21o_1
XFILLER_45_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10399__B _10399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _14157_/Q _07754_/B vssd1 vssd1 vccd1 vccd1 _07737_/X sky130_fd_sc_hd__and2_1
XANTENNA__12455__A1 _08896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07989__A _13874_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ _14140_/Q _07740_/A vssd1 vssd1 vccd1 vccd1 _07668_/X sky130_fd_sc_hd__or2_1
XANTENNA__06893__A _07090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09871__A2 _10083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09407_ _09404_/X _09405_/Y _09345_/A _09345_/Y vssd1 vssd1 vccd1 vccd1 _09411_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_111_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07599_ _07599_/A vssd1 vssd1 vccd1 vccd1 _14084_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09338_ _09345_/A _09345_/B _09345_/C vssd1 vssd1 vccd1 vccd1 _09338_/X sky130_fd_sc_hd__and3_1
XFILLER_51_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ _09187_/X _09189_/X _09049_/A _09188_/X vssd1 vssd1 vccd1 vccd1 _09271_/B
+ sky130_fd_sc_hd__a211oi_2
X_11300_ _11300_/A _11300_/B vssd1 vssd1 vccd1 vccd1 _11317_/A sky130_fd_sc_hd__xnor2_1
X_12280_ _12286_/A vssd1 vssd1 vccd1 vccd1 _12285_/A sky130_fd_sc_hd__buf_2
XFILLER_107_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11231_ _13902_/Q vssd1 vssd1 vccd1 vccd1 _11285_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12135__A input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11162_ _13920_/Q _13921_/Q _13922_/Q _13923_/Q _10679_/A _10721_/C vssd1 vssd1 vccd1
+ vccd1 _11181_/B sky130_fd_sc_hd__mux4_1
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _10064_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10114_/B sky130_fd_sc_hd__and2b_1
X_11093_ _11093_/A _11093_/B vssd1 vssd1 vccd1 vccd1 _11093_/Y sky130_fd_sc_hd__nand2_1
XFILLER_96_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input32_A dout1[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _10045_/A _10122_/A vssd1 vssd1 vccd1 vccd1 _10044_/X sky130_fd_sc_hd__and2_1
XANTENNA__14356__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13803_ _14348_/CLK _13803_/D vssd1 vssd1 vccd1 vccd1 _13803_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13643__A0 _13084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12446__A1 _08946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11995_ _13113_/B _12211_/A input65/X vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__or3b_4
XFILLER_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13734_ _13734_/A vssd1 vssd1 vccd1 vccd1 _14463_/D sky130_fd_sc_hd__clkbuf_1
X_10946_ _10946_/A _10946_/B _13894_/Q vssd1 vssd1 vccd1 vccd1 _10946_/X sky130_fd_sc_hd__or3_1
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13665_ _13678_/A _13665_/B vssd1 vssd1 vccd1 vccd1 _13666_/A sky130_fd_sc_hd__and2_1
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10877_ _13934_/Q _10875_/X _10897_/S vssd1 vssd1 vccd1 vccd1 _10878_/A sky130_fd_sc_hd__mux2_1
X_12616_ _12616_/A vssd1 vssd1 vccd1 vccd1 _14037_/D sky130_fd_sc_hd__clkbuf_1
X_13596_ _13614_/A vssd1 vssd1 vccd1 vccd1 _13611_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12547_ _12930_/A _08317_/A _12555_/S vssd1 vssd1 vccd1 vccd1 _12548_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11868__B _11870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ _14033_/Q _12464_/X _12477_/X _12473_/X vssd1 vssd1 vccd1 vccd1 _12478_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08523__A _08828_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14217_ _14217_/CLK _14217_/D _13013_/Y vssd1 vssd1 vccd1 vccd1 _14217_/Q sky130_fd_sc_hd__dfrtp_1
X_11429_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11493_/A sky130_fd_sc_hd__nor2_1
XFILLER_99_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14148_ _14164_/CLK _14148_/D vssd1 vssd1 vccd1 vccd1 _14148_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09057__C _09218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06970_ _06970_/A vssd1 vssd1 vccd1 vccd1 _06970_/X sky130_fd_sc_hd__clkbuf_2
X_14079_ _14283_/CLK _14079_/D _12724_/Y vssd1 vssd1 vccd1 vccd1 _14079_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12685__A1 _14054_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14469__181 vssd1 vssd1 vccd1 vccd1 _14469__181/HI io_oeb[1] sky130_fd_sc_hd__conb_1
XFILLER_6_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08640_ _08639_/A _08639_/C _08639_/B vssd1 vssd1 vccd1 vccd1 _08641_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09550__B2 _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08571_ _08571_/A _08944_/D vssd1 vssd1 vccd1 vccd1 _08576_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13634__A0 input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _14186_/Q _07519_/X _07541_/B _07521_/X vssd1 vssd1 vccd1 vccd1 _14178_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07453_ _14199_/Q _14201_/Q _07469_/S vssd1 vssd1 vccd1 vccd1 _07454_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07959__D _09842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07384_ _07376_/X _07382_/X _07383_/X _07379_/X vssd1 vssd1 vccd1 vccd1 _07384_/X
+ sky130_fd_sc_hd__a22o_1
X_09123_ _09457_/A _09457_/B _09123_/C _09803_/A vssd1 vssd1 vccd1 vccd1 _09127_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_109_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09054_ _09054_/A _09054_/B vssd1 vssd1 vccd1 vccd1 _09056_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08433__A _08791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14229__CLK _14256_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08005_ _08005_/A _08053_/A vssd1 vssd1 vccd1 vccd1 _08054_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11176__A1 _10722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11176__B2 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09956_ _09956_/A _09957_/A vssd1 vssd1 vccd1 vccd1 _09997_/B sky130_fd_sc_hd__xnor2_2
XFILLER_104_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08907_ _08872_/A _08872_/C _08872_/B vssd1 vssd1 vccd1 vccd1 _08908_/B sky130_fd_sc_hd__a21oi_1
XFILLER_83_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09887_ _09887_/A _09887_/B vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__xnor2_4
XFILLER_100_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08344__A2 _09848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ _08848_/A _08848_/B vssd1 vssd1 vccd1 vccd1 _08839_/B sky130_fd_sc_hd__or2b_1
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07552__A0 _14105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08769_ _08774_/B _08769_/B vssd1 vssd1 vccd1 vccd1 _08770_/B sky130_fd_sc_hd__xnor2_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12829__S _12853_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10800_ _13934_/Q _10800_/B vssd1 vssd1 vccd1 vccd1 _10801_/B sky130_fd_sc_hd__nor2_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _12193_/A input59/X _12762_/B vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10731_ _11220_/A _10746_/A _10731_/S vssd1 vssd1 vccd1 vccd1 _10812_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ _13450_/A vssd1 vssd1 vccd1 vccd1 _14381_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10662_ _10662_/A vssd1 vssd1 vccd1 vccd1 _10777_/B sky130_fd_sc_hd__buf_2
XFILLER_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12401_ _12403_/A vssd1 vssd1 vccd1 vccd1 _12401_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13381_ _13381_/A vssd1 vssd1 vccd1 vccd1 _14361_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12600__A1 _14033_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ _10622_/A _10593_/B vssd1 vssd1 vccd1 vccd1 _10593_/Y sky130_fd_sc_hd__nor2_1
X_12332_ _12335_/A vssd1 vssd1 vccd1 vccd1 _12332_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10611__B1 _09788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12263_ _12267_/A vssd1 vssd1 vccd1 vccd1 _12263_/Y sky130_fd_sc_hd__inv_2
X_14002_ _14396_/CLK _14002_/D vssd1 vssd1 vccd1 vccd1 _14002_/Q sky130_fd_sc_hd__dfxtp_1
X_11214_ _11214_/A _11300_/B vssd1 vssd1 vccd1 vccd1 _11315_/B sky130_fd_sc_hd__or2_1
X_12194_ _12213_/A _12900_/A vssd1 vssd1 vccd1 vccd1 _12201_/A sky130_fd_sc_hd__nor2_1
X_11145_ _13915_/Q _13916_/Q _13917_/Q _13918_/Q _10679_/A _10721_/C vssd1 vssd1 vccd1
+ vccd1 _11145_/X sky130_fd_sc_hd__mux4_1
XFILLER_68_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11076_ _11076_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11077_/B sky130_fd_sc_hd__or2_1
XFILLER_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10027_ _10028_/B _10027_/B vssd1 vssd1 vccd1 vccd1 _10244_/B sky130_fd_sc_hd__xnor2_2
XFILLER_62_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11875__C1 _11874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11978_ _12252_/A vssd1 vssd1 vccd1 vccd1 _12233_/A sky130_fd_sc_hd__buf_6
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10929_ _10929_/A vssd1 vssd1 vccd1 vccd1 _10993_/A sky130_fd_sc_hd__inv_2
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13717_ _13717_/A vssd1 vssd1 vccd1 vccd1 _14458_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13648_ _13661_/A _13648_/B vssd1 vssd1 vccd1 vccd1 _13649_/A sky130_fd_sc_hd__and2_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13579_ _13614_/A vssd1 vssd1 vccd1 vccd1 _13593_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09349__A _09349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09810_ _13867_/Q _13866_/Q vssd1 vssd1 vccd1 vccd1 _09875_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08574__A2 _08824_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _09741_/A _09741_/B vssd1 vssd1 vccd1 vccd1 _09741_/X sky130_fd_sc_hd__and2_1
X_06953_ _06953_/A vssd1 vssd1 vccd1 vccd1 _14316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11119__A _11119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _09712_/A _09673_/B vssd1 vssd1 vccd1 vccd1 _09672_/X sky130_fd_sc_hd__or2_1
X_06884_ _14395_/Q _06855_/Y _06864_/Y _14390_/Q vssd1 vssd1 vccd1 vccd1 _06884_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08623_ _08623_/A _08623_/B _09085_/B _09941_/A vssd1 vssd1 vccd1 vccd1 _08623_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11881__A2 _11872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _09543_/A vssd1 vssd1 vccd1 vccd1 _09001_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07505_ _07505_/A vssd1 vssd1 vccd1 vccd1 _14185_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07332__A _14105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08485_ _09865_/B vssd1 vssd1 vccd1 vccd1 _09199_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_39_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ _07425_/X _07431_/X _07434_/X _07435_/X _14204_/Q vssd1 vssd1 vccd1 vccd1
+ _14204_/D sky130_fd_sc_hd__a32o_1
XANTENNA__09039__B1 _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07367_ _07349_/X _07364_/X _07366_/X _07352_/X vssd1 vssd1 vccd1 vccd1 _07367_/X
+ sky130_fd_sc_hd__a22o_1
X_09106_ _09119_/B _09106_/B _09106_/C _09106_/D vssd1 vssd1 vccd1 vccd1 _09106_/Y
+ sky130_fd_sc_hd__nor4_4
X_07298_ _14226_/Q vssd1 vssd1 vccd1 vccd1 _07298_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09037_ _09034_/X _09035_/Y _08964_/Y _08965_/X vssd1 vssd1 vccd1 vccd1 _09037_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_102_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12897__A1 _14147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09939_ _10394_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _10013_/A sky130_fd_sc_hd__xor2_2
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12950_ _12950_/A vssd1 vssd1 vccd1 vccd1 _12950_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11901_ _13815_/Q _11882_/X _11899_/X _11900_/Y _11885_/X vssd1 vssd1 vccd1 vccd1
+ _13755_/D sky130_fd_sc_hd__o221a_1
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _12924_/A _12883_/B vssd1 vssd1 vccd1 vccd1 _12881_/X sky130_fd_sc_hd__or2_1
XANTENNA__06879__A2 _06873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11832_ _14335_/Q _11808_/X _11823_/X _13794_/Q _11831_/X vssd1 vssd1 vccd1 vccd1
+ _11832_/X sky130_fd_sc_hd__a221o_2
XANTENNA__08983__D _10007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _12426_/A vssd1 vssd1 vccd1 vccd1 _12440_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12821__B2 _14148_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10765_/B vssd1 vssd1 vccd1 vccd1 _10761_/B sky130_fd_sc_hd__clkbuf_2
X_13502_ _13502_/A _13502_/B vssd1 vssd1 vccd1 vccd1 _13503_/A sky130_fd_sc_hd__and2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _13749_/Q _13748_/Q _13747_/Q vssd1 vssd1 vccd1 vccd1 _11883_/B sky130_fd_sc_hd__or3_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13433_ _13433_/A vssd1 vssd1 vccd1 vccd1 _14376_/D sky130_fd_sc_hd__clkbuf_1
X_10645_ _10645_/A _10645_/B vssd1 vssd1 vccd1 vccd1 _10645_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13364_ _13364_/A vssd1 vssd1 vccd1 vccd1 _14356_/D sky130_fd_sc_hd__clkbuf_1
X_10576_ _10576_/A _10576_/B _10576_/C vssd1 vssd1 vccd1 vccd1 _10578_/B sky130_fd_sc_hd__and3_1
XFILLER_6_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12315_ _12316_/A vssd1 vssd1 vccd1 vccd1 _12315_/Y sky130_fd_sc_hd__inv_2
X_13295_ _14372_/Q _13215_/A _13294_/X _14452_/Q vssd1 vssd1 vccd1 vccd1 _13295_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12246_ _12252_/A vssd1 vssd1 vccd1 vccd1 _12251_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12177_ input66/X _13113_/B _13359_/A _12828_/C vssd1 vssd1 vccd1 vccd1 _12179_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_3_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11128_ _11108_/A _11124_/C _11127_/X _11319_/A _11052_/A vssd1 vssd1 vccd1 vccd1
+ _13914_/D sky130_fd_sc_hd__o32ai_1
XANTENNA__07417__A _07471_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11059_ _11117_/B _11059_/B vssd1 vssd1 vccd1 vccd1 _11059_/X sky130_fd_sc_hd__and2_1
XFILLER_110_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13154__A _13178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08270_ _09712_/A _08270_/B vssd1 vssd1 vccd1 vccd1 _08271_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07221_ _07258_/S vssd1 vssd1 vccd1 vccd1 _07235_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_34_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07152_ _07259_/S vssd1 vssd1 vccd1 vccd1 _07165_/S sky130_fd_sc_hd__buf_6
XFILLER_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08795__A2 _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ _07080_/X _14299_/Q _07083_/S vssd1 vssd1 vccd1 vccd1 _07084_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10018__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09807__A _09807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12233__A _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13915_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_102_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07327__A _14106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07985_ _07985_/A _07985_/B vssd1 vssd1 vccd1 vccd1 _07994_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09724_ _09724_/A _09724_/B vssd1 vssd1 vccd1 vccd1 _10566_/B sky130_fd_sc_hd__nand2_1
X_06936_ _06934_/X _06935_/X _14382_/Q vssd1 vssd1 vccd1 vccd1 _06937_/S sky130_fd_sc_hd__o21a_1
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14417__CLK _14417_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _10576_/A _09655_/B _10592_/A _10596_/A vssd1 vssd1 vccd1 vccd1 _09662_/A
+ sky130_fd_sc_hd__or4_1
X_06867_ _14398_/Q _06864_/Y _06865_/Y _14397_/Q _06866_/X vssd1 vssd1 vccd1 vccd1
+ _06869_/C sky130_fd_sc_hd__a221o_1
XFILLER_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11854__A2 _11808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08606_ _09434_/B _08604_/X _08605_/X vssd1 vssd1 vccd1 vccd1 _08607_/B sky130_fd_sc_hd__a21bo_1
XFILLER_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _09586_/A _09586_/B _09586_/C vssd1 vssd1 vccd1 vccd1 _09586_/Y sky130_fd_sc_hd__nand3_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08537_/A _08566_/B _08537_/C vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__and3_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08468_ _09053_/A _08468_/B _08983_/C _08703_/B vssd1 vssd1 vccd1 vccd1 _08469_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07419_ _07399_/X _07416_/X _07418_/X _07408_/X _14207_/Q vssd1 vssd1 vccd1 vccd1
+ _14207_/D sky130_fd_sc_hd__a32o_1
X_08399_ _09729_/A _09729_/B _09729_/C vssd1 vssd1 vccd1 vccd1 _08399_/Y sky130_fd_sc_hd__nor3_1
XFILLER_12_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10430_ _09766_/A _10429_/Y _10430_/S vssd1 vssd1 vccd1 vccd1 _10432_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_66_io_wbs_clk clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _14441_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_10361_ _10361_/A _10361_/B vssd1 vssd1 vccd1 vccd1 _10414_/S sky130_fd_sc_hd__nor2_1
X_12100_ _12924_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12100_/X sky130_fd_sc_hd__or2_1
XFILLER_88_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13080_ _13105_/S vssd1 vssd1 vccd1 vccd1 _13096_/S sky130_fd_sc_hd__clkbuf_2
X_10292_ _10315_/B _10292_/B vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08621__A _08621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _12031_/A vssd1 vssd1 vccd1 vccd1 _13791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12143__A input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13982_ _13982_/CLK _13982_/D _12409_/Y vssd1 vssd1 vccd1 vccd1 _13982_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14097__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12933_ _12933_/A vssd1 vssd1 vccd1 vccd1 _13254_/A sky130_fd_sc_hd__buf_2
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12909_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _12864_/X sky130_fd_sc_hd__or2_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _14329_/Q _11833_/A _11797_/X _13994_/Q _11814_/X vssd1 vssd1 vccd1 vccd1
+ _11815_/X sky130_fd_sc_hd__a221o_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _14139_/Q _12776_/A _12791_/X vssd1 vssd1 vccd1 vccd1 _12795_/X sky130_fd_sc_hd__a21o_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11746_ _07146_/Y _14226_/Q _11746_/S vssd1 vssd1 vccd1 vccd1 _11746_/X sky130_fd_sc_hd__mux2_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13934__CLK _14102_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11677_ _13775_/Q vssd1 vssd1 vccd1 vccd1 _11682_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14465_ _14465_/CLK _14465_/D vssd1 vssd1 vccd1 vccd1 _14465_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12558__A0 _12938_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13416_ input73/X _14372_/Q _13425_/S vssd1 vssd1 vccd1 vccd1 _13417_/B sky130_fd_sc_hd__mux2_1
X_10628_ _10625_/X _10626_/Y _10528_/X _10627_/X vssd1 vssd1 vccd1 vccd1 _10628_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_14396_ _14396_/CLK _14396_/D vssd1 vssd1 vccd1 vccd1 _14396_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13347_ _14352_/Q _13332_/X _13346_/X _13343_/X vssd1 vssd1 vccd1 vccd1 _14352_/D
+ sky130_fd_sc_hd__o211a_1
X_10559_ _09724_/A _10558_/X _09718_/X vssd1 vssd1 vccd1 vccd1 _10561_/A sky130_fd_sc_hd__a21oi_1
XFILLER_52_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13278_ _13343_/A vssd1 vssd1 vccd1 vccd1 _13278_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12229_ _12906_/A _12205_/A _12229_/S vssd1 vssd1 vccd1 vccd1 _12230_/B sky130_fd_sc_hd__mux2_1
XFILLER_64_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08250__B _08621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__A2 _10186_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07770_ _14259_/Q _07185_/A _07769_/X vssd1 vssd1 vccd1 vccd1 _07921_/C sky130_fd_sc_hd__o21a_2
XFILLER_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09362__A _09362_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09440_ _09440_/A _09440_/B _09440_/C vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__nand3_2
XFILLER_18_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09371_ _09371_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _09373_/B sky130_fd_sc_hd__xor2_2
XFILLER_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10020__B _10191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08322_ _08322_/A _08322_/B _08322_/C vssd1 vssd1 vccd1 vccd1 _08380_/B sky130_fd_sc_hd__nand3_2
XFILLER_75_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08465__B2 _08925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10272__A1 _09962_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08253_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _09755_/B sky130_fd_sc_hd__xnor2_2
XFILLER_119_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07204_ _07258_/S vssd1 vssd1 vccd1 vccd1 _07218_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ _09055_/A vssd1 vssd1 vccd1 vccd1 _08937_/B sky130_fd_sc_hd__buf_4
X_07135_ _06973_/A _07134_/X _14375_/Q vssd1 vssd1 vccd1 vccd1 _07136_/S sky130_fd_sc_hd__o21a_1
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07066_ _07105_/A vssd1 vssd1 vccd1 vccd1 _07098_/B sky130_fd_sc_hd__buf_2
XFILLER_88_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11524__A1 _08941_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12898__A _12942_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07968_ _08004_/B _07968_/B vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06919_ _06894_/X _06918_/X _14384_/Q vssd1 vssd1 vccd1 vccd1 _06920_/S sky130_fd_sc_hd__o21a_1
X_09707_ _09704_/X _09705_/Y _09672_/X _09674_/X vssd1 vssd1 vccd1 vccd1 _09707_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11827__A2 _11808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07899_ _07899_/A vssd1 vssd1 vccd1 vccd1 _13976_/D sky130_fd_sc_hd__clkbuf_1
X_09638_ _09638_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09665_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13957__CLK _14020_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ _09586_/A _09586_/B _09586_/C vssd1 vssd1 vccd1 vccd1 _09569_/X sky130_fd_sc_hd__and3_1
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11600_ _11600_/A vssd1 vssd1 vccd1 vccd1 _13854_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _12579_/X _14027_/Q _12583_/S vssd1 vssd1 vccd1 vccd1 _12581_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11531_ _11048_/A _11513_/X _11499_/A _13895_/Q _11514_/X vssd1 vssd1 vccd1 vccd1
+ _11531_/X sky130_fd_sc_hd__o221a_1
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14250_ _14250_/CLK _14250_/D vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_2
X_11462_ _11456_/X _11458_/Y _11460_/X _11092_/A _11461_/X vssd1 vssd1 vccd1 vccd1
+ _11462_/X sky130_fd_sc_hd__o221a_1
X_13201_ _13637_/A vssd1 vssd1 vccd1 vccd1 _13201_/X sky130_fd_sc_hd__buf_4
XANTENNA__11977__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _10413_/A _10413_/B vssd1 vssd1 vccd1 vccd1 _10416_/A sky130_fd_sc_hd__xor2_1
X_14181_ _14256_/CLK _14181_/D _12968_/Y vssd1 vssd1 vccd1 vccd1 _14181_/Q sky130_fd_sc_hd__dfrtp_1
X_11393_ _11407_/B vssd1 vssd1 vccd1 vccd1 _11403_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_87_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13132_ _13134_/A vssd1 vssd1 vccd1 vccd1 _13132_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input62_A io_wbs_adr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ _10345_/A _10345_/B vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__or2_1
XFILLER_87_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13063_ _12218_/X _14241_/Q _13076_/S vssd1 vssd1 vccd1 vccd1 _13064_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09166__B _09875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10275_ _10273_/X _10275_/B vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__and2b_1
XFILLER_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11515__A1 _11056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _13787_/Q _12000_/X _12003_/X _13827_/Q vssd1 vssd1 vccd1 vccd1 _12015_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10105__B _10106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output149_A _14305_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__A2 _10061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13965_ _14031_/CLK _13965_/D _12389_/Y vssd1 vssd1 vccd1 vccd1 _13965_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12916_ _12942_/B vssd1 vssd1 vccd1 vccd1 _12926_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13896_ _13897_/CLK _13896_/D _12303_/Y vssd1 vssd1 vccd1 vccd1 _13896_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_111_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12847_ _12847_/A _12847_/B vssd1 vssd1 vccd1 vccd1 _12848_/A sky130_fd_sc_hd__and2_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08526__A _08796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12778_ _14109_/Q _12771_/X _12775_/X _12777_/X _12207_/X vssd1 vssd1 vccd1 vccd1
+ _14109_/D sky130_fd_sc_hd__o221a_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11729_ _13767_/Q _11729_/B vssd1 vssd1 vccd1 vccd1 _11729_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_31_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14448_ _14449_/CLK _14448_/D vssd1 vssd1 vccd1 vccd1 _14448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07407__C1 _07521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14379_ _14467_/CLK _14379_/D vssd1 vssd1 vccd1 vccd1 _14379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14262__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08940_ _08940_/A _08940_/B vssd1 vssd1 vccd1 vccd1 _08950_/B sky130_fd_sc_hd__nor2_1
X_08871_ _08861_/A _08861_/B _08861_/C vssd1 vssd1 vccd1 vccd1 _08872_/C sky130_fd_sc_hd__a21o_1
XFILLER_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07822_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07847_/A sky130_fd_sc_hd__inv_2
XFILLER_96_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13259__A1 _14364_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__A _12562_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06933__A1 _14286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _14064_/Q _07720_/X _07751_/X _07752_/Y vssd1 vssd1 vccd1 vccd1 _14064_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07684_ _07684_/A _07684_/B vssd1 vssd1 vccd1 vccd1 _07685_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ _09423_/A _09423_/B _09423_/C vssd1 vssd1 vccd1 vccd1 _09423_/Y sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_leaf_12_io_wbs_clk_A clkbuf_3_1_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_80_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09354_ _09354_/A _09354_/B _09354_/C vssd1 vssd1 vccd1 vccd1 _09455_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08436__A _08789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08305_ _14022_/Q vssd1 vssd1 vccd1 vccd1 _09361_/B sky130_fd_sc_hd__clkbuf_2
X_09285_ _09482_/A _10007_/A vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__nand2_1
X_08236_ _08173_/Y _08194_/X _08274_/B _08235_/X vssd1 vssd1 vccd1 vccd1 _09749_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_119_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ _08243_/A _08167_/B _08167_/C vssd1 vssd1 vccd1 vccd1 _08168_/B sky130_fd_sc_hd__and3_1
XFILLER_109_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07118_ _14435_/Q _07117_/Y _07087_/X vssd1 vssd1 vccd1 vccd1 _07118_/X sky130_fd_sc_hd__a21o_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08098_ _09459_/A vssd1 vssd1 vccd1 vccd1 _08098_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__07267__D_N _14240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07049_ _14415_/Q _07047_/Y _07048_/X vssd1 vssd1 vccd1 vccd1 _07049_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13498__A1 _14396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10206__A _10206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _10069_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10060_/X sky130_fd_sc_hd__or2_1
XFILLER_47_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06924__A1 _14287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10962_ _10769_/A _10958_/X _10959_/X _10744_/A _10961_/X vssd1 vssd1 vccd1 vccd1
+ _11039_/A sky130_fd_sc_hd__a221oi_4
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13750_ _13826_/CLK _13750_/D _11938_/Y vssd1 vssd1 vccd1 vccd1 _13750_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12701_ _12703_/A vssd1 vssd1 vccd1 vccd1 _12701_/Y sky130_fd_sc_hd__inv_2
X_13681_ _12610_/X _14448_/Q _13687_/S vssd1 vssd1 vccd1 vccd1 _13682_/B sky130_fd_sc_hd__mux2_1
X_10893_ _10893_/A vssd1 vssd1 vccd1 vccd1 _13931_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12632_ _12632_/A vssd1 vssd1 vccd1 vccd1 _14041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12563_ _13184_/A _12563_/B vssd1 vssd1 vccd1 vccd1 _12564_/A sky130_fd_sc_hd__or2_1
XFILLER_106_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _11534_/S vssd1 vssd1 vccd1 vccd1 _11514_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14302_ _14304_/CLK _14302_/D _13169_/Y vssd1 vssd1 vccd1 vccd1 _14302_/Q sky130_fd_sc_hd__dfrtp_4
X_12494_ _14037_/Q _12485_/X _12493_/X _12473_/A vssd1 vssd1 vccd1 vccd1 _12494_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14285__CLK _14365_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09929__A1 _08893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11445_ _11466_/A _11466_/B vssd1 vssd1 vccd1 vccd1 _11465_/B sky130_fd_sc_hd__nor2_1
X_14233_ _14239_/CLK _14233_/D vssd1 vssd1 vccd1 vccd1 _14233_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14164_ _14164_/CLK _14164_/D vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_2
X_11376_ hold39/A _11363_/X _11370_/X _11375_/X vssd1 vssd1 vccd1 vccd1 _13889_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13115_ _13115_/A vssd1 vssd1 vccd1 vccd1 _13115_/Y sky130_fd_sc_hd__inv_2
X_10327_ _10589_/A _10598_/C vssd1 vssd1 vccd1 vccd1 _10327_/X sky130_fd_sc_hd__or2_1
XFILLER_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14095_ _14102_/CLK _14095_/D _12744_/Y vssd1 vssd1 vccd1 vccd1 _14095_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13046_ _14234_/Q _13041_/X _13045_/X _13039_/X vssd1 vssd1 vccd1 vccd1 _14234_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10258_ _10259_/A _10259_/B vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__or2_1
XFILLER_61_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10189_ _10191_/A _10191_/B _09897_/X vssd1 vssd1 vccd1 vccd1 _10226_/A sky130_fd_sc_hd__a21oi_1
XFILLER_39_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07425__A _07452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13948_ _13949_/CLK _13948_/D _12368_/Y vssd1 vssd1 vccd1 vccd1 _13948_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_3_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13879_ _14198_/CLK _13879_/D _12282_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09093__A1 _08573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__B2 _08012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ _09119_/A _09068_/Y _08991_/B _08993_/B vssd1 vssd1 vccd1 vccd1 _09106_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_78_io_wbs_clk_A clkbuf_3_0_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_08021_ _08021_/A _08078_/C vssd1 vssd1 vccd1 vccd1 _08054_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08703__B _08703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__B2 _13828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09972_ _10151_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _10274_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08923_ _09188_/A _08918_/B _08919_/A _08954_/A vssd1 vssd1 vccd1 vccd1 _08924_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__14008__CLK _14008_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09815__A _10271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__A1 _07158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12152__A1 _13823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08854_ _08859_/A _08852_/Y _08858_/A vssd1 vssd1 vccd1 vccd1 _08856_/B sky130_fd_sc_hd__a21o_1
XFILLER_44_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07805_ _10727_/B vssd1 vssd1 vccd1 vccd1 _10705_/B sky130_fd_sc_hd__clkbuf_4
X_08785_ _08785_/A _08785_/B _08785_/C vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__nand3_1
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07736_ _07736_/A vssd1 vssd1 vccd1 vccd1 _14069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07667_ _07667_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07740_/A sky130_fd_sc_hd__xnor2_4
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10696__A _11240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13072__A _13072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09406_ _09345_/A _09345_/Y _09404_/X _09405_/Y vssd1 vssd1 vccd1 vccd1 _09411_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07598_ _14084_/Q input31/X _07604_/S vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10218__A1 _10067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09337_ _09345_/A _09345_/C _09345_/B vssd1 vssd1 vccd1 vccd1 _09337_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ _09049_/A _09188_/X _09187_/A _09189_/X vssd1 vssd1 vccd1 vccd1 _09271_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08219_ _09771_/B _08219_/B vssd1 vssd1 vccd1 vccd1 _08221_/A sky130_fd_sc_hd__xnor2_1
XFILLER_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09199_ _09472_/A _09361_/B _09866_/A _09199_/D vssd1 vssd1 vccd1 vccd1 _09202_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_14_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12416__A input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ _11288_/A _11288_/B vssd1 vssd1 vccd1 vccd1 _11327_/A sky130_fd_sc_hd__and2_1
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11161_ _10769_/A _11158_/X _11160_/X vssd1 vssd1 vccd1 vccd1 _11256_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12850__S _12853_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10112_ _10063_/B _10112_/B vssd1 vssd1 vccd1 vccd1 _10114_/A sky130_fd_sc_hd__and2b_1
XFILLER_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11092_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11093_/B sky130_fd_sc_hd__or2_1
XFILLER_103_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10043_ _10354_/B _10073_/B _10042_/X vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__a21o_1
XFILLER_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12151__A _12904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_input25_A dout1[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13802_ _13820_/CLK _13802_/D vssd1 vssd1 vccd1 vccd1 _13802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11994_ _11994_/A _12952_/B vssd1 vssd1 vccd1 vccd1 _13113_/B sky130_fd_sc_hd__or2_1
XFILLER_1_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13733_ _13745_/A _13733_/B vssd1 vssd1 vccd1 vccd1 _13734_/A sky130_fd_sc_hd__and2_1
X_10945_ _10946_/A _13895_/Q _10946_/B vssd1 vssd1 vccd1 vccd1 _10945_/X sky130_fd_sc_hd__or3b_1
XFILLER_95_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13664_ input95/X _14443_/Q _13670_/S vssd1 vssd1 vccd1 vccd1 _13665_/B sky130_fd_sc_hd__mux2_1
XFILLER_108_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10876_ _10902_/S vssd1 vssd1 vccd1 vccd1 _10897_/S sky130_fd_sc_hd__buf_2
XANTENNA__11214__B _11300_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12615_ _12615_/A _12615_/B vssd1 vssd1 vccd1 vccd1 _12616_/A sky130_fd_sc_hd__and2_1
XANTENNA__09075__A1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13595_ _13595_/A vssd1 vssd1 vccd1 vccd1 _14423_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_2_3_0_io_wbs_clk_A clkbuf_2_3_0_io_wbs_clk/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_118_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12546_ _12546_/A vssd1 vssd1 vccd1 vccd1 _14017_/D sky130_fd_sc_hd__clkbuf_1
X_12477_ _08632_/A _12465_/X _12476_/X _14049_/Q vssd1 vssd1 vccd1 vccd1 _12477_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14216_ _14224_/CLK _14216_/D _13012_/Y vssd1 vssd1 vccd1 vccd1 _14216_/Q sky130_fd_sc_hd__dfrtp_2
X_11428_ _11285_/A _11014_/B _11436_/S vssd1 vssd1 vccd1 vccd1 _11497_/B sky130_fd_sc_hd__mux2_1
XFILLER_6_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14147_ _14164_/CLK _14147_/D vssd1 vssd1 vccd1 vccd1 _14147_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_4_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11359_ _14057_/Q _13969_/Q vssd1 vssd1 vccd1 vccd1 _11536_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09057__D _09848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09635__A _09635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14078_ _14283_/CLK _14078_/D _12723_/Y vssd1 vssd1 vccd1 vccd1 _14078_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06978__B _14280_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _13116_/A vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08570_ _10081_/A vssd1 vssd1 vccd1 vccd1 _08944_/D sky130_fd_sc_hd__buf_4
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07521_ _07520_/Y _07521_/B _14178_/Q _07521_/D vssd1 vssd1 vccd1 vccd1 _07521_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07452_ _07452_/A vssd1 vssd1 vccd1 vccd1 _07452_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07383_ _14212_/Q _14214_/Q _07387_/S vssd1 vssd1 vccd1 vccd1 _07383_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09122_ _09336_/A _09192_/B vssd1 vssd1 vccd1 vccd1 _09184_/A sky130_fd_sc_hd__xor2_1
XFILLER_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09053_ _09053_/A _09053_/B _09824_/A _09857_/A vssd1 vssd1 vccd1 vccd1 _09054_/B
+ sky130_fd_sc_hd__and4_1
X_08004_ _08004_/A _08004_/B vssd1 vssd1 vccd1 vccd1 _08053_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09955_ _10003_/A _10003_/B _09954_/X vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__o21a_1
XFILLER_44_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08906_ _08906_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08915_/A sky130_fd_sc_hd__xnor2_1
XFILLER_106_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09886_ _09906_/A _09884_/X _09885_/X vssd1 vssd1 vccd1 vccd1 _10050_/B sky130_fd_sc_hd__a21oi_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10687__A1 _10686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08837_ _08844_/B _08837_/B vssd1 vssd1 vccd1 vccd1 _08848_/B sky130_fd_sc_hd__xnor2_1
XFILLER_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07552__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _08707_/A _08706_/A _08706_/B vssd1 vssd1 vccd1 vccd1 _08769_/B sky130_fd_sc_hd__o21ba_1
XFILLER_73_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07719_ _07719_/A vssd1 vssd1 vccd1 vccd1 _14072_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _08745_/B _08745_/C _08745_/A vssd1 vssd1 vccd1 vccd1 _08701_/B sky130_fd_sc_hd__a21bo_1
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10730_ _10730_/A _10730_/B vssd1 vssd1 vccd1 vccd1 _10731_/S sky130_fd_sc_hd__nand2_1
XFILLER_14_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10661_ _10954_/A vssd1 vssd1 vccd1 vccd1 _10662_/A sky130_fd_sc_hd__buf_2
XFILLER_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13530__A _13539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07068__B1 _14356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ _12403_/A vssd1 vssd1 vccd1 vccd1 _12400_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12061__B1 _12060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13380_ _13392_/A _13380_/B vssd1 vssd1 vccd1 vccd1 _13381_/A sky130_fd_sc_hd__and2_1
X_10592_ _10592_/A _10592_/B vssd1 vssd1 vccd1 vccd1 _10593_/B sky130_fd_sc_hd__xnor2_1
XFILLER_51_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10611__A1 _10634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12331_ _12335_/A vssd1 vssd1 vccd1 vccd1 _12331_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12146__A _12146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12262_ _12286_/A vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__buf_2
X_11213_ _11213_/A _11213_/B vssd1 vssd1 vccd1 vccd1 _11300_/B sky130_fd_sc_hd__xnor2_2
X_14001_ _14396_/CLK _14001_/D vssd1 vssd1 vccd1 vccd1 _14001_/Q sky130_fd_sc_hd__dfxtp_1
X_12193_ _12193_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12213_/A sky130_fd_sc_hd__nand2_1
X_11144_ _10652_/X _11141_/X _11143_/X vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11075_ _11104_/B _11108_/B _11104_/A vssd1 vssd1 vccd1 vccd1 _11105_/B sky130_fd_sc_hd__o21a_1
XFILLER_62_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10026_ _10111_/A _10024_/X _10025_/X vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11977_ _12223_/A vssd1 vssd1 vccd1 vccd1 _12252_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_91_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13716_ _13729_/A _13716_/B vssd1 vssd1 vccd1 vccd1 _13717_/A sky130_fd_sc_hd__and2_1
X_10928_ _11142_/A _10927_/Y _10920_/X vssd1 vssd1 vccd1 vccd1 _10929_/A sky130_fd_sc_hd__a21boi_1
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13647_ input88/X _14438_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13648_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10859_ _13979_/Q _10906_/A vssd1 vssd1 vccd1 vccd1 _10859_/Y sky130_fd_sc_hd__nand2_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13578_ _13578_/A vssd1 vssd1 vccd1 vccd1 _14418_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12529_ _12529_/A vssd1 vssd1 vccd1 vccd1 _14012_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09349__B _09821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13552__A0 input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_io_wbs_clk clkbuf_3_2_0_io_wbs_clk/X vssd1 vssd1 vccd1 vccd1 _13982_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold33_A hold33/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06952_ _06948_/X _14316_/Q _06952_/S vssd1 vssd1 vccd1 vccd1 _06953_/A sky130_fd_sc_hd__mux2_1
X_09740_ _09742_/A _10540_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09741_/B sky130_fd_sc_hd__o21bai_2
XANTENNA__10304__A _10333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

