VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO merge_memory
  CLASS BLOCK ;
  FOREIGN merge_memory ;
  ORIGIN 0.000 0.000 ;
  SIZE 750.000 BY 200.000 ;
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 17.720 750.000 18.320 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 21.800 750.000 22.400 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 25.880 750.000 26.480 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 29.960 750.000 30.560 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 34.040 750.000 34.640 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 38.120 750.000 38.720 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 42.200 750.000 42.800 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 46.280 750.000 46.880 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 50.360 750.000 50.960 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 54.440 750.000 55.040 ;
    END
  END addr[9]
  PIN addr_mem0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END addr_mem0[0]
  PIN addr_mem0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END addr_mem0[1]
  PIN addr_mem0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END addr_mem0[2]
  PIN addr_mem0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END addr_mem0[3]
  PIN addr_mem0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END addr_mem0[4]
  PIN addr_mem0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END addr_mem0[5]
  PIN addr_mem0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END addr_mem0[6]
  PIN addr_mem0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END addr_mem0[7]
  PIN addr_mem0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END addr_mem0[8]
  PIN addr_mem1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END addr_mem1[0]
  PIN addr_mem1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END addr_mem1[1]
  PIN addr_mem1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END addr_mem1[2]
  PIN addr_mem1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END addr_mem1[3]
  PIN addr_mem1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END addr_mem1[4]
  PIN addr_mem1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END addr_mem1[5]
  PIN addr_mem1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END addr_mem1[6]
  PIN addr_mem1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END addr_mem1[7]
  PIN addr_mem1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END addr_mem1[8]
  PIN csb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 13.640 750.000 14.240 ;
    END
  END csb
  PIN csb_mem0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END csb_mem0
  PIN csb_mem1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END csb_mem1
  PIN dout[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 58.520 750.000 59.120 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 99.320 750.000 99.920 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 103.400 750.000 104.000 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 107.480 750.000 108.080 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 111.560 750.000 112.160 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 115.640 750.000 116.240 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 119.720 750.000 120.320 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 123.800 750.000 124.400 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 127.880 750.000 128.480 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 131.960 750.000 132.560 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 136.040 750.000 136.640 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 62.600 750.000 63.200 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 140.120 750.000 140.720 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 144.200 750.000 144.800 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 148.280 750.000 148.880 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 152.360 750.000 152.960 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 156.440 750.000 157.040 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 160.520 750.000 161.120 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 164.600 750.000 165.200 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 168.680 750.000 169.280 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 172.760 750.000 173.360 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 176.840 750.000 177.440 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 66.680 750.000 67.280 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 180.920 750.000 181.520 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 185.000 750.000 185.600 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 70.760 750.000 71.360 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 74.840 750.000 75.440 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 78.920 750.000 79.520 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 83.000 750.000 83.600 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 87.080 750.000 87.680 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 91.160 750.000 91.760 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 746.000 95.240 750.000 95.840 ;
    END
  END dout[9]
  PIN dout_mem0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END dout_mem0[0]
  PIN dout_mem0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END dout_mem0[10]
  PIN dout_mem0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END dout_mem0[11]
  PIN dout_mem0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END dout_mem0[12]
  PIN dout_mem0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END dout_mem0[13]
  PIN dout_mem0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END dout_mem0[14]
  PIN dout_mem0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END dout_mem0[15]
  PIN dout_mem0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END dout_mem0[16]
  PIN dout_mem0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END dout_mem0[17]
  PIN dout_mem0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END dout_mem0[18]
  PIN dout_mem0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END dout_mem0[19]
  PIN dout_mem0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END dout_mem0[1]
  PIN dout_mem0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END dout_mem0[20]
  PIN dout_mem0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END dout_mem0[21]
  PIN dout_mem0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END dout_mem0[22]
  PIN dout_mem0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END dout_mem0[23]
  PIN dout_mem0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END dout_mem0[24]
  PIN dout_mem0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END dout_mem0[25]
  PIN dout_mem0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END dout_mem0[26]
  PIN dout_mem0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END dout_mem0[27]
  PIN dout_mem0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END dout_mem0[28]
  PIN dout_mem0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END dout_mem0[29]
  PIN dout_mem0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END dout_mem0[2]
  PIN dout_mem0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 4.000 ;
    END
  END dout_mem0[30]
  PIN dout_mem0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END dout_mem0[31]
  PIN dout_mem0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END dout_mem0[3]
  PIN dout_mem0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END dout_mem0[4]
  PIN dout_mem0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END dout_mem0[5]
  PIN dout_mem0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END dout_mem0[6]
  PIN dout_mem0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END dout_mem0[7]
  PIN dout_mem0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END dout_mem0[8]
  PIN dout_mem0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END dout_mem0[9]
  PIN dout_mem1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END dout_mem1[0]
  PIN dout_mem1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END dout_mem1[10]
  PIN dout_mem1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END dout_mem1[11]
  PIN dout_mem1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END dout_mem1[12]
  PIN dout_mem1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END dout_mem1[13]
  PIN dout_mem1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END dout_mem1[14]
  PIN dout_mem1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 4.000 ;
    END
  END dout_mem1[15]
  PIN dout_mem1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END dout_mem1[16]
  PIN dout_mem1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END dout_mem1[17]
  PIN dout_mem1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END dout_mem1[18]
  PIN dout_mem1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END dout_mem1[19]
  PIN dout_mem1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END dout_mem1[1]
  PIN dout_mem1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END dout_mem1[20]
  PIN dout_mem1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END dout_mem1[21]
  PIN dout_mem1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END dout_mem1[22]
  PIN dout_mem1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END dout_mem1[23]
  PIN dout_mem1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END dout_mem1[24]
  PIN dout_mem1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 0.000 685.310 4.000 ;
    END
  END dout_mem1[25]
  PIN dout_mem1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 4.000 ;
    END
  END dout_mem1[26]
  PIN dout_mem1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END dout_mem1[27]
  PIN dout_mem1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END dout_mem1[28]
  PIN dout_mem1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 0.000 720.270 4.000 ;
    END
  END dout_mem1[29]
  PIN dout_mem1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END dout_mem1[2]
  PIN dout_mem1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 0.000 729.010 4.000 ;
    END
  END dout_mem1[30]
  PIN dout_mem1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END dout_mem1[31]
  PIN dout_mem1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END dout_mem1[3]
  PIN dout_mem1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END dout_mem1[4]
  PIN dout_mem1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 0.000 510.510 4.000 ;
    END
  END dout_mem1[5]
  PIN dout_mem1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END dout_mem1[6]
  PIN dout_mem1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END dout_mem1[7]
  PIN dout_mem1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END dout_mem1[8]
  PIN dout_mem1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END dout_mem1[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 187.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 187.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 187.920 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 186.265 744.470 187.870 ;
        RECT 5.330 180.825 744.470 183.655 ;
        RECT 5.330 175.385 744.470 178.215 ;
        RECT 5.330 169.945 744.470 172.775 ;
        RECT 5.330 164.505 744.470 167.335 ;
        RECT 5.330 159.065 744.470 161.895 ;
        RECT 5.330 153.625 744.470 156.455 ;
        RECT 5.330 148.185 744.470 151.015 ;
        RECT 5.330 142.745 744.470 145.575 ;
        RECT 5.330 137.305 744.470 140.135 ;
        RECT 5.330 131.865 744.470 134.695 ;
        RECT 5.330 126.425 744.470 129.255 ;
        RECT 5.330 120.985 744.470 123.815 ;
        RECT 5.330 115.545 744.470 118.375 ;
        RECT 5.330 110.105 744.470 112.935 ;
        RECT 5.330 104.665 744.470 107.495 ;
        RECT 5.330 99.225 744.470 102.055 ;
        RECT 5.330 93.785 744.470 96.615 ;
        RECT 5.330 88.345 744.470 91.175 ;
        RECT 5.330 82.905 744.470 85.735 ;
        RECT 5.330 77.465 744.470 80.295 ;
        RECT 5.330 72.025 744.470 74.855 ;
        RECT 5.330 66.585 744.470 69.415 ;
        RECT 5.330 61.145 744.470 63.975 ;
        RECT 5.330 55.705 744.470 58.535 ;
        RECT 5.330 50.265 744.470 53.095 ;
        RECT 5.330 44.825 744.470 47.655 ;
        RECT 5.330 39.385 744.470 42.215 ;
        RECT 5.330 33.945 744.470 36.775 ;
        RECT 5.330 28.505 744.470 31.335 ;
        RECT 5.330 23.065 744.470 25.895 ;
        RECT 5.330 17.625 744.470 20.455 ;
        RECT 5.330 12.185 744.470 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 744.280 187.765 ;
      LAYER met1 ;
        RECT 5.520 2.420 744.280 187.920 ;
      LAYER met2 ;
        RECT 12.060 4.280 740.970 187.865 ;
        RECT 12.610 2.390 20.510 4.280 ;
        RECT 21.350 2.390 29.250 4.280 ;
        RECT 30.090 2.390 37.990 4.280 ;
        RECT 38.830 2.390 46.730 4.280 ;
        RECT 47.570 2.390 55.470 4.280 ;
        RECT 56.310 2.390 64.210 4.280 ;
        RECT 65.050 2.390 72.950 4.280 ;
        RECT 73.790 2.390 81.690 4.280 ;
        RECT 82.530 2.390 90.430 4.280 ;
        RECT 91.270 2.390 99.170 4.280 ;
        RECT 100.010 2.390 107.910 4.280 ;
        RECT 108.750 2.390 116.650 4.280 ;
        RECT 117.490 2.390 125.390 4.280 ;
        RECT 126.230 2.390 134.130 4.280 ;
        RECT 134.970 2.390 142.870 4.280 ;
        RECT 143.710 2.390 151.610 4.280 ;
        RECT 152.450 2.390 160.350 4.280 ;
        RECT 161.190 2.390 169.090 4.280 ;
        RECT 169.930 2.390 177.830 4.280 ;
        RECT 178.670 2.390 186.570 4.280 ;
        RECT 187.410 2.390 195.310 4.280 ;
        RECT 196.150 2.390 204.050 4.280 ;
        RECT 204.890 2.390 212.790 4.280 ;
        RECT 213.630 2.390 221.530 4.280 ;
        RECT 222.370 2.390 230.270 4.280 ;
        RECT 231.110 2.390 239.010 4.280 ;
        RECT 239.850 2.390 247.750 4.280 ;
        RECT 248.590 2.390 256.490 4.280 ;
        RECT 257.330 2.390 265.230 4.280 ;
        RECT 266.070 2.390 273.970 4.280 ;
        RECT 274.810 2.390 282.710 4.280 ;
        RECT 283.550 2.390 291.450 4.280 ;
        RECT 292.290 2.390 300.190 4.280 ;
        RECT 301.030 2.390 308.930 4.280 ;
        RECT 309.770 2.390 317.670 4.280 ;
        RECT 318.510 2.390 326.410 4.280 ;
        RECT 327.250 2.390 335.150 4.280 ;
        RECT 335.990 2.390 343.890 4.280 ;
        RECT 344.730 2.390 352.630 4.280 ;
        RECT 353.470 2.390 361.370 4.280 ;
        RECT 362.210 2.390 370.110 4.280 ;
        RECT 370.950 2.390 378.850 4.280 ;
        RECT 379.690 2.390 387.590 4.280 ;
        RECT 388.430 2.390 396.330 4.280 ;
        RECT 397.170 2.390 405.070 4.280 ;
        RECT 405.910 2.390 413.810 4.280 ;
        RECT 414.650 2.390 422.550 4.280 ;
        RECT 423.390 2.390 431.290 4.280 ;
        RECT 432.130 2.390 440.030 4.280 ;
        RECT 440.870 2.390 448.770 4.280 ;
        RECT 449.610 2.390 457.510 4.280 ;
        RECT 458.350 2.390 466.250 4.280 ;
        RECT 467.090 2.390 474.990 4.280 ;
        RECT 475.830 2.390 483.730 4.280 ;
        RECT 484.570 2.390 492.470 4.280 ;
        RECT 493.310 2.390 501.210 4.280 ;
        RECT 502.050 2.390 509.950 4.280 ;
        RECT 510.790 2.390 518.690 4.280 ;
        RECT 519.530 2.390 527.430 4.280 ;
        RECT 528.270 2.390 536.170 4.280 ;
        RECT 537.010 2.390 544.910 4.280 ;
        RECT 545.750 2.390 553.650 4.280 ;
        RECT 554.490 2.390 562.390 4.280 ;
        RECT 563.230 2.390 571.130 4.280 ;
        RECT 571.970 2.390 579.870 4.280 ;
        RECT 580.710 2.390 588.610 4.280 ;
        RECT 589.450 2.390 597.350 4.280 ;
        RECT 598.190 2.390 606.090 4.280 ;
        RECT 606.930 2.390 614.830 4.280 ;
        RECT 615.670 2.390 623.570 4.280 ;
        RECT 624.410 2.390 632.310 4.280 ;
        RECT 633.150 2.390 641.050 4.280 ;
        RECT 641.890 2.390 649.790 4.280 ;
        RECT 650.630 2.390 658.530 4.280 ;
        RECT 659.370 2.390 667.270 4.280 ;
        RECT 668.110 2.390 676.010 4.280 ;
        RECT 676.850 2.390 684.750 4.280 ;
        RECT 685.590 2.390 693.490 4.280 ;
        RECT 694.330 2.390 702.230 4.280 ;
        RECT 703.070 2.390 710.970 4.280 ;
        RECT 711.810 2.390 719.710 4.280 ;
        RECT 720.550 2.390 728.450 4.280 ;
        RECT 729.290 2.390 737.190 4.280 ;
        RECT 738.030 2.390 740.970 4.280 ;
      LAYER met3 ;
        RECT 21.050 186.000 746.000 187.845 ;
        RECT 21.050 184.600 745.600 186.000 ;
        RECT 21.050 181.920 746.000 184.600 ;
        RECT 21.050 180.520 745.600 181.920 ;
        RECT 21.050 177.840 746.000 180.520 ;
        RECT 21.050 176.440 745.600 177.840 ;
        RECT 21.050 173.760 746.000 176.440 ;
        RECT 21.050 172.360 745.600 173.760 ;
        RECT 21.050 169.680 746.000 172.360 ;
        RECT 21.050 168.280 745.600 169.680 ;
        RECT 21.050 165.600 746.000 168.280 ;
        RECT 21.050 164.200 745.600 165.600 ;
        RECT 21.050 161.520 746.000 164.200 ;
        RECT 21.050 160.120 745.600 161.520 ;
        RECT 21.050 157.440 746.000 160.120 ;
        RECT 21.050 156.040 745.600 157.440 ;
        RECT 21.050 153.360 746.000 156.040 ;
        RECT 21.050 151.960 745.600 153.360 ;
        RECT 21.050 149.280 746.000 151.960 ;
        RECT 21.050 147.880 745.600 149.280 ;
        RECT 21.050 145.200 746.000 147.880 ;
        RECT 21.050 143.800 745.600 145.200 ;
        RECT 21.050 141.120 746.000 143.800 ;
        RECT 21.050 139.720 745.600 141.120 ;
        RECT 21.050 137.040 746.000 139.720 ;
        RECT 21.050 135.640 745.600 137.040 ;
        RECT 21.050 132.960 746.000 135.640 ;
        RECT 21.050 131.560 745.600 132.960 ;
        RECT 21.050 128.880 746.000 131.560 ;
        RECT 21.050 127.480 745.600 128.880 ;
        RECT 21.050 124.800 746.000 127.480 ;
        RECT 21.050 123.400 745.600 124.800 ;
        RECT 21.050 120.720 746.000 123.400 ;
        RECT 21.050 119.320 745.600 120.720 ;
        RECT 21.050 116.640 746.000 119.320 ;
        RECT 21.050 115.240 745.600 116.640 ;
        RECT 21.050 112.560 746.000 115.240 ;
        RECT 21.050 111.160 745.600 112.560 ;
        RECT 21.050 108.480 746.000 111.160 ;
        RECT 21.050 107.080 745.600 108.480 ;
        RECT 21.050 104.400 746.000 107.080 ;
        RECT 21.050 103.000 745.600 104.400 ;
        RECT 21.050 100.320 746.000 103.000 ;
        RECT 21.050 98.920 745.600 100.320 ;
        RECT 21.050 96.240 746.000 98.920 ;
        RECT 21.050 94.840 745.600 96.240 ;
        RECT 21.050 92.160 746.000 94.840 ;
        RECT 21.050 90.760 745.600 92.160 ;
        RECT 21.050 88.080 746.000 90.760 ;
        RECT 21.050 86.680 745.600 88.080 ;
        RECT 21.050 84.000 746.000 86.680 ;
        RECT 21.050 82.600 745.600 84.000 ;
        RECT 21.050 79.920 746.000 82.600 ;
        RECT 21.050 78.520 745.600 79.920 ;
        RECT 21.050 75.840 746.000 78.520 ;
        RECT 21.050 74.440 745.600 75.840 ;
        RECT 21.050 71.760 746.000 74.440 ;
        RECT 21.050 70.360 745.600 71.760 ;
        RECT 21.050 67.680 746.000 70.360 ;
        RECT 21.050 66.280 745.600 67.680 ;
        RECT 21.050 63.600 746.000 66.280 ;
        RECT 21.050 62.200 745.600 63.600 ;
        RECT 21.050 59.520 746.000 62.200 ;
        RECT 21.050 58.120 745.600 59.520 ;
        RECT 21.050 55.440 746.000 58.120 ;
        RECT 21.050 54.040 745.600 55.440 ;
        RECT 21.050 51.360 746.000 54.040 ;
        RECT 21.050 49.960 745.600 51.360 ;
        RECT 21.050 47.280 746.000 49.960 ;
        RECT 21.050 45.880 745.600 47.280 ;
        RECT 21.050 43.200 746.000 45.880 ;
        RECT 21.050 41.800 745.600 43.200 ;
        RECT 21.050 39.120 746.000 41.800 ;
        RECT 21.050 37.720 745.600 39.120 ;
        RECT 21.050 35.040 746.000 37.720 ;
        RECT 21.050 33.640 745.600 35.040 ;
        RECT 21.050 30.960 746.000 33.640 ;
        RECT 21.050 29.560 745.600 30.960 ;
        RECT 21.050 26.880 746.000 29.560 ;
        RECT 21.050 25.480 745.600 26.880 ;
        RECT 21.050 22.800 746.000 25.480 ;
        RECT 21.050 21.400 745.600 22.800 ;
        RECT 21.050 18.720 746.000 21.400 ;
        RECT 21.050 17.320 745.600 18.720 ;
        RECT 21.050 14.640 746.000 17.320 ;
        RECT 21.050 13.240 745.600 14.640 ;
        RECT 21.050 4.255 746.000 13.240 ;
  END
END merge_memory
END LIBRARY

