magic
tech sky130A
magscale 1 2
timestamp 1657783833
<< viali >>
rect 1685 75293 1719 75327
rect 2145 75293 2179 75327
rect 77861 75293 77895 75327
rect 1501 75157 1535 75191
rect 77309 75157 77343 75191
rect 78045 75157 78079 75191
rect 1409 74817 1443 74851
rect 77861 74817 77895 74851
rect 77677 74681 77711 74715
rect 1593 74613 1627 74647
rect 1409 74341 1443 74375
rect 78137 74341 78171 74375
rect 1685 73729 1719 73763
rect 77677 73729 77711 73763
rect 1501 73593 1535 73627
rect 77861 73593 77895 73627
rect 2237 73525 2271 73559
rect 77125 73525 77159 73559
rect 1685 73117 1719 73151
rect 77861 73117 77895 73151
rect 1501 72981 1535 73015
rect 2237 72981 2271 73015
rect 78045 72981 78079 73015
rect 1685 72641 1719 72675
rect 77677 72641 77711 72675
rect 1501 72437 1535 72471
rect 2237 72437 2271 72471
rect 77861 72437 77895 72471
rect 1685 72029 1719 72063
rect 77861 72029 77895 72063
rect 1501 71893 1535 71927
rect 2237 71893 2271 71927
rect 78045 71893 78079 71927
rect 76205 71689 76239 71723
rect 72617 71553 72651 71587
rect 73445 71553 73479 71587
rect 76021 71553 76055 71587
rect 72433 71349 72467 71383
rect 76665 71349 76699 71383
rect 76113 71145 76147 71179
rect 1685 70941 1719 70975
rect 72065 70941 72099 70975
rect 72617 70941 72651 70975
rect 75929 70941 75963 70975
rect 76573 70941 76607 70975
rect 77861 70941 77895 70975
rect 1501 70805 1535 70839
rect 2237 70805 2271 70839
rect 71881 70805 71915 70839
rect 78045 70805 78079 70839
rect 71237 70601 71271 70635
rect 74825 70601 74859 70635
rect 1685 70465 1719 70499
rect 71421 70465 71455 70499
rect 71973 70465 72007 70499
rect 74641 70465 74675 70499
rect 75285 70465 75319 70499
rect 77677 70465 77711 70499
rect 2237 70397 2271 70431
rect 1501 70261 1535 70295
rect 77861 70261 77895 70295
rect 74089 70057 74123 70091
rect 1409 69853 1443 69887
rect 2145 69853 2179 69887
rect 71053 69853 71087 69887
rect 71605 69853 71639 69887
rect 73905 69853 73939 69887
rect 77493 69853 77527 69887
rect 78137 69853 78171 69887
rect 1593 69717 1627 69751
rect 70869 69717 70903 69751
rect 74549 69717 74583 69751
rect 77953 69717 77987 69751
rect 1409 69377 1443 69411
rect 2145 69377 2179 69411
rect 77309 69377 77343 69411
rect 77953 69377 77987 69411
rect 1593 69173 1627 69207
rect 77769 69173 77803 69207
rect 73353 68969 73387 69003
rect 70133 68765 70167 68799
rect 70869 68765 70903 68799
rect 73169 68765 73203 68799
rect 1409 68629 1443 68663
rect 69949 68629 69983 68663
rect 73813 68629 73847 68663
rect 78045 68629 78079 68663
rect 1409 68289 1443 68323
rect 77953 68289 77987 68323
rect 1593 68085 1627 68119
rect 77769 68085 77803 68119
rect 1593 67813 1627 67847
rect 77953 67813 77987 67847
rect 1409 67677 1443 67711
rect 2145 67677 2179 67711
rect 77493 67677 77527 67711
rect 78137 67677 78171 67711
rect 1409 67201 1443 67235
rect 2145 67201 2179 67235
rect 77309 67201 77343 67235
rect 77953 67201 77987 67235
rect 77769 67065 77803 67099
rect 1593 66997 1627 67031
rect 1409 66589 1443 66623
rect 2145 66589 2179 66623
rect 77493 66589 77527 66623
rect 78137 66589 78171 66623
rect 1593 66453 1627 66487
rect 77953 66453 77987 66487
rect 1409 65909 1443 65943
rect 1409 65501 1443 65535
rect 77493 65501 77527 65535
rect 78137 65501 78171 65535
rect 1593 65365 1627 65399
rect 77953 65365 77987 65399
rect 1593 65161 1627 65195
rect 1409 65025 1443 65059
rect 2145 65025 2179 65059
rect 77309 65025 77343 65059
rect 77953 65025 77987 65059
rect 77769 64889 77803 64923
rect 1409 64413 1443 64447
rect 2145 64413 2179 64447
rect 77493 64413 77527 64447
rect 78137 64413 78171 64447
rect 1593 64277 1627 64311
rect 77953 64277 77987 64311
rect 1409 63937 1443 63971
rect 2145 63937 2179 63971
rect 77309 63937 77343 63971
rect 77953 63937 77987 63971
rect 77769 63801 77803 63835
rect 1593 63733 1627 63767
rect 1409 63189 1443 63223
rect 78045 63189 78079 63223
rect 1409 62849 1443 62883
rect 77953 62849 77987 62883
rect 1593 62645 1627 62679
rect 77769 62645 77803 62679
rect 65717 62441 65751 62475
rect 1409 62237 1443 62271
rect 2145 62237 2179 62271
rect 77493 62237 77527 62271
rect 78137 62237 78171 62271
rect 1593 62101 1627 62135
rect 64245 62101 64279 62135
rect 77953 62101 77987 62135
rect 64521 61897 64555 61931
rect 66177 61897 66211 61931
rect 65717 61829 65751 61863
rect 1409 61761 1443 61795
rect 2145 61761 2179 61795
rect 64061 61761 64095 61795
rect 77309 61761 77343 61795
rect 77953 61761 77987 61795
rect 65073 61625 65107 61659
rect 1593 61557 1627 61591
rect 63877 61557 63911 61591
rect 66729 61557 66763 61591
rect 77769 61557 77803 61591
rect 63141 61353 63175 61387
rect 64981 61285 65015 61319
rect 66177 61285 66211 61319
rect 1409 61149 1443 61183
rect 2145 61149 2179 61183
rect 63969 61149 64003 61183
rect 64429 61149 64463 61183
rect 64849 61149 64883 61183
rect 65625 61149 65659 61183
rect 65998 61149 66032 61183
rect 66729 61149 66763 61183
rect 67465 61149 67499 61183
rect 77493 61149 77527 61183
rect 78137 61149 78171 61183
rect 64613 61081 64647 61115
rect 64705 61081 64739 61115
rect 65809 61081 65843 61115
rect 65901 61081 65935 61115
rect 1593 61013 1627 61047
rect 63785 61013 63819 61047
rect 66913 61013 66947 61047
rect 77953 61013 77987 61047
rect 63969 60809 64003 60843
rect 63785 60673 63819 60707
rect 64429 60673 64463 60707
rect 64613 60673 64647 60707
rect 64705 60673 64739 60707
rect 64802 60673 64836 60707
rect 65717 60673 65751 60707
rect 63601 60605 63635 60639
rect 65533 60605 65567 60639
rect 65901 60605 65935 60639
rect 66361 60605 66395 60639
rect 66637 60605 66671 60639
rect 62497 60537 62531 60571
rect 1409 60469 1443 60503
rect 63049 60469 63083 60503
rect 64981 60469 65015 60503
rect 62681 60265 62715 60299
rect 63969 60265 64003 60299
rect 66729 60265 66763 60299
rect 64981 60197 65015 60231
rect 66177 60197 66211 60231
rect 68109 60197 68143 60231
rect 68661 60129 68695 60163
rect 1409 60061 1443 60095
rect 62129 60061 62163 60095
rect 63601 60061 63635 60095
rect 63785 60061 63819 60095
rect 64429 60061 64463 60095
rect 64802 60061 64836 60095
rect 65625 60061 65659 60095
rect 65809 60061 65843 60095
rect 65901 60061 65935 60095
rect 65998 60061 66032 60095
rect 66913 60061 66947 60095
rect 67097 60061 67131 60095
rect 77493 60061 77527 60095
rect 78137 60061 78171 60095
rect 64613 59993 64647 60027
rect 64705 59993 64739 60027
rect 67649 59993 67683 60027
rect 1593 59925 1627 59959
rect 77953 59925 77987 59959
rect 62497 59721 62531 59755
rect 63509 59653 63543 59687
rect 64705 59653 64739 59687
rect 1409 59585 1443 59619
rect 2145 59585 2179 59619
rect 63325 59585 63359 59619
rect 63601 59585 63635 59619
rect 63745 59585 63779 59619
rect 64429 59585 64463 59619
rect 64613 59585 64647 59619
rect 64843 59585 64877 59619
rect 65553 59585 65587 59619
rect 65717 59585 65751 59619
rect 65809 59585 65843 59619
rect 65953 59585 65987 59619
rect 77309 59585 77343 59619
rect 77953 59585 77987 59619
rect 64998 59517 65032 59551
rect 66637 59449 66671 59483
rect 1593 59381 1627 59415
rect 61669 59381 61703 59415
rect 63877 59381 63911 59415
rect 66085 59381 66119 59415
rect 67189 59381 67223 59415
rect 77769 59381 77803 59415
rect 63325 59177 63359 59211
rect 64383 59177 64417 59211
rect 65809 59177 65843 59211
rect 62405 59109 62439 59143
rect 60749 59041 60783 59075
rect 1409 58973 1443 59007
rect 2145 58973 2179 59007
rect 61853 58973 61887 59007
rect 62226 58973 62260 59007
rect 63141 58973 63175 59007
rect 64613 58973 64647 59007
rect 65625 58973 65659 59007
rect 66821 58973 66855 59007
rect 77493 58973 77527 59007
rect 78137 58973 78171 59007
rect 62037 58905 62071 58939
rect 62129 58905 62163 58939
rect 66269 58905 66303 58939
rect 1593 58837 1627 58871
rect 59829 58837 59863 58871
rect 61301 58837 61335 58871
rect 67373 58837 67407 58871
rect 77953 58837 77987 58871
rect 59553 58633 59587 58667
rect 65993 58633 66027 58667
rect 66545 58633 66579 58667
rect 60289 58565 60323 58599
rect 62129 58565 62163 58599
rect 1409 58497 1443 58531
rect 2145 58497 2179 58531
rect 60013 58497 60047 58531
rect 60197 58497 60231 58531
rect 60386 58497 60420 58531
rect 61853 58497 61887 58531
rect 62037 58497 62071 58531
rect 62226 58497 62260 58531
rect 64705 58497 64739 58531
rect 77309 58497 77343 58531
rect 77953 58497 77987 58531
rect 63049 58429 63083 58463
rect 64981 58429 65015 58463
rect 65441 58429 65475 58463
rect 1593 58293 1627 58327
rect 60565 58293 60599 58327
rect 61117 58293 61151 58327
rect 62405 58293 62439 58327
rect 63601 58293 63635 58327
rect 77769 58293 77803 58327
rect 59277 57885 59311 57919
rect 59553 57885 59587 57919
rect 59697 57885 59731 57919
rect 60697 57885 60731 57919
rect 60841 57885 60875 57919
rect 61117 57885 61151 57919
rect 61761 57885 61795 57919
rect 62134 57885 62168 57919
rect 62330 57885 62364 57919
rect 62865 57885 62899 57919
rect 63238 57885 63272 57919
rect 65625 57885 65659 57919
rect 58725 57817 58759 57851
rect 59461 57817 59495 57851
rect 60933 57817 60967 57851
rect 61945 57817 61979 57851
rect 62037 57817 62071 57851
rect 63049 57817 63083 57851
rect 63141 57817 63175 57851
rect 64613 57817 64647 57851
rect 1409 57749 1443 57783
rect 59837 57749 59871 57783
rect 60557 57749 60591 57783
rect 63425 57749 63459 57783
rect 64061 57749 64095 57783
rect 78045 57749 78079 57783
rect 59645 57477 59679 57511
rect 1409 57409 1443 57443
rect 59369 57409 59403 57443
rect 59553 57409 59587 57443
rect 59742 57409 59776 57443
rect 62129 57409 62163 57443
rect 63049 57409 63083 57443
rect 63233 57409 63267 57443
rect 63325 57409 63359 57443
rect 63422 57409 63456 57443
rect 77953 57409 77987 57443
rect 61393 57341 61427 57375
rect 61669 57341 61703 57375
rect 64245 57341 64279 57375
rect 58817 57273 58851 57307
rect 63601 57273 63635 57307
rect 1593 57205 1627 57239
rect 58357 57205 58391 57239
rect 59921 57205 59955 57239
rect 77769 57205 77803 57239
rect 63049 57001 63083 57035
rect 59829 56933 59863 56967
rect 60749 56865 60783 56899
rect 1409 56797 1443 56831
rect 2145 56797 2179 56831
rect 59277 56797 59311 56831
rect 59461 56797 59495 56831
rect 59697 56797 59731 56831
rect 60473 56797 60507 56831
rect 61761 56797 61795 56831
rect 62037 56797 62071 56831
rect 77493 56797 77527 56831
rect 78137 56797 78171 56831
rect 58725 56729 58759 56763
rect 59553 56729 59587 56763
rect 1593 56661 1627 56695
rect 77953 56661 77987 56695
rect 59461 56457 59495 56491
rect 58541 56389 58575 56423
rect 1409 56321 1443 56355
rect 2145 56321 2179 56355
rect 60473 56321 60507 56355
rect 77309 56321 77343 56355
rect 77953 56321 77987 56355
rect 60749 56253 60783 56287
rect 61209 56253 61243 56287
rect 1593 56185 1627 56219
rect 57989 56185 58023 56219
rect 77769 56185 77803 56219
rect 57069 56117 57103 56151
rect 61439 56117 61473 56151
rect 55965 55913 55999 55947
rect 77953 55913 77987 55947
rect 57069 55845 57103 55879
rect 58173 55845 58207 55879
rect 58725 55777 58759 55811
rect 61025 55777 61059 55811
rect 56517 55709 56551 55743
rect 56793 55709 56827 55743
rect 56890 55709 56924 55743
rect 57621 55709 57655 55743
rect 57897 55709 57931 55743
rect 57994 55709 58028 55743
rect 60749 55709 60783 55743
rect 77493 55709 77527 55743
rect 78137 55709 78171 55743
rect 1501 55641 1535 55675
rect 1685 55641 1719 55675
rect 56701 55641 56735 55675
rect 57805 55641 57839 55675
rect 2145 55573 2179 55607
rect 55689 55369 55723 55403
rect 56517 55301 56551 55335
rect 58081 55301 58115 55335
rect 56241 55233 56275 55267
rect 56425 55233 56459 55267
rect 56661 55233 56695 55267
rect 57897 55233 57931 55267
rect 58173 55233 58207 55267
rect 58270 55233 58304 55267
rect 58466 55233 58500 55267
rect 60565 55233 60599 55267
rect 61209 55233 61243 55267
rect 59001 55097 59035 55131
rect 1501 55029 1535 55063
rect 56793 55029 56827 55063
rect 77953 55029 77987 55063
rect 59001 54825 59035 54859
rect 56333 54689 56367 54723
rect 57897 54689 57931 54723
rect 1501 54621 1535 54655
rect 56609 54621 56643 54655
rect 57621 54621 57655 54655
rect 77493 54621 77527 54655
rect 78137 54621 78171 54655
rect 1593 54485 1627 54519
rect 77953 54485 77987 54519
rect 55505 54281 55539 54315
rect 56241 54213 56275 54247
rect 1501 54145 1535 54179
rect 2145 54145 2179 54179
rect 56057 54145 56091 54179
rect 56333 54145 56367 54179
rect 56477 54145 56511 54179
rect 77677 54077 77711 54111
rect 77953 54077 77987 54111
rect 1685 54009 1719 54043
rect 56609 53941 56643 53975
rect 57253 53941 57287 53975
rect 76849 53533 76883 53567
rect 77309 53533 77343 53567
rect 77585 53533 77619 53567
rect 1501 53465 1535 53499
rect 2145 53465 2179 53499
rect 53849 53465 53883 53499
rect 1593 53397 1627 53431
rect 54309 53397 54343 53431
rect 53297 53125 53331 53159
rect 1501 53057 1535 53091
rect 2145 53057 2179 53091
rect 53021 53057 53055 53091
rect 53205 53057 53239 53091
rect 53441 53057 53475 53091
rect 54125 53057 54159 53091
rect 54309 53057 54343 53091
rect 54401 53057 54435 53091
rect 54498 53057 54532 53091
rect 77677 53057 77711 53091
rect 77953 52989 77987 53023
rect 1685 52921 1719 52955
rect 53573 52853 53607 52887
rect 54677 52853 54711 52887
rect 55321 52853 55355 52887
rect 52837 52649 52871 52683
rect 77585 52581 77619 52615
rect 52377 52513 52411 52547
rect 53389 52445 53423 52479
rect 53665 52445 53699 52479
rect 1501 52309 1535 52343
rect 54769 52309 54803 52343
rect 78045 52309 78079 52343
rect 51825 52037 51859 52071
rect 54861 52037 54895 52071
rect 1501 51969 1535 52003
rect 51549 51969 51583 52003
rect 51733 51969 51767 52003
rect 51969 51969 52003 52003
rect 53389 51969 53423 52003
rect 54625 51969 54659 52003
rect 54769 51969 54803 52003
rect 55045 51969 55079 52003
rect 53113 51901 53147 51935
rect 77677 51901 77711 51935
rect 77953 51901 77987 51935
rect 51089 51833 51123 51867
rect 1593 51765 1627 51799
rect 52101 51765 52135 51799
rect 54493 51765 54527 51799
rect 55597 51765 55631 51799
rect 52377 51493 52411 51527
rect 52929 51425 52963 51459
rect 51365 51357 51399 51391
rect 51825 51357 51859 51391
rect 52009 51357 52043 51391
rect 52198 51357 52232 51391
rect 53205 51357 53239 51391
rect 76849 51357 76883 51391
rect 77309 51357 77343 51391
rect 77585 51357 77619 51391
rect 1501 51289 1535 51323
rect 1685 51289 1719 51323
rect 52101 51289 52135 51323
rect 54309 51289 54343 51323
rect 2145 51221 2179 51255
rect 1501 50881 1535 50915
rect 2145 50881 2179 50915
rect 53205 50881 53239 50915
rect 53481 50813 53515 50847
rect 76665 50813 76699 50847
rect 77125 50813 77159 50847
rect 77401 50813 77435 50847
rect 1685 50745 1719 50779
rect 50261 50473 50295 50507
rect 52009 50473 52043 50507
rect 51365 50405 51399 50439
rect 53389 50405 53423 50439
rect 50813 50269 50847 50303
rect 51089 50269 51123 50303
rect 51233 50269 51267 50303
rect 52837 50269 52871 50303
rect 53257 50269 53291 50303
rect 77309 50269 77343 50303
rect 77585 50269 77619 50303
rect 1501 50201 1535 50235
rect 1685 50201 1719 50235
rect 50997 50201 51031 50235
rect 53021 50201 53055 50235
rect 53113 50201 53147 50235
rect 2145 50133 2179 50167
rect 54033 50133 54067 50167
rect 49801 49929 49835 49963
rect 52745 49929 52779 49963
rect 50537 49861 50571 49895
rect 50629 49861 50663 49895
rect 77401 49861 77435 49895
rect 50353 49793 50387 49827
rect 50773 49793 50807 49827
rect 51549 49725 51583 49759
rect 50905 49657 50939 49691
rect 1501 49589 1535 49623
rect 77953 49589 77987 49623
rect 50721 49317 50755 49351
rect 1501 49181 1535 49215
rect 50169 49181 50203 49215
rect 50353 49181 50387 49215
rect 50589 49181 50623 49215
rect 77861 49181 77895 49215
rect 78137 49181 78171 49215
rect 50445 49113 50479 49147
rect 1593 49045 1627 49079
rect 49525 49045 49559 49079
rect 51365 49045 51399 49079
rect 50353 48773 50387 48807
rect 1501 48705 1535 48739
rect 2145 48705 2179 48739
rect 50169 48705 50203 48739
rect 50445 48705 50479 48739
rect 50589 48705 50623 48739
rect 76665 48637 76699 48671
rect 77125 48637 77159 48671
rect 77401 48637 77435 48671
rect 1685 48569 1719 48603
rect 49709 48501 49743 48535
rect 50721 48501 50755 48535
rect 51365 48501 51399 48535
rect 1685 48093 1719 48127
rect 77861 48093 77895 48127
rect 2237 48025 2271 48059
rect 1501 47957 1535 47991
rect 48145 47957 48179 47991
rect 77309 47957 77343 47991
rect 78045 47957 78079 47991
rect 47777 47753 47811 47787
rect 1685 47617 1719 47651
rect 2237 47617 2271 47651
rect 47869 47617 47903 47651
rect 48881 47617 48915 47651
rect 77677 47617 77711 47651
rect 49065 47481 49099 47515
rect 1501 47413 1535 47447
rect 49525 47413 49559 47447
rect 77125 47413 77159 47447
rect 77861 47413 77895 47447
rect 47133 47209 47167 47243
rect 47225 47005 47259 47039
rect 48145 47005 48179 47039
rect 48789 47005 48823 47039
rect 48329 46937 48363 46971
rect 47685 46665 47719 46699
rect 1685 46529 1719 46563
rect 2237 46529 2271 46563
rect 77677 46529 77711 46563
rect 1501 46393 1535 46427
rect 77861 46393 77895 46427
rect 46765 46325 46799 46359
rect 77125 46325 77159 46359
rect 46397 46121 46431 46155
rect 1685 45917 1719 45951
rect 46489 45917 46523 45951
rect 47409 45917 47443 45951
rect 48053 45917 48087 45951
rect 77309 45917 77343 45951
rect 77861 45917 77895 45951
rect 47593 45849 47627 45883
rect 1501 45781 1535 45815
rect 2237 45781 2271 45815
rect 78045 45781 78079 45815
rect 46857 45509 46891 45543
rect 1685 45441 1719 45475
rect 2237 45441 2271 45475
rect 45753 45441 45787 45475
rect 46673 45441 46707 45475
rect 47593 45441 47627 45475
rect 77677 45441 77711 45475
rect 45109 45373 45143 45407
rect 45569 45305 45603 45339
rect 1501 45237 1535 45271
rect 77125 45237 77159 45271
rect 77861 45237 77895 45271
rect 45109 45033 45143 45067
rect 1685 44829 1719 44863
rect 2237 44829 2271 44863
rect 77861 44829 77895 44863
rect 45201 44761 45235 44795
rect 45937 44761 45971 44795
rect 46121 44761 46155 44795
rect 1501 44693 1535 44727
rect 46581 44693 46615 44727
rect 77309 44693 77343 44727
rect 78045 44693 78079 44727
rect 44281 44489 44315 44523
rect 43729 44353 43763 44387
rect 44373 44353 44407 44387
rect 45201 44353 45235 44387
rect 45845 44353 45879 44387
rect 45385 44217 45419 44251
rect 46397 44149 46431 44183
rect 1685 43741 1719 43775
rect 2237 43741 2271 43775
rect 77861 43741 77895 43775
rect 1501 43605 1535 43639
rect 43913 43605 43947 43639
rect 44373 43605 44407 43639
rect 77309 43605 77343 43639
rect 78045 43605 78079 43639
rect 43545 43401 43579 43435
rect 1685 43265 1719 43299
rect 43637 43265 43671 43299
rect 44465 43265 44499 43299
rect 77677 43265 77711 43299
rect 44649 43129 44683 43163
rect 1501 43061 1535 43095
rect 2237 43061 2271 43095
rect 77125 43061 77159 43095
rect 77861 43061 77895 43095
rect 1685 42653 1719 42687
rect 42717 42653 42751 42687
rect 77861 42653 77895 42687
rect 2237 42585 2271 42619
rect 42901 42585 42935 42619
rect 43729 42585 43763 42619
rect 43913 42585 43947 42619
rect 1501 42517 1535 42551
rect 42257 42517 42291 42551
rect 44373 42517 44407 42551
rect 77309 42517 77343 42551
rect 78045 42517 78079 42551
rect 42533 42313 42567 42347
rect 1685 42177 1719 42211
rect 42625 42177 42659 42211
rect 43269 42177 43303 42211
rect 43913 42177 43947 42211
rect 77677 42177 77711 42211
rect 2237 42041 2271 42075
rect 43453 42041 43487 42075
rect 1501 41973 1535 42007
rect 77125 41973 77159 42007
rect 77861 41973 77895 42007
rect 41337 41701 41371 41735
rect 41521 41565 41555 41599
rect 42349 41565 42383 41599
rect 42533 41497 42567 41531
rect 43085 41429 43119 41463
rect 1685 41089 1719 41123
rect 77677 41089 77711 41123
rect 1501 40953 1535 40987
rect 2237 40953 2271 40987
rect 77861 40953 77895 40987
rect 41061 40885 41095 40919
rect 41797 40885 41831 40919
rect 42625 40885 42659 40919
rect 77125 40885 77159 40919
rect 40693 40681 40727 40715
rect 1685 40477 1719 40511
rect 77861 40477 77895 40511
rect 40785 40409 40819 40443
rect 41613 40409 41647 40443
rect 41797 40409 41831 40443
rect 1501 40341 1535 40375
rect 2237 40341 2271 40375
rect 77309 40341 77343 40375
rect 78045 40341 78079 40375
rect 1685 40001 1719 40035
rect 39405 40001 39439 40035
rect 40049 40001 40083 40035
rect 40877 40001 40911 40035
rect 41061 40001 41095 40035
rect 77677 40001 77711 40035
rect 39865 39933 39899 39967
rect 2237 39865 2271 39899
rect 1501 39797 1535 39831
rect 41521 39797 41555 39831
rect 77125 39797 77159 39831
rect 77861 39797 77895 39831
rect 39129 39593 39163 39627
rect 1685 39389 1719 39423
rect 77861 39389 77895 39423
rect 2237 39321 2271 39355
rect 38577 39321 38611 39355
rect 39221 39321 39255 39355
rect 40141 39321 40175 39355
rect 40325 39321 40359 39355
rect 1501 39253 1535 39287
rect 40785 39253 40819 39287
rect 77309 39253 77343 39287
rect 78045 39253 78079 39287
rect 38485 39049 38519 39083
rect 37933 38913 37967 38947
rect 38577 38913 38611 38947
rect 39405 38913 39439 38947
rect 39589 38777 39623 38811
rect 40049 38709 40083 38743
rect 1685 38301 1719 38335
rect 77861 38301 77895 38335
rect 2237 38233 2271 38267
rect 1501 38165 1535 38199
rect 38393 38165 38427 38199
rect 39129 38165 39163 38199
rect 77309 38165 77343 38199
rect 78045 38165 78079 38199
rect 37749 37961 37783 37995
rect 1685 37825 1719 37859
rect 37841 37825 37875 37859
rect 38669 37825 38703 37859
rect 77677 37825 77711 37859
rect 2237 37689 2271 37723
rect 38853 37689 38887 37723
rect 1501 37621 1535 37655
rect 77125 37621 77159 37655
rect 77861 37621 77895 37655
rect 37013 37417 37047 37451
rect 38577 37349 38611 37383
rect 38117 37281 38151 37315
rect 1685 37213 1719 37247
rect 77861 37213 77895 37247
rect 2237 37145 2271 37179
rect 36461 37145 36495 37179
rect 37105 37145 37139 37179
rect 37933 37145 37967 37179
rect 1501 37077 1535 37111
rect 77309 37077 77343 37111
rect 78045 37077 78079 37111
rect 36277 36873 36311 36907
rect 38025 36873 38059 36907
rect 1685 36737 1719 36771
rect 2237 36737 2271 36771
rect 35725 36737 35759 36771
rect 36369 36737 36403 36771
rect 37381 36737 37415 36771
rect 77677 36737 77711 36771
rect 37565 36601 37599 36635
rect 1501 36533 1535 36567
rect 77125 36533 77159 36567
rect 77861 36533 77895 36567
rect 35633 36329 35667 36363
rect 37197 36329 37231 36363
rect 35081 36057 35115 36091
rect 35725 36057 35759 36091
rect 36553 36057 36587 36091
rect 36737 36057 36771 36091
rect 1685 35649 1719 35683
rect 77677 35649 77711 35683
rect 1501 35513 1535 35547
rect 2237 35513 2271 35547
rect 77861 35513 77895 35547
rect 35633 35445 35667 35479
rect 36277 35445 36311 35479
rect 77125 35445 77159 35479
rect 34897 35241 34931 35275
rect 1685 35037 1719 35071
rect 2237 35037 2271 35071
rect 77861 35037 77895 35071
rect 34989 34969 35023 35003
rect 35817 34969 35851 35003
rect 1501 34901 1535 34935
rect 35909 34901 35943 34935
rect 77309 34901 77343 34935
rect 78045 34901 78079 34935
rect 34161 34697 34195 34731
rect 35725 34697 35759 34731
rect 35265 34629 35299 34663
rect 1685 34561 1719 34595
rect 33609 34561 33643 34595
rect 34253 34561 34287 34595
rect 35081 34561 35115 34595
rect 77677 34561 77711 34595
rect 2237 34493 2271 34527
rect 77125 34493 77159 34527
rect 1501 34357 1535 34391
rect 77861 34357 77895 34391
rect 1685 33949 1719 33983
rect 33333 33949 33367 33983
rect 77861 33949 77895 33983
rect 2237 33881 2271 33915
rect 33517 33881 33551 33915
rect 34805 33881 34839 33915
rect 34989 33881 35023 33915
rect 1501 33813 1535 33847
rect 32873 33813 32907 33847
rect 34069 33813 34103 33847
rect 35449 33813 35483 33847
rect 77309 33813 77343 33847
rect 78045 33813 78079 33847
rect 32689 33609 32723 33643
rect 32781 33473 32815 33507
rect 33701 33473 33735 33507
rect 34345 33473 34379 33507
rect 33885 33337 33919 33371
rect 1685 32861 1719 32895
rect 77861 32861 77895 32895
rect 2237 32793 2271 32827
rect 1501 32725 1535 32759
rect 32781 32725 32815 32759
rect 33425 32725 33459 32759
rect 77309 32725 77343 32759
rect 78045 32725 78079 32759
rect 32229 32521 32263 32555
rect 1685 32385 1719 32419
rect 2237 32385 2271 32419
rect 32321 32385 32355 32419
rect 32965 32385 32999 32419
rect 77677 32385 77711 32419
rect 33149 32249 33183 32283
rect 1501 32181 1535 32215
rect 77125 32181 77159 32215
rect 77861 32181 77895 32215
rect 31217 31977 31251 32011
rect 77309 31909 77343 31943
rect 78045 31909 78079 31943
rect 32505 31841 32539 31875
rect 1685 31773 1719 31807
rect 2237 31773 2271 31807
rect 32965 31773 32999 31807
rect 77861 31773 77895 31807
rect 31309 31705 31343 31739
rect 32321 31705 32355 31739
rect 1501 31637 1535 31671
rect 32413 31365 32447 31399
rect 1685 31297 1719 31331
rect 29929 31297 29963 31331
rect 30573 31297 30607 31331
rect 32229 31297 32263 31331
rect 77677 31297 77711 31331
rect 30389 31229 30423 31263
rect 2237 31161 2271 31195
rect 1501 31093 1535 31127
rect 31585 31093 31619 31127
rect 32873 31093 32907 31127
rect 77125 31093 77159 31127
rect 77861 31093 77895 31127
rect 29745 30889 29779 30923
rect 29837 30617 29871 30651
rect 30941 30617 30975 30651
rect 31125 30617 31159 30651
rect 31953 30549 31987 30583
rect 1685 30209 1719 30243
rect 77677 30209 77711 30243
rect 1501 30073 1535 30107
rect 2237 30073 2271 30107
rect 77861 30073 77895 30107
rect 29193 30005 29227 30039
rect 30113 30005 30147 30039
rect 30665 30005 30699 30039
rect 77125 30005 77159 30039
rect 28825 29801 28859 29835
rect 1685 29597 1719 29631
rect 2237 29597 2271 29631
rect 77861 29597 77895 29631
rect 28917 29529 28951 29563
rect 30205 29529 30239 29563
rect 30389 29529 30423 29563
rect 1501 29461 1535 29495
rect 29561 29461 29595 29495
rect 77309 29461 77343 29495
rect 78045 29461 78079 29495
rect 28273 29257 28307 29291
rect 1685 29121 1719 29155
rect 27721 29121 27755 29155
rect 28365 29121 28399 29155
rect 29561 29121 29595 29155
rect 29745 29121 29779 29155
rect 77677 29121 77711 29155
rect 2237 29053 2271 29087
rect 1501 28985 1535 29019
rect 28917 28985 28951 29019
rect 77125 28985 77159 29019
rect 77861 28985 77895 29019
rect 27445 28645 27479 28679
rect 1685 28509 1719 28543
rect 2237 28509 2271 28543
rect 77861 28509 77895 28543
rect 26985 28441 27019 28475
rect 27629 28441 27663 28475
rect 28825 28441 28859 28475
rect 29009 28441 29043 28475
rect 1501 28373 1535 28407
rect 28181 28373 28215 28407
rect 77309 28373 77343 28407
rect 78045 28373 78079 28407
rect 27077 28169 27111 28203
rect 27169 28033 27203 28067
rect 28181 28033 28215 28067
rect 28273 27829 28307 27863
rect 1685 27421 1719 27455
rect 2237 27421 2271 27455
rect 77861 27421 77895 27455
rect 1501 27285 1535 27319
rect 26341 27285 26375 27319
rect 27445 27285 27479 27319
rect 27905 27285 27939 27319
rect 77309 27285 77343 27319
rect 78045 27285 78079 27319
rect 26065 27081 26099 27115
rect 1685 26945 1719 26979
rect 2237 26945 2271 26979
rect 26157 26945 26191 26979
rect 27445 26945 27479 26979
rect 77677 26945 77711 26979
rect 27629 26809 27663 26843
rect 1501 26741 1535 26775
rect 77125 26741 77159 26775
rect 77861 26741 77895 26775
rect 25237 26537 25271 26571
rect 78045 26469 78079 26503
rect 27353 26401 27387 26435
rect 1685 26333 1719 26367
rect 2237 26333 2271 26367
rect 26893 26333 26927 26367
rect 77401 26333 77435 26367
rect 77861 26333 77895 26367
rect 25329 26265 25363 26299
rect 26709 26265 26743 26299
rect 1501 26197 1535 26231
rect 26065 26197 26099 26231
rect 32505 26197 32539 26231
rect 22845 25925 22879 25959
rect 32689 25925 32723 25959
rect 1685 25857 1719 25891
rect 23029 25857 23063 25891
rect 23581 25857 23615 25891
rect 77677 25857 77711 25891
rect 2237 25721 2271 25755
rect 77125 25721 77159 25755
rect 1501 25653 1535 25687
rect 25605 25653 25639 25687
rect 32781 25653 32815 25687
rect 77861 25653 77895 25687
rect 22293 25449 22327 25483
rect 22477 25245 22511 25279
rect 22937 25245 22971 25279
rect 32597 25177 32631 25211
rect 31953 25109 31987 25143
rect 32689 25109 32723 25143
rect 41622 24837 41656 24871
rect 1685 24769 1719 24803
rect 2237 24769 2271 24803
rect 41245 24769 41279 24803
rect 77677 24769 77711 24803
rect 1501 24633 1535 24667
rect 40785 24633 40819 24667
rect 41797 24633 41831 24667
rect 77861 24633 77895 24667
rect 41613 24565 41647 24599
rect 77125 24565 77159 24599
rect 22293 24361 22327 24395
rect 41705 24361 41739 24395
rect 1685 24157 1719 24191
rect 2237 24157 2271 24191
rect 22477 24157 22511 24191
rect 32229 24157 32263 24191
rect 41981 24157 42015 24191
rect 77861 24157 77895 24191
rect 23029 24089 23063 24123
rect 31493 24089 31527 24123
rect 32045 24089 32079 24123
rect 40969 24089 41003 24123
rect 41521 24089 41555 24123
rect 1501 24021 1535 24055
rect 41705 24021 41739 24055
rect 77309 24021 77343 24055
rect 78045 24021 78079 24055
rect 21833 23817 21867 23851
rect 30849 23817 30883 23851
rect 1685 23681 1719 23715
rect 22017 23681 22051 23715
rect 31401 23681 31435 23715
rect 31585 23681 31619 23715
rect 32229 23681 32263 23715
rect 32873 23681 32907 23715
rect 41705 23681 41739 23715
rect 77677 23681 77711 23715
rect 32413 23613 32447 23647
rect 2237 23545 2271 23579
rect 31585 23545 31619 23579
rect 1501 23477 1535 23511
rect 22569 23477 22603 23511
rect 41245 23477 41279 23511
rect 77125 23477 77159 23511
rect 77861 23477 77895 23511
rect 19717 23273 19751 23307
rect 31401 23273 31435 23307
rect 31585 23273 31619 23307
rect 27997 23137 28031 23171
rect 1685 23069 1719 23103
rect 19901 23069 19935 23103
rect 31585 23069 31619 23103
rect 31953 23069 31987 23103
rect 32045 23069 32079 23103
rect 77861 23069 77895 23103
rect 2237 23001 2271 23035
rect 27813 23001 27847 23035
rect 30941 23001 30975 23035
rect 1501 22933 1535 22967
rect 20453 22933 20487 22967
rect 27169 22933 27203 22967
rect 30389 22933 30423 22967
rect 77309 22933 77343 22967
rect 78045 22933 78079 22967
rect 19993 22729 20027 22763
rect 31125 22729 31159 22763
rect 20177 22593 20211 22627
rect 27813 22593 27847 22627
rect 27997 22457 28031 22491
rect 20729 22389 20763 22423
rect 27169 22389 27203 22423
rect 1685 21981 1719 22015
rect 77861 21981 77895 22015
rect 27445 21913 27479 21947
rect 27997 21913 28031 21947
rect 1501 21845 1535 21879
rect 28089 21845 28123 21879
rect 77309 21845 77343 21879
rect 78045 21845 78079 21879
rect 19073 21641 19107 21675
rect 1685 21505 1719 21539
rect 19257 21505 19291 21539
rect 77677 21505 77711 21539
rect 1501 21301 1535 21335
rect 19809 21301 19843 21335
rect 77125 21301 77159 21335
rect 77861 21301 77895 21335
rect 17877 21097 17911 21131
rect 1685 20893 1719 20927
rect 18061 20893 18095 20927
rect 18613 20893 18647 20927
rect 77309 20893 77343 20927
rect 77861 20893 77895 20927
rect 27813 20825 27847 20859
rect 1501 20757 1535 20791
rect 27169 20757 27203 20791
rect 27905 20757 27939 20791
rect 78045 20757 78079 20791
rect 18521 20553 18555 20587
rect 32413 20485 32447 20519
rect 1685 20417 1719 20451
rect 18705 20417 18739 20451
rect 32229 20417 32263 20451
rect 77677 20417 77711 20451
rect 1501 20213 1535 20247
rect 19257 20213 19291 20247
rect 31493 20213 31527 20247
rect 77125 20213 77159 20247
rect 77861 20213 77895 20247
rect 17049 20009 17083 20043
rect 17233 19805 17267 19839
rect 31585 19737 31619 19771
rect 31769 19737 31803 19771
rect 17785 19669 17819 19703
rect 30941 19669 30975 19703
rect 16681 19465 16715 19499
rect 77861 19465 77895 19499
rect 1685 19329 1719 19363
rect 16865 19329 16899 19363
rect 30573 19329 30607 19363
rect 32229 19329 32263 19363
rect 77677 19329 77711 19363
rect 1501 19193 1535 19227
rect 17417 19125 17451 19159
rect 31493 19125 31527 19159
rect 32321 19125 32355 19159
rect 77125 19125 77159 19159
rect 31125 18921 31159 18955
rect 31585 18921 31619 18955
rect 31217 18785 31251 18819
rect 1685 18717 1719 18751
rect 16313 18717 16347 18751
rect 31125 18717 31159 18751
rect 31401 18717 31435 18751
rect 77861 18717 77895 18751
rect 30021 18649 30055 18683
rect 32137 18649 32171 18683
rect 1501 18581 1535 18615
rect 16129 18581 16163 18615
rect 16865 18581 16899 18615
rect 26341 18581 26375 18615
rect 26985 18581 27019 18615
rect 30573 18581 30607 18615
rect 32229 18581 32263 18615
rect 77309 18581 77343 18615
rect 78045 18581 78079 18615
rect 32137 18377 32171 18411
rect 26433 18309 26467 18343
rect 30849 18309 30883 18343
rect 1685 18241 1719 18275
rect 27077 18241 27111 18275
rect 27353 18241 27387 18275
rect 77677 18241 77711 18275
rect 27169 18173 27203 18207
rect 1501 18037 1535 18071
rect 27077 18037 27111 18071
rect 27537 18037 27571 18071
rect 77125 18037 77159 18071
rect 77861 18037 77895 18071
rect 14841 17833 14875 17867
rect 27721 17697 27755 17731
rect 1685 17629 1719 17663
rect 15025 17629 15059 17663
rect 27353 17629 27387 17663
rect 27537 17629 27571 17663
rect 77861 17629 77895 17663
rect 1501 17493 1535 17527
rect 15577 17493 15611 17527
rect 26525 17493 26559 17527
rect 27813 17493 27847 17527
rect 77309 17493 77343 17527
rect 78045 17493 78079 17527
rect 14473 17289 14507 17323
rect 14657 17153 14691 17187
rect 26433 17153 26467 17187
rect 27537 17153 27571 17187
rect 27721 17017 27755 17051
rect 15209 16949 15243 16983
rect 28181 16949 28215 16983
rect 26249 16745 26283 16779
rect 28181 16745 28215 16779
rect 27537 16677 27571 16711
rect 77309 16677 77343 16711
rect 1685 16541 1719 16575
rect 28089 16541 28123 16575
rect 77861 16541 77895 16575
rect 27353 16473 27387 16507
rect 1501 16405 1535 16439
rect 26709 16405 26743 16439
rect 78045 16405 78079 16439
rect 12725 16201 12759 16235
rect 25881 16201 25915 16235
rect 27445 16201 27479 16235
rect 26985 16133 27019 16167
rect 1685 16065 1719 16099
rect 12909 16065 12943 16099
rect 13645 16065 13679 16099
rect 27261 16065 27295 16099
rect 27997 16065 28031 16099
rect 77677 16065 77711 16099
rect 27077 15997 27111 16031
rect 13461 15929 13495 15963
rect 1501 15861 1535 15895
rect 14105 15861 14139 15895
rect 26433 15861 26467 15895
rect 27261 15861 27295 15895
rect 28089 15861 28123 15895
rect 77125 15861 77159 15895
rect 77861 15861 77895 15895
rect 27721 15657 27755 15691
rect 26709 15589 26743 15623
rect 1685 15453 1719 15487
rect 77861 15453 77895 15487
rect 77309 15385 77343 15419
rect 1501 15317 1535 15351
rect 13093 15317 13127 15351
rect 78045 15317 78079 15351
rect 11529 15113 11563 15147
rect 27721 15045 27755 15079
rect 1685 14977 1719 15011
rect 11713 14977 11747 15011
rect 26433 14977 26467 15011
rect 27537 14977 27571 15011
rect 77677 14977 77711 15011
rect 1501 14773 1535 14807
rect 12265 14773 12299 14807
rect 77125 14773 77159 14807
rect 77861 14773 77895 14807
rect 11529 14569 11563 14603
rect 11713 14365 11747 14399
rect 26801 14297 26835 14331
rect 27353 14297 27387 14331
rect 12265 14229 12299 14263
rect 27445 14229 27479 14263
rect 10425 14025 10459 14059
rect 27353 14025 27387 14059
rect 77861 14025 77895 14059
rect 1685 13889 1719 13923
rect 10609 13889 10643 13923
rect 25789 13889 25823 13923
rect 26985 13889 27019 13923
rect 27077 13889 27111 13923
rect 27905 13889 27939 13923
rect 77677 13889 77711 13923
rect 11621 13821 11655 13855
rect 26433 13821 26467 13855
rect 28089 13821 28123 13855
rect 77125 13821 77159 13855
rect 1501 13753 1535 13787
rect 26985 13685 27019 13719
rect 26709 13481 26743 13515
rect 27721 13481 27755 13515
rect 1685 13277 1719 13311
rect 9597 13277 9631 13311
rect 77861 13277 77895 13311
rect 10149 13209 10183 13243
rect 42165 13209 42199 13243
rect 1501 13141 1535 13175
rect 9413 13141 9447 13175
rect 41521 13141 41555 13175
rect 42257 13141 42291 13175
rect 77309 13141 77343 13175
rect 78045 13141 78079 13175
rect 1685 12801 1719 12835
rect 77677 12801 77711 12835
rect 1501 12597 1535 12631
rect 77125 12597 77159 12631
rect 77861 12597 77895 12631
rect 9689 12393 9723 12427
rect 1685 12189 1719 12223
rect 9873 12189 9907 12223
rect 12633 12189 12667 12223
rect 77861 12189 77895 12223
rect 1501 12053 1535 12087
rect 12817 12053 12851 12087
rect 77309 12053 77343 12087
rect 78045 12053 78079 12087
rect 9045 11849 9079 11883
rect 9229 11713 9263 11747
rect 11989 11713 12023 11747
rect 12173 11509 12207 11543
rect 1501 11237 1535 11271
rect 78045 11237 78079 11271
rect 1685 11101 1719 11135
rect 77861 11101 77895 11135
rect 77309 11033 77343 11067
rect 8309 10761 8343 10795
rect 11713 10761 11747 10795
rect 1685 10625 1719 10659
rect 8493 10625 8527 10659
rect 11529 10625 11563 10659
rect 77677 10625 77711 10659
rect 1501 10421 1535 10455
rect 77125 10421 77159 10455
rect 77861 10421 77895 10455
rect 7573 10217 7607 10251
rect 1685 10013 1719 10047
rect 7757 10013 7791 10047
rect 10701 10013 10735 10047
rect 77861 10013 77895 10047
rect 1501 9877 1535 9911
rect 10885 9877 10919 9911
rect 77309 9877 77343 9911
rect 78045 9877 78079 9911
rect 6745 9673 6779 9707
rect 10149 9673 10183 9707
rect 1685 9537 1719 9571
rect 6929 9537 6963 9571
rect 9965 9537 9999 9571
rect 77677 9537 77711 9571
rect 1501 9333 1535 9367
rect 77125 9333 77159 9367
rect 77861 9333 77895 9367
rect 6009 9129 6043 9163
rect 6193 8925 6227 8959
rect 9321 8925 9355 8959
rect 9505 8789 9539 8823
rect 1685 8449 1719 8483
rect 77677 8449 77711 8483
rect 1501 8313 1535 8347
rect 77125 8313 77159 8347
rect 77861 8313 77895 8347
rect 5273 8041 5307 8075
rect 1685 7837 1719 7871
rect 5457 7837 5491 7871
rect 8953 7837 8987 7871
rect 77861 7837 77895 7871
rect 77309 7769 77343 7803
rect 1501 7701 1535 7735
rect 9137 7701 9171 7735
rect 78045 7701 78079 7735
rect 4537 7497 4571 7531
rect 1685 7361 1719 7395
rect 4721 7361 4755 7395
rect 8033 7361 8067 7395
rect 77677 7361 77711 7395
rect 8217 7225 8251 7259
rect 1501 7157 1535 7191
rect 77125 7157 77159 7191
rect 77861 7157 77895 7191
rect 3893 6953 3927 6987
rect 1685 6749 1719 6783
rect 4077 6749 4111 6783
rect 7481 6749 7515 6783
rect 77861 6749 77895 6783
rect 1501 6613 1535 6647
rect 7665 6613 7699 6647
rect 77309 6613 77343 6647
rect 78045 6613 78079 6647
rect 3249 6409 3283 6443
rect 3433 6273 3467 6307
rect 6929 6273 6963 6307
rect 7113 6069 7147 6103
rect 1685 5661 1719 5695
rect 77309 5661 77343 5695
rect 77861 5661 77895 5695
rect 1501 5525 1535 5559
rect 78045 5525 78079 5559
rect 2605 5321 2639 5355
rect 6653 5321 6687 5355
rect 1685 5185 1719 5219
rect 2789 5185 2823 5219
rect 6469 5185 6503 5219
rect 77677 5185 77711 5219
rect 1501 4981 1535 5015
rect 77125 4981 77159 5015
rect 77861 4981 77895 5015
rect 2053 4777 2087 4811
rect 2237 4573 2271 4607
rect 6009 4573 6043 4607
rect 6193 4437 6227 4471
rect 53849 3689 53883 3723
rect 64337 3689 64371 3723
rect 27445 3553 27479 3587
rect 69489 3553 69523 3587
rect 26709 3485 26743 3519
rect 27169 3485 27203 3519
rect 30481 3417 30515 3451
rect 28457 3349 28491 3383
rect 30021 3349 30055 3383
rect 32229 3349 32263 3383
rect 32965 3349 32999 3383
rect 33701 3349 33735 3383
rect 43729 3349 43763 3383
rect 74733 3349 74767 3383
rect 78045 3349 78079 3383
rect 3801 3145 3835 3179
rect 8953 3145 8987 3179
rect 14105 3145 14139 3179
rect 24409 3145 24443 3179
rect 32505 3145 32539 3179
rect 33241 3145 33275 3179
rect 34713 3145 34747 3179
rect 39865 3145 39899 3179
rect 44281 3145 44315 3179
rect 49985 3145 50019 3179
rect 50629 3145 50663 3179
rect 51273 3145 51307 3179
rect 51825 3145 51859 3179
rect 52745 3145 52779 3179
rect 53297 3145 53331 3179
rect 55229 3145 55263 3179
rect 56517 3145 56551 3179
rect 57161 3145 57195 3179
rect 58449 3145 58483 3179
rect 59001 3145 59035 3179
rect 60289 3145 60323 3179
rect 60841 3145 60875 3179
rect 64153 3145 64187 3179
rect 66913 3145 66947 3179
rect 69305 3145 69339 3179
rect 70593 3145 70627 3179
rect 72065 3145 72099 3179
rect 75193 3145 75227 3179
rect 77769 3145 77803 3179
rect 19349 3077 19383 3111
rect 53849 3077 53883 3111
rect 57989 3077 58023 3111
rect 61393 3077 61427 3111
rect 63601 3077 63635 3111
rect 68201 3077 68235 3111
rect 3617 3009 3651 3043
rect 4261 3009 4295 3043
rect 8309 3009 8343 3043
rect 8769 3009 8803 3043
rect 13461 3009 13495 3043
rect 14013 3009 14047 3043
rect 18613 3009 18647 3043
rect 19165 3009 19199 3043
rect 23765 3009 23799 3043
rect 24317 3009 24351 3043
rect 26157 3009 26191 3043
rect 28089 3009 28123 3043
rect 29377 3009 29411 3043
rect 30389 3009 30423 3043
rect 32413 3009 32447 3043
rect 33149 3009 33183 3043
rect 34069 3009 34103 3043
rect 34621 3009 34655 3043
rect 39221 3009 39255 3043
rect 39773 3009 39807 3043
rect 43637 3009 43671 3043
rect 44189 3009 44223 3043
rect 49525 3009 49559 3043
rect 54401 3009 54435 3043
rect 59829 3009 59863 3043
rect 64705 3009 64739 3043
rect 68753 3009 68787 3043
rect 69857 3009 69891 3043
rect 74549 3009 74583 3043
rect 75009 3009 75043 3043
rect 77953 3009 77987 3043
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 28365 2941 28399 2975
rect 29653 2941 29687 2975
rect 30113 2941 30147 2975
rect 61945 2941 61979 2975
rect 65441 2941 65475 2975
rect 66269 2873 66303 2907
rect 71329 2873 71363 2907
rect 77125 2873 77159 2907
rect 2789 2805 2823 2839
rect 5181 2805 5215 2839
rect 5733 2805 5767 2839
rect 6469 2805 6503 2839
rect 7205 2805 7239 2839
rect 7757 2805 7791 2839
rect 9689 2805 9723 2839
rect 10333 2805 10367 2839
rect 10885 2805 10919 2839
rect 11621 2805 11655 2839
rect 12357 2805 12391 2839
rect 12909 2805 12943 2839
rect 14749 2805 14783 2839
rect 15485 2805 15519 2839
rect 16037 2805 16071 2839
rect 16773 2805 16807 2839
rect 17509 2805 17543 2839
rect 18061 2805 18095 2839
rect 19993 2805 20027 2839
rect 20729 2805 20763 2839
rect 21189 2805 21223 2839
rect 21925 2805 21959 2839
rect 22661 2805 22695 2839
rect 23213 2805 23247 2839
rect 25053 2805 25087 2839
rect 31493 2805 31527 2839
rect 35357 2805 35391 2839
rect 36093 2805 36127 2839
rect 36645 2805 36679 2839
rect 37381 2805 37415 2839
rect 38117 2805 38151 2839
rect 38669 2805 38703 2839
rect 41061 2805 41095 2839
rect 42441 2805 42475 2839
rect 42993 2805 43027 2839
rect 44833 2805 44867 2839
rect 45661 2805 45695 2839
rect 46305 2805 46339 2839
rect 47593 2805 47627 2839
rect 48145 2805 48179 2839
rect 48789 2805 48823 2839
rect 49341 2805 49375 2839
rect 54585 2805 54619 2839
rect 59645 2805 59679 2839
rect 63049 2805 63083 2839
rect 64889 2805 64923 2839
rect 70041 2805 70075 2839
rect 73353 2805 73387 2839
rect 73905 2805 73939 2839
rect 75745 2805 75779 2839
rect 76481 2805 76515 2839
rect 2329 2601 2363 2635
rect 3065 2601 3099 2635
rect 4537 2601 4571 2635
rect 5181 2601 5215 2635
rect 5641 2601 5675 2635
rect 6745 2601 6779 2635
rect 7481 2601 7515 2635
rect 8217 2601 8251 2635
rect 9597 2601 9631 2635
rect 10057 2601 10091 2635
rect 10793 2601 10827 2635
rect 11897 2601 11931 2635
rect 12633 2601 12667 2635
rect 13369 2601 13403 2635
rect 14473 2601 14507 2635
rect 15945 2601 15979 2635
rect 17049 2601 17083 2635
rect 17785 2601 17819 2635
rect 18521 2601 18555 2635
rect 20361 2601 20395 2635
rect 22937 2601 22971 2635
rect 23673 2601 23707 2635
rect 24961 2601 24995 2635
rect 33977 2601 34011 2635
rect 35817 2601 35851 2635
rect 36553 2601 36587 2635
rect 37657 2601 37691 2635
rect 38393 2601 38427 2635
rect 39129 2601 39163 2635
rect 40601 2601 40635 2635
rect 42625 2601 42659 2635
rect 43361 2601 43395 2635
rect 45201 2601 45235 2635
rect 45937 2601 45971 2635
rect 46673 2601 46707 2635
rect 47777 2601 47811 2635
rect 49249 2601 49283 2635
rect 73537 2601 73571 2635
rect 74273 2601 74307 2635
rect 75009 2601 75043 2635
rect 76113 2601 76147 2635
rect 15117 2533 15151 2567
rect 19533 2533 19567 2567
rect 22293 2533 22327 2567
rect 34989 2533 35023 2567
rect 41429 2533 41463 2567
rect 44189 2533 44223 2567
rect 48605 2533 48639 2567
rect 53573 2533 53607 2567
rect 58817 2533 58851 2567
rect 64705 2533 64739 2567
rect 69857 2533 69891 2567
rect 26157 2465 26191 2499
rect 28733 2465 28767 2499
rect 31033 2465 31067 2499
rect 32413 2465 32447 2499
rect 1685 2397 1719 2431
rect 2145 2397 2179 2431
rect 2881 2397 2915 2431
rect 3893 2397 3927 2431
rect 4353 2397 4387 2431
rect 4997 2397 5031 2431
rect 5825 2397 5859 2431
rect 6561 2397 6595 2431
rect 7297 2397 7331 2431
rect 8033 2397 8067 2431
rect 9413 2397 9447 2431
rect 10241 2397 10275 2431
rect 10977 2397 11011 2431
rect 22109 2397 22143 2431
rect 23581 2397 23615 2431
rect 26433 2397 26467 2431
rect 26985 2397 27019 2431
rect 29009 2397 29043 2431
rect 29561 2397 29595 2431
rect 30297 2397 30331 2431
rect 30757 2397 30791 2431
rect 32137 2397 32171 2431
rect 45845 2397 45879 2431
rect 48421 2397 48455 2431
rect 50445 2397 50479 2431
rect 51181 2397 51215 2431
rect 51917 2397 51951 2431
rect 52745 2397 52779 2431
rect 53757 2397 53791 2431
rect 54217 2397 54251 2431
rect 55321 2397 55355 2431
rect 56333 2397 56367 2431
rect 57069 2397 57103 2431
rect 57897 2397 57931 2431
rect 58633 2397 58667 2431
rect 59369 2397 59403 2431
rect 60749 2397 60783 2431
rect 61485 2397 61519 2431
rect 61945 2397 61979 2431
rect 63049 2397 63083 2431
rect 63785 2397 63819 2431
rect 64521 2397 64555 2431
rect 65625 2397 65659 2431
rect 66361 2397 66395 2431
rect 67097 2397 67131 2431
rect 68201 2397 68235 2431
rect 68937 2397 68971 2431
rect 69673 2397 69707 2431
rect 70777 2397 70811 2431
rect 71513 2397 71547 2431
rect 72249 2397 72283 2431
rect 73353 2397 73387 2431
rect 74089 2397 74123 2431
rect 74825 2397 74859 2431
rect 75929 2397 75963 2431
rect 76665 2397 76699 2431
rect 77401 2397 77435 2431
rect 11805 2329 11839 2363
rect 12541 2329 12575 2363
rect 13277 2329 13311 2363
rect 14565 2329 14599 2363
rect 15301 2329 15335 2363
rect 16037 2329 16071 2363
rect 16957 2329 16991 2363
rect 17693 2329 17727 2363
rect 18429 2329 18463 2363
rect 19717 2329 19751 2363
rect 20453 2329 20487 2363
rect 21189 2329 21223 2363
rect 22845 2329 22879 2363
rect 25053 2329 25087 2363
rect 33885 2329 33919 2363
rect 35173 2329 35207 2363
rect 35909 2329 35943 2363
rect 36645 2329 36679 2363
rect 37565 2329 37599 2363
rect 38301 2329 38335 2363
rect 39037 2329 39071 2363
rect 39957 2329 39991 2363
rect 40509 2329 40543 2363
rect 41245 2329 41279 2363
rect 42533 2329 42567 2363
rect 43269 2329 43303 2363
rect 44005 2329 44039 2363
rect 45109 2329 45143 2363
rect 46581 2329 46615 2363
rect 47685 2329 47719 2363
rect 49157 2329 49191 2363
rect 21097 2261 21131 2295
rect 50261 2261 50295 2295
rect 50997 2261 51031 2295
rect 51733 2261 51767 2295
rect 52929 2261 52963 2295
rect 54401 2261 54435 2295
rect 55505 2261 55539 2295
rect 56149 2261 56183 2295
rect 56885 2261 56919 2295
rect 58081 2261 58115 2295
rect 59553 2261 59587 2295
rect 60565 2261 60599 2295
rect 61301 2261 61335 2295
rect 62129 2261 62163 2295
rect 63233 2261 63267 2295
rect 63969 2261 64003 2295
rect 65809 2261 65843 2295
rect 66545 2261 66579 2295
rect 67281 2261 67315 2295
rect 68385 2261 68419 2295
rect 69121 2261 69155 2295
rect 70961 2261 70995 2295
rect 71697 2261 71731 2295
rect 72433 2261 72467 2295
rect 76849 2261 76883 2295
rect 77585 2261 77619 2295
<< metal1 >>
rect 1104 77818 78844 77840
rect 1104 77766 4214 77818
rect 4266 77766 4278 77818
rect 4330 77766 4342 77818
rect 4394 77766 4406 77818
rect 4458 77766 4470 77818
rect 4522 77766 34934 77818
rect 34986 77766 34998 77818
rect 35050 77766 35062 77818
rect 35114 77766 35126 77818
rect 35178 77766 35190 77818
rect 35242 77766 65654 77818
rect 65706 77766 65718 77818
rect 65770 77766 65782 77818
rect 65834 77766 65846 77818
rect 65898 77766 65910 77818
rect 65962 77766 78844 77818
rect 1104 77744 78844 77766
rect 1104 77274 78844 77296
rect 1104 77222 19574 77274
rect 19626 77222 19638 77274
rect 19690 77222 19702 77274
rect 19754 77222 19766 77274
rect 19818 77222 19830 77274
rect 19882 77222 50294 77274
rect 50346 77222 50358 77274
rect 50410 77222 50422 77274
rect 50474 77222 50486 77274
rect 50538 77222 50550 77274
rect 50602 77222 78844 77274
rect 1104 77200 78844 77222
rect 1104 76730 78844 76752
rect 1104 76678 4214 76730
rect 4266 76678 4278 76730
rect 4330 76678 4342 76730
rect 4394 76678 4406 76730
rect 4458 76678 4470 76730
rect 4522 76678 34934 76730
rect 34986 76678 34998 76730
rect 35050 76678 35062 76730
rect 35114 76678 35126 76730
rect 35178 76678 35190 76730
rect 35242 76678 65654 76730
rect 65706 76678 65718 76730
rect 65770 76678 65782 76730
rect 65834 76678 65846 76730
rect 65898 76678 65910 76730
rect 65962 76678 78844 76730
rect 1104 76656 78844 76678
rect 1104 76186 78844 76208
rect 1104 76134 19574 76186
rect 19626 76134 19638 76186
rect 19690 76134 19702 76186
rect 19754 76134 19766 76186
rect 19818 76134 19830 76186
rect 19882 76134 50294 76186
rect 50346 76134 50358 76186
rect 50410 76134 50422 76186
rect 50474 76134 50486 76186
rect 50538 76134 50550 76186
rect 50602 76134 78844 76186
rect 1104 76112 78844 76134
rect 1104 75642 78844 75664
rect 1104 75590 4214 75642
rect 4266 75590 4278 75642
rect 4330 75590 4342 75642
rect 4394 75590 4406 75642
rect 4458 75590 4470 75642
rect 4522 75590 34934 75642
rect 34986 75590 34998 75642
rect 35050 75590 35062 75642
rect 35114 75590 35126 75642
rect 35178 75590 35190 75642
rect 35242 75590 65654 75642
rect 65706 75590 65718 75642
rect 65770 75590 65782 75642
rect 65834 75590 65846 75642
rect 65898 75590 65910 75642
rect 65962 75590 78844 75642
rect 1104 75568 78844 75590
rect 1670 75324 1676 75336
rect 1631 75296 1676 75324
rect 1670 75284 1676 75296
rect 1728 75324 1734 75336
rect 2133 75327 2191 75333
rect 2133 75324 2145 75327
rect 1728 75296 2145 75324
rect 1728 75284 1734 75296
rect 2133 75293 2145 75296
rect 2179 75293 2191 75327
rect 77849 75327 77907 75333
rect 77849 75324 77861 75327
rect 2133 75287 2191 75293
rect 77312 75296 77861 75324
rect 1486 75188 1492 75200
rect 1447 75160 1492 75188
rect 1486 75148 1492 75160
rect 1544 75148 1550 75200
rect 76558 75148 76564 75200
rect 76616 75188 76622 75200
rect 77312 75197 77340 75296
rect 77849 75293 77861 75296
rect 77895 75293 77907 75327
rect 77849 75287 77907 75293
rect 77297 75191 77355 75197
rect 77297 75188 77309 75191
rect 76616 75160 77309 75188
rect 76616 75148 76622 75160
rect 77297 75157 77309 75160
rect 77343 75157 77355 75191
rect 78030 75188 78036 75200
rect 77991 75160 78036 75188
rect 77297 75151 77355 75157
rect 78030 75148 78036 75160
rect 78088 75148 78094 75200
rect 1104 75098 78844 75120
rect 1104 75046 19574 75098
rect 19626 75046 19638 75098
rect 19690 75046 19702 75098
rect 19754 75046 19766 75098
rect 19818 75046 19830 75098
rect 19882 75046 50294 75098
rect 50346 75046 50358 75098
rect 50410 75046 50422 75098
rect 50474 75046 50486 75098
rect 50538 75046 50550 75098
rect 50602 75046 78844 75098
rect 1104 75024 78844 75046
rect 1394 74848 1400 74860
rect 1355 74820 1400 74848
rect 1394 74808 1400 74820
rect 1452 74808 1458 74860
rect 77849 74851 77907 74857
rect 77849 74817 77861 74851
rect 77895 74848 77907 74851
rect 78122 74848 78128 74860
rect 77895 74820 78128 74848
rect 77895 74817 77907 74820
rect 77849 74811 77907 74817
rect 78122 74808 78128 74820
rect 78180 74808 78186 74860
rect 77570 74672 77576 74724
rect 77628 74712 77634 74724
rect 77665 74715 77723 74721
rect 77665 74712 77677 74715
rect 77628 74684 77677 74712
rect 77628 74672 77634 74684
rect 77665 74681 77677 74684
rect 77711 74681 77723 74715
rect 77665 74675 77723 74681
rect 1581 74647 1639 74653
rect 1581 74613 1593 74647
rect 1627 74644 1639 74647
rect 2406 74644 2412 74656
rect 1627 74616 2412 74644
rect 1627 74613 1639 74616
rect 1581 74607 1639 74613
rect 2406 74604 2412 74616
rect 2464 74604 2470 74656
rect 1104 74554 78844 74576
rect 1104 74502 4214 74554
rect 4266 74502 4278 74554
rect 4330 74502 4342 74554
rect 4394 74502 4406 74554
rect 4458 74502 4470 74554
rect 4522 74502 34934 74554
rect 34986 74502 34998 74554
rect 35050 74502 35062 74554
rect 35114 74502 35126 74554
rect 35178 74502 35190 74554
rect 35242 74502 65654 74554
rect 65706 74502 65718 74554
rect 65770 74502 65782 74554
rect 65834 74502 65846 74554
rect 65898 74502 65910 74554
rect 65962 74502 78844 74554
rect 1104 74480 78844 74502
rect 1394 74372 1400 74384
rect 1355 74344 1400 74372
rect 1394 74332 1400 74344
rect 1452 74332 1458 74384
rect 78122 74372 78128 74384
rect 78083 74344 78128 74372
rect 78122 74332 78128 74344
rect 78180 74332 78186 74384
rect 1104 74010 78844 74032
rect 1104 73958 19574 74010
rect 19626 73958 19638 74010
rect 19690 73958 19702 74010
rect 19754 73958 19766 74010
rect 19818 73958 19830 74010
rect 19882 73958 50294 74010
rect 50346 73958 50358 74010
rect 50410 73958 50422 74010
rect 50474 73958 50486 74010
rect 50538 73958 50550 74010
rect 50602 73958 78844 74010
rect 1104 73936 78844 73958
rect 1673 73763 1731 73769
rect 1673 73729 1685 73763
rect 1719 73760 1731 73763
rect 77665 73763 77723 73769
rect 77665 73760 77677 73763
rect 1719 73732 2268 73760
rect 1719 73729 1731 73732
rect 1673 73723 1731 73729
rect 1486 73624 1492 73636
rect 1447 73596 1492 73624
rect 1486 73584 1492 73596
rect 1544 73584 1550 73636
rect 2240 73565 2268 73732
rect 77128 73732 77677 73760
rect 2225 73559 2283 73565
rect 2225 73525 2237 73559
rect 2271 73556 2283 73559
rect 2682 73556 2688 73568
rect 2271 73528 2688 73556
rect 2271 73525 2283 73528
rect 2225 73519 2283 73525
rect 2682 73516 2688 73528
rect 2740 73516 2746 73568
rect 77018 73516 77024 73568
rect 77076 73556 77082 73568
rect 77128 73565 77156 73732
rect 77665 73729 77677 73732
rect 77711 73729 77723 73763
rect 77665 73723 77723 73729
rect 77846 73624 77852 73636
rect 77807 73596 77852 73624
rect 77846 73584 77852 73596
rect 77904 73584 77910 73636
rect 77113 73559 77171 73565
rect 77113 73556 77125 73559
rect 77076 73528 77125 73556
rect 77076 73516 77082 73528
rect 77113 73525 77125 73528
rect 77159 73525 77171 73559
rect 77113 73519 77171 73525
rect 1104 73466 78844 73488
rect 1104 73414 4214 73466
rect 4266 73414 4278 73466
rect 4330 73414 4342 73466
rect 4394 73414 4406 73466
rect 4458 73414 4470 73466
rect 4522 73414 34934 73466
rect 34986 73414 34998 73466
rect 35050 73414 35062 73466
rect 35114 73414 35126 73466
rect 35178 73414 35190 73466
rect 35242 73414 65654 73466
rect 65706 73414 65718 73466
rect 65770 73414 65782 73466
rect 65834 73414 65846 73466
rect 65898 73414 65910 73466
rect 65962 73414 78844 73466
rect 1104 73392 78844 73414
rect 1673 73151 1731 73157
rect 1673 73117 1685 73151
rect 1719 73148 1731 73151
rect 1719 73120 2268 73148
rect 1719 73117 1731 73120
rect 1673 73111 1731 73117
rect 1486 73012 1492 73024
rect 1447 72984 1492 73012
rect 1486 72972 1492 72984
rect 1544 72972 1550 73024
rect 2240 73021 2268 73120
rect 76190 73108 76196 73160
rect 76248 73148 76254 73160
rect 77849 73151 77907 73157
rect 77849 73148 77861 73151
rect 76248 73120 77861 73148
rect 76248 73108 76254 73120
rect 77849 73117 77861 73120
rect 77895 73117 77907 73151
rect 77849 73111 77907 73117
rect 2225 73015 2283 73021
rect 2225 72981 2237 73015
rect 2271 73012 2283 73015
rect 2314 73012 2320 73024
rect 2271 72984 2320 73012
rect 2271 72981 2283 72984
rect 2225 72975 2283 72981
rect 2314 72972 2320 72984
rect 2372 72972 2378 73024
rect 78030 73012 78036 73024
rect 77991 72984 78036 73012
rect 78030 72972 78036 72984
rect 78088 72972 78094 73024
rect 1104 72922 78844 72944
rect 1104 72870 19574 72922
rect 19626 72870 19638 72922
rect 19690 72870 19702 72922
rect 19754 72870 19766 72922
rect 19818 72870 19830 72922
rect 19882 72870 50294 72922
rect 50346 72870 50358 72922
rect 50410 72870 50422 72922
rect 50474 72870 50486 72922
rect 50538 72870 50550 72922
rect 50602 72870 78844 72922
rect 1104 72848 78844 72870
rect 1673 72675 1731 72681
rect 1673 72641 1685 72675
rect 1719 72672 1731 72675
rect 1719 72644 2268 72672
rect 1719 72641 1731 72644
rect 1673 72635 1731 72641
rect 1486 72468 1492 72480
rect 1447 72440 1492 72468
rect 1486 72428 1492 72440
rect 1544 72428 1550 72480
rect 2240 72477 2268 72644
rect 76098 72632 76104 72684
rect 76156 72672 76162 72684
rect 77665 72675 77723 72681
rect 77665 72672 77677 72675
rect 76156 72644 77677 72672
rect 76156 72632 76162 72644
rect 77665 72641 77677 72644
rect 77711 72641 77723 72675
rect 77665 72635 77723 72641
rect 2225 72471 2283 72477
rect 2225 72437 2237 72471
rect 2271 72468 2283 72471
rect 2406 72468 2412 72480
rect 2271 72440 2412 72468
rect 2271 72437 2283 72440
rect 2225 72431 2283 72437
rect 2406 72428 2412 72440
rect 2464 72428 2470 72480
rect 77846 72468 77852 72480
rect 77807 72440 77852 72468
rect 77846 72428 77852 72440
rect 77904 72428 77910 72480
rect 1104 72378 78844 72400
rect 1104 72326 4214 72378
rect 4266 72326 4278 72378
rect 4330 72326 4342 72378
rect 4394 72326 4406 72378
rect 4458 72326 4470 72378
rect 4522 72326 34934 72378
rect 34986 72326 34998 72378
rect 35050 72326 35062 72378
rect 35114 72326 35126 72378
rect 35178 72326 35190 72378
rect 35242 72326 65654 72378
rect 65706 72326 65718 72378
rect 65770 72326 65782 72378
rect 65834 72326 65846 72378
rect 65898 72326 65910 72378
rect 65962 72326 78844 72378
rect 1104 72304 78844 72326
rect 1673 72063 1731 72069
rect 1673 72029 1685 72063
rect 1719 72060 1731 72063
rect 1719 72032 2268 72060
rect 1719 72029 1731 72032
rect 1673 72023 1731 72029
rect 2240 71936 2268 72032
rect 75914 72020 75920 72072
rect 75972 72060 75978 72072
rect 77849 72063 77907 72069
rect 77849 72060 77861 72063
rect 75972 72032 77861 72060
rect 75972 72020 75978 72032
rect 77849 72029 77861 72032
rect 77895 72029 77907 72063
rect 77849 72023 77907 72029
rect 1486 71924 1492 71936
rect 1447 71896 1492 71924
rect 1486 71884 1492 71896
rect 1544 71884 1550 71936
rect 2222 71924 2228 71936
rect 2183 71896 2228 71924
rect 2222 71884 2228 71896
rect 2280 71884 2286 71936
rect 78030 71924 78036 71936
rect 77991 71896 78036 71924
rect 78030 71884 78036 71896
rect 78088 71884 78094 71936
rect 1104 71834 78844 71856
rect 1104 71782 19574 71834
rect 19626 71782 19638 71834
rect 19690 71782 19702 71834
rect 19754 71782 19766 71834
rect 19818 71782 19830 71834
rect 19882 71782 50294 71834
rect 50346 71782 50358 71834
rect 50410 71782 50422 71834
rect 50474 71782 50486 71834
rect 50538 71782 50550 71834
rect 50602 71782 78844 71834
rect 1104 71760 78844 71782
rect 76190 71720 76196 71732
rect 76151 71692 76196 71720
rect 76190 71680 76196 71692
rect 76248 71680 76254 71732
rect 72605 71587 72663 71593
rect 72605 71553 72617 71587
rect 72651 71584 72663 71587
rect 73433 71587 73491 71593
rect 73433 71584 73445 71587
rect 72651 71556 73445 71584
rect 72651 71553 72663 71556
rect 72605 71547 72663 71553
rect 73433 71553 73445 71556
rect 73479 71584 73491 71587
rect 76009 71587 76067 71593
rect 76009 71584 76021 71587
rect 73479 71556 76021 71584
rect 73479 71553 73491 71556
rect 73433 71547 73491 71553
rect 76009 71553 76021 71556
rect 76055 71584 76067 71587
rect 76282 71584 76288 71596
rect 76055 71556 76288 71584
rect 76055 71553 76067 71556
rect 76009 71547 76067 71553
rect 76282 71544 76288 71556
rect 76340 71544 76346 71596
rect 2314 71340 2320 71392
rect 2372 71380 2378 71392
rect 72421 71383 72479 71389
rect 72421 71380 72433 71383
rect 2372 71352 72433 71380
rect 2372 71340 2378 71352
rect 72421 71349 72433 71352
rect 72467 71349 72479 71383
rect 72421 71343 72479 71349
rect 76282 71340 76288 71392
rect 76340 71380 76346 71392
rect 76653 71383 76711 71389
rect 76653 71380 76665 71383
rect 76340 71352 76665 71380
rect 76340 71340 76346 71352
rect 76653 71349 76665 71352
rect 76699 71349 76711 71383
rect 76653 71343 76711 71349
rect 1104 71290 78844 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 34934 71290
rect 34986 71238 34998 71290
rect 35050 71238 35062 71290
rect 35114 71238 35126 71290
rect 35178 71238 35190 71290
rect 35242 71238 65654 71290
rect 65706 71238 65718 71290
rect 65770 71238 65782 71290
rect 65834 71238 65846 71290
rect 65898 71238 65910 71290
rect 65962 71238 78844 71290
rect 1104 71216 78844 71238
rect 76098 71176 76104 71188
rect 76059 71148 76104 71176
rect 76098 71136 76104 71148
rect 76156 71136 76162 71188
rect 1673 70975 1731 70981
rect 1673 70941 1685 70975
rect 1719 70972 1731 70975
rect 72053 70975 72111 70981
rect 1719 70944 2268 70972
rect 1719 70941 1731 70944
rect 1673 70935 1731 70941
rect 1486 70836 1492 70848
rect 1447 70808 1492 70836
rect 1486 70796 1492 70808
rect 1544 70796 1550 70848
rect 2240 70845 2268 70944
rect 72053 70941 72065 70975
rect 72099 70972 72111 70975
rect 72605 70975 72663 70981
rect 72605 70972 72617 70975
rect 72099 70944 72617 70972
rect 72099 70941 72111 70944
rect 72053 70935 72111 70941
rect 72605 70941 72617 70944
rect 72651 70972 72663 70975
rect 75917 70975 75975 70981
rect 75917 70972 75929 70975
rect 72651 70944 75929 70972
rect 72651 70941 72663 70944
rect 72605 70935 72663 70941
rect 75917 70941 75929 70944
rect 75963 70972 75975 70975
rect 76006 70972 76012 70984
rect 75963 70944 76012 70972
rect 75963 70941 75975 70944
rect 75917 70935 75975 70941
rect 76006 70932 76012 70944
rect 76064 70972 76070 70984
rect 76561 70975 76619 70981
rect 76561 70972 76573 70975
rect 76064 70944 76573 70972
rect 76064 70932 76070 70944
rect 76561 70941 76573 70944
rect 76607 70941 76619 70975
rect 76561 70935 76619 70941
rect 77849 70975 77907 70981
rect 77849 70941 77861 70975
rect 77895 70941 77907 70975
rect 77849 70935 77907 70941
rect 2406 70864 2412 70916
rect 2464 70904 2470 70916
rect 2464 70876 64874 70904
rect 2464 70864 2470 70876
rect 2225 70839 2283 70845
rect 2225 70805 2237 70839
rect 2271 70836 2283 70839
rect 2314 70836 2320 70848
rect 2271 70808 2320 70836
rect 2271 70805 2283 70808
rect 2225 70799 2283 70805
rect 2314 70796 2320 70808
rect 2372 70796 2378 70848
rect 64846 70836 64874 70876
rect 75822 70864 75828 70916
rect 75880 70904 75886 70916
rect 77864 70904 77892 70935
rect 75880 70876 77892 70904
rect 75880 70864 75886 70876
rect 71869 70839 71927 70845
rect 71869 70836 71881 70839
rect 64846 70808 71881 70836
rect 71869 70805 71881 70808
rect 71915 70805 71927 70839
rect 78030 70836 78036 70848
rect 77991 70808 78036 70836
rect 71869 70799 71927 70805
rect 78030 70796 78036 70808
rect 78088 70796 78094 70848
rect 1104 70746 78844 70768
rect 1104 70694 19574 70746
rect 19626 70694 19638 70746
rect 19690 70694 19702 70746
rect 19754 70694 19766 70746
rect 19818 70694 19830 70746
rect 19882 70694 50294 70746
rect 50346 70694 50358 70746
rect 50410 70694 50422 70746
rect 50474 70694 50486 70746
rect 50538 70694 50550 70746
rect 50602 70694 78844 70746
rect 1104 70672 78844 70694
rect 71225 70635 71283 70641
rect 71225 70632 71237 70635
rect 64846 70604 71237 70632
rect 2222 70524 2228 70576
rect 2280 70564 2286 70576
rect 64846 70564 64874 70604
rect 71225 70601 71237 70604
rect 71271 70601 71283 70635
rect 71225 70595 71283 70601
rect 74813 70635 74871 70641
rect 74813 70601 74825 70635
rect 74859 70632 74871 70635
rect 75914 70632 75920 70644
rect 74859 70604 75920 70632
rect 74859 70601 74871 70604
rect 74813 70595 74871 70601
rect 75914 70592 75920 70604
rect 75972 70592 75978 70644
rect 2280 70536 64874 70564
rect 2280 70524 2286 70536
rect 1673 70499 1731 70505
rect 1673 70465 1685 70499
rect 1719 70496 1731 70499
rect 71409 70499 71467 70505
rect 1719 70468 2268 70496
rect 1719 70465 1731 70468
rect 1673 70459 1731 70465
rect 2240 70440 2268 70468
rect 71409 70465 71421 70499
rect 71455 70496 71467 70499
rect 71961 70499 72019 70505
rect 71961 70496 71973 70499
rect 71455 70468 71973 70496
rect 71455 70465 71467 70468
rect 71409 70459 71467 70465
rect 71961 70465 71973 70468
rect 72007 70496 72019 70499
rect 74629 70499 74687 70505
rect 74629 70496 74641 70499
rect 72007 70468 74641 70496
rect 72007 70465 72019 70468
rect 71961 70459 72019 70465
rect 74629 70465 74641 70468
rect 74675 70496 74687 70499
rect 74994 70496 75000 70508
rect 74675 70468 75000 70496
rect 74675 70465 74687 70468
rect 74629 70459 74687 70465
rect 74994 70456 75000 70468
rect 75052 70496 75058 70508
rect 75273 70499 75331 70505
rect 75273 70496 75285 70499
rect 75052 70468 75285 70496
rect 75052 70456 75058 70468
rect 75273 70465 75285 70468
rect 75319 70465 75331 70499
rect 75273 70459 75331 70465
rect 77665 70499 77723 70505
rect 77665 70465 77677 70499
rect 77711 70465 77723 70499
rect 77665 70459 77723 70465
rect 2222 70428 2228 70440
rect 2183 70400 2228 70428
rect 2222 70388 2228 70400
rect 2280 70388 2286 70440
rect 73338 70388 73344 70440
rect 73396 70428 73402 70440
rect 77680 70428 77708 70459
rect 73396 70400 77708 70428
rect 73396 70388 73402 70400
rect 1486 70292 1492 70304
rect 1447 70264 1492 70292
rect 1486 70252 1492 70264
rect 1544 70252 1550 70304
rect 77846 70292 77852 70304
rect 77807 70264 77852 70292
rect 77846 70252 77852 70264
rect 77904 70252 77910 70304
rect 1104 70202 78844 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 34934 70202
rect 34986 70150 34998 70202
rect 35050 70150 35062 70202
rect 35114 70150 35126 70202
rect 35178 70150 35190 70202
rect 35242 70150 65654 70202
rect 65706 70150 65718 70202
rect 65770 70150 65782 70202
rect 65834 70150 65846 70202
rect 65898 70150 65910 70202
rect 65962 70150 78844 70202
rect 1104 70128 78844 70150
rect 74077 70091 74135 70097
rect 74077 70057 74089 70091
rect 74123 70088 74135 70091
rect 75822 70088 75828 70100
rect 74123 70060 75828 70088
rect 74123 70057 74135 70060
rect 74077 70051 74135 70057
rect 75822 70048 75828 70060
rect 75880 70048 75886 70100
rect 1394 69884 1400 69896
rect 1355 69856 1400 69884
rect 1394 69844 1400 69856
rect 1452 69884 1458 69896
rect 2133 69887 2191 69893
rect 2133 69884 2145 69887
rect 1452 69856 2145 69884
rect 1452 69844 1458 69856
rect 2133 69853 2145 69856
rect 2179 69853 2191 69887
rect 2133 69847 2191 69853
rect 71041 69887 71099 69893
rect 71041 69853 71053 69887
rect 71087 69884 71099 69887
rect 71593 69887 71651 69893
rect 71593 69884 71605 69887
rect 71087 69856 71605 69884
rect 71087 69853 71099 69856
rect 71041 69847 71099 69853
rect 71593 69853 71605 69856
rect 71639 69884 71651 69887
rect 73893 69887 73951 69893
rect 73893 69884 73905 69887
rect 71639 69856 73905 69884
rect 71639 69853 71651 69856
rect 71593 69847 71651 69853
rect 73893 69853 73905 69856
rect 73939 69884 73951 69887
rect 77481 69887 77539 69893
rect 73939 69856 74304 69884
rect 73939 69853 73951 69856
rect 73893 69847 73951 69853
rect 2314 69776 2320 69828
rect 2372 69816 2378 69828
rect 2372 69788 64874 69816
rect 2372 69776 2378 69788
rect 1581 69751 1639 69757
rect 1581 69717 1593 69751
rect 1627 69748 1639 69751
rect 1762 69748 1768 69760
rect 1627 69720 1768 69748
rect 1627 69717 1639 69720
rect 1581 69711 1639 69717
rect 1762 69708 1768 69720
rect 1820 69708 1826 69760
rect 64846 69748 64874 69788
rect 74276 69760 74304 69856
rect 77481 69853 77493 69887
rect 77527 69884 77539 69887
rect 78122 69884 78128 69896
rect 77527 69856 78128 69884
rect 77527 69853 77539 69856
rect 77481 69847 77539 69853
rect 78122 69844 78128 69856
rect 78180 69844 78186 69896
rect 70857 69751 70915 69757
rect 70857 69748 70869 69751
rect 64846 69720 70869 69748
rect 70857 69717 70869 69720
rect 70903 69717 70915 69751
rect 70857 69711 70915 69717
rect 74258 69708 74264 69760
rect 74316 69748 74322 69760
rect 74537 69751 74595 69757
rect 74537 69748 74549 69751
rect 74316 69720 74549 69748
rect 74316 69708 74322 69720
rect 74537 69717 74549 69720
rect 74583 69717 74595 69751
rect 77938 69748 77944 69760
rect 77899 69720 77944 69748
rect 74537 69711 74595 69717
rect 77938 69708 77944 69720
rect 77996 69708 78002 69760
rect 1104 69658 78844 69680
rect 1104 69606 19574 69658
rect 19626 69606 19638 69658
rect 19690 69606 19702 69658
rect 19754 69606 19766 69658
rect 19818 69606 19830 69658
rect 19882 69606 50294 69658
rect 50346 69606 50358 69658
rect 50410 69606 50422 69658
rect 50474 69606 50486 69658
rect 50538 69606 50550 69658
rect 50602 69606 78844 69658
rect 1104 69584 78844 69606
rect 65978 69504 65984 69556
rect 66036 69544 66042 69556
rect 77938 69544 77944 69556
rect 66036 69516 77944 69544
rect 66036 69504 66042 69516
rect 77938 69504 77944 69516
rect 77996 69504 78002 69556
rect 1394 69408 1400 69420
rect 1355 69380 1400 69408
rect 1394 69368 1400 69380
rect 1452 69408 1458 69420
rect 2133 69411 2191 69417
rect 2133 69408 2145 69411
rect 1452 69380 2145 69408
rect 1452 69368 1458 69380
rect 2133 69377 2145 69380
rect 2179 69377 2191 69411
rect 2133 69371 2191 69377
rect 77297 69411 77355 69417
rect 77297 69377 77309 69411
rect 77343 69408 77355 69411
rect 77938 69408 77944 69420
rect 77343 69380 77944 69408
rect 77343 69377 77355 69380
rect 77297 69371 77355 69377
rect 77938 69368 77944 69380
rect 77996 69368 78002 69420
rect 1581 69207 1639 69213
rect 1581 69173 1593 69207
rect 1627 69204 1639 69207
rect 1670 69204 1676 69216
rect 1627 69176 1676 69204
rect 1627 69173 1639 69176
rect 1581 69167 1639 69173
rect 1670 69164 1676 69176
rect 1728 69164 1734 69216
rect 76650 69164 76656 69216
rect 76708 69204 76714 69216
rect 77757 69207 77815 69213
rect 77757 69204 77769 69207
rect 76708 69176 77769 69204
rect 76708 69164 76714 69176
rect 77757 69173 77769 69176
rect 77803 69173 77815 69207
rect 77757 69167 77815 69173
rect 1104 69114 78844 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 34934 69114
rect 34986 69062 34998 69114
rect 35050 69062 35062 69114
rect 35114 69062 35126 69114
rect 35178 69062 35190 69114
rect 35242 69062 65654 69114
rect 65706 69062 65718 69114
rect 65770 69062 65782 69114
rect 65834 69062 65846 69114
rect 65898 69062 65910 69114
rect 65962 69062 78844 69114
rect 1104 69040 78844 69062
rect 73338 69000 73344 69012
rect 73299 68972 73344 69000
rect 73338 68960 73344 68972
rect 73396 68960 73402 69012
rect 70121 68799 70179 68805
rect 70121 68765 70133 68799
rect 70167 68796 70179 68799
rect 70857 68799 70915 68805
rect 70857 68796 70869 68799
rect 70167 68768 70869 68796
rect 70167 68765 70179 68768
rect 70121 68759 70179 68765
rect 70857 68765 70869 68768
rect 70903 68796 70915 68799
rect 73157 68799 73215 68805
rect 73157 68796 73169 68799
rect 70903 68768 73169 68796
rect 70903 68765 70915 68768
rect 70857 68759 70915 68765
rect 73157 68765 73169 68768
rect 73203 68796 73215 68799
rect 73203 68768 73568 68796
rect 73203 68765 73215 68768
rect 73157 68759 73215 68765
rect 73540 68672 73568 68768
rect 1394 68660 1400 68672
rect 1355 68632 1400 68660
rect 1394 68620 1400 68632
rect 1452 68620 1458 68672
rect 2222 68620 2228 68672
rect 2280 68660 2286 68672
rect 69937 68663 69995 68669
rect 69937 68660 69949 68663
rect 2280 68632 69949 68660
rect 2280 68620 2286 68632
rect 69937 68629 69949 68632
rect 69983 68629 69995 68663
rect 69937 68623 69995 68629
rect 73522 68620 73528 68672
rect 73580 68660 73586 68672
rect 73801 68663 73859 68669
rect 73801 68660 73813 68663
rect 73580 68632 73813 68660
rect 73580 68620 73586 68632
rect 73801 68629 73813 68632
rect 73847 68629 73859 68663
rect 73801 68623 73859 68629
rect 77938 68620 77944 68672
rect 77996 68660 78002 68672
rect 78033 68663 78091 68669
rect 78033 68660 78045 68663
rect 77996 68632 78045 68660
rect 77996 68620 78002 68632
rect 78033 68629 78045 68632
rect 78079 68629 78091 68663
rect 78033 68623 78091 68629
rect 1104 68570 78844 68592
rect 1104 68518 19574 68570
rect 19626 68518 19638 68570
rect 19690 68518 19702 68570
rect 19754 68518 19766 68570
rect 19818 68518 19830 68570
rect 19882 68518 50294 68570
rect 50346 68518 50358 68570
rect 50410 68518 50422 68570
rect 50474 68518 50486 68570
rect 50538 68518 50550 68570
rect 50602 68518 78844 68570
rect 1104 68496 78844 68518
rect 1394 68320 1400 68332
rect 1355 68292 1400 68320
rect 1394 68280 1400 68292
rect 1452 68280 1458 68332
rect 77938 68320 77944 68332
rect 77899 68292 77944 68320
rect 77938 68280 77944 68292
rect 77996 68280 78002 68332
rect 1581 68119 1639 68125
rect 1581 68085 1593 68119
rect 1627 68116 1639 68119
rect 66162 68116 66168 68128
rect 1627 68088 66168 68116
rect 1627 68085 1639 68088
rect 1581 68079 1639 68085
rect 66162 68076 66168 68088
rect 66220 68076 66226 68128
rect 75178 68076 75184 68128
rect 75236 68116 75242 68128
rect 77757 68119 77815 68125
rect 77757 68116 77769 68119
rect 75236 68088 77769 68116
rect 75236 68076 75242 68088
rect 77757 68085 77769 68088
rect 77803 68085 77815 68119
rect 77757 68079 77815 68085
rect 1104 68026 78844 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 34934 68026
rect 34986 67974 34998 68026
rect 35050 67974 35062 68026
rect 35114 67974 35126 68026
rect 35178 67974 35190 68026
rect 35242 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 78844 68026
rect 1104 67952 78844 67974
rect 1581 67847 1639 67853
rect 1581 67813 1593 67847
rect 1627 67844 1639 67847
rect 1854 67844 1860 67856
rect 1627 67816 1860 67844
rect 1627 67813 1639 67816
rect 1581 67807 1639 67813
rect 1854 67804 1860 67816
rect 1912 67804 1918 67856
rect 66990 67804 66996 67856
rect 67048 67844 67054 67856
rect 77941 67847 77999 67853
rect 77941 67844 77953 67847
rect 67048 67816 77953 67844
rect 67048 67804 67054 67816
rect 77941 67813 77953 67816
rect 77987 67813 77999 67847
rect 77941 67807 77999 67813
rect 1394 67708 1400 67720
rect 1355 67680 1400 67708
rect 1394 67668 1400 67680
rect 1452 67708 1458 67720
rect 2133 67711 2191 67717
rect 2133 67708 2145 67711
rect 1452 67680 2145 67708
rect 1452 67668 1458 67680
rect 2133 67677 2145 67680
rect 2179 67677 2191 67711
rect 2133 67671 2191 67677
rect 77481 67711 77539 67717
rect 77481 67677 77493 67711
rect 77527 67708 77539 67711
rect 78122 67708 78128 67720
rect 77527 67680 78128 67708
rect 77527 67677 77539 67680
rect 77481 67671 77539 67677
rect 78122 67668 78128 67680
rect 78180 67668 78186 67720
rect 1104 67482 78844 67504
rect 1104 67430 19574 67482
rect 19626 67430 19638 67482
rect 19690 67430 19702 67482
rect 19754 67430 19766 67482
rect 19818 67430 19830 67482
rect 19882 67430 50294 67482
rect 50346 67430 50358 67482
rect 50410 67430 50422 67482
rect 50474 67430 50486 67482
rect 50538 67430 50550 67482
rect 50602 67430 78844 67482
rect 1104 67408 78844 67430
rect 1394 67232 1400 67244
rect 1355 67204 1400 67232
rect 1394 67192 1400 67204
rect 1452 67232 1458 67244
rect 2133 67235 2191 67241
rect 2133 67232 2145 67235
rect 1452 67204 2145 67232
rect 1452 67192 1458 67204
rect 2133 67201 2145 67204
rect 2179 67201 2191 67235
rect 2133 67195 2191 67201
rect 77297 67235 77355 67241
rect 77297 67201 77309 67235
rect 77343 67232 77355 67235
rect 77938 67232 77944 67244
rect 77343 67204 77944 67232
rect 77343 67201 77355 67204
rect 77297 67195 77355 67201
rect 77938 67192 77944 67204
rect 77996 67192 78002 67244
rect 72326 67056 72332 67108
rect 72384 67096 72390 67108
rect 77757 67099 77815 67105
rect 77757 67096 77769 67099
rect 72384 67068 77769 67096
rect 72384 67056 72390 67068
rect 77757 67065 77769 67068
rect 77803 67065 77815 67099
rect 77757 67059 77815 67065
rect 1578 67028 1584 67040
rect 1539 67000 1584 67028
rect 1578 66988 1584 67000
rect 1636 66988 1642 67040
rect 1104 66938 78844 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 78844 66938
rect 1104 66864 78844 66886
rect 1578 66784 1584 66836
rect 1636 66824 1642 66836
rect 63126 66824 63132 66836
rect 1636 66796 63132 66824
rect 1636 66784 1642 66796
rect 63126 66784 63132 66796
rect 63184 66784 63190 66836
rect 1394 66620 1400 66632
rect 1355 66592 1400 66620
rect 1394 66580 1400 66592
rect 1452 66620 1458 66632
rect 2133 66623 2191 66629
rect 2133 66620 2145 66623
rect 1452 66592 2145 66620
rect 1452 66580 1458 66592
rect 2133 66589 2145 66592
rect 2179 66589 2191 66623
rect 2133 66583 2191 66589
rect 77481 66623 77539 66629
rect 77481 66589 77493 66623
rect 77527 66620 77539 66623
rect 78122 66620 78128 66632
rect 77527 66592 78128 66620
rect 77527 66589 77539 66592
rect 77481 66583 77539 66589
rect 78122 66580 78128 66592
rect 78180 66580 78186 66632
rect 1578 66484 1584 66496
rect 1539 66456 1584 66484
rect 1578 66444 1584 66456
rect 1636 66444 1642 66496
rect 77938 66484 77944 66496
rect 77899 66456 77944 66484
rect 77938 66444 77944 66456
rect 77996 66444 78002 66496
rect 1104 66394 78844 66416
rect 1104 66342 19574 66394
rect 19626 66342 19638 66394
rect 19690 66342 19702 66394
rect 19754 66342 19766 66394
rect 19818 66342 19830 66394
rect 19882 66342 50294 66394
rect 50346 66342 50358 66394
rect 50410 66342 50422 66394
rect 50474 66342 50486 66394
rect 50538 66342 50550 66394
rect 50602 66342 78844 66394
rect 1104 66320 78844 66342
rect 66070 66240 66076 66292
rect 66128 66280 66134 66292
rect 77938 66280 77944 66292
rect 66128 66252 77944 66280
rect 66128 66240 66134 66252
rect 77938 66240 77944 66252
rect 77996 66240 78002 66292
rect 1394 65940 1400 65952
rect 1355 65912 1400 65940
rect 1394 65900 1400 65912
rect 1452 65900 1458 65952
rect 1104 65850 78844 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 78844 65850
rect 1104 65776 78844 65798
rect 1394 65532 1400 65544
rect 1355 65504 1400 65532
rect 1394 65492 1400 65504
rect 1452 65492 1458 65544
rect 77481 65535 77539 65541
rect 77481 65501 77493 65535
rect 77527 65532 77539 65535
rect 78122 65532 78128 65544
rect 77527 65504 78128 65532
rect 77527 65501 77539 65504
rect 77481 65495 77539 65501
rect 78122 65492 78128 65504
rect 78180 65492 78186 65544
rect 1581 65399 1639 65405
rect 1581 65365 1593 65399
rect 1627 65396 1639 65399
rect 64506 65396 64512 65408
rect 1627 65368 64512 65396
rect 1627 65365 1639 65368
rect 1581 65359 1639 65365
rect 64506 65356 64512 65368
rect 64564 65356 64570 65408
rect 76006 65356 76012 65408
rect 76064 65396 76070 65408
rect 77941 65399 77999 65405
rect 77941 65396 77953 65399
rect 76064 65368 77953 65396
rect 76064 65356 76070 65368
rect 77941 65365 77953 65368
rect 77987 65365 77999 65399
rect 77941 65359 77999 65365
rect 1104 65306 78844 65328
rect 1104 65254 19574 65306
rect 19626 65254 19638 65306
rect 19690 65254 19702 65306
rect 19754 65254 19766 65306
rect 19818 65254 19830 65306
rect 19882 65254 50294 65306
rect 50346 65254 50358 65306
rect 50410 65254 50422 65306
rect 50474 65254 50486 65306
rect 50538 65254 50550 65306
rect 50602 65254 78844 65306
rect 1104 65232 78844 65254
rect 1581 65195 1639 65201
rect 1581 65161 1593 65195
rect 1627 65192 1639 65195
rect 2314 65192 2320 65204
rect 1627 65164 2320 65192
rect 1627 65161 1639 65164
rect 1581 65155 1639 65161
rect 2314 65152 2320 65164
rect 2372 65152 2378 65204
rect 1394 65056 1400 65068
rect 1307 65028 1400 65056
rect 1394 65016 1400 65028
rect 1452 65056 1458 65068
rect 2133 65059 2191 65065
rect 2133 65056 2145 65059
rect 1452 65028 2145 65056
rect 1452 65016 1458 65028
rect 2133 65025 2145 65028
rect 2179 65025 2191 65059
rect 2133 65019 2191 65025
rect 77297 65059 77355 65065
rect 77297 65025 77309 65059
rect 77343 65056 77355 65059
rect 77938 65056 77944 65068
rect 77343 65028 77944 65056
rect 77343 65025 77355 65028
rect 77297 65019 77355 65025
rect 77938 65016 77944 65028
rect 77996 65016 78002 65068
rect 72418 64948 72424 65000
rect 72476 64988 72482 65000
rect 72476 64960 77800 64988
rect 72476 64948 72482 64960
rect 77772 64929 77800 64960
rect 77757 64923 77815 64929
rect 77757 64889 77769 64923
rect 77803 64889 77815 64923
rect 77757 64883 77815 64889
rect 1104 64762 78844 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 34934 64762
rect 34986 64710 34998 64762
rect 35050 64710 35062 64762
rect 35114 64710 35126 64762
rect 35178 64710 35190 64762
rect 35242 64710 65654 64762
rect 65706 64710 65718 64762
rect 65770 64710 65782 64762
rect 65834 64710 65846 64762
rect 65898 64710 65910 64762
rect 65962 64710 78844 64762
rect 1104 64688 78844 64710
rect 1394 64444 1400 64456
rect 1355 64416 1400 64444
rect 1394 64404 1400 64416
rect 1452 64444 1458 64456
rect 2133 64447 2191 64453
rect 2133 64444 2145 64447
rect 1452 64416 2145 64444
rect 1452 64404 1458 64416
rect 2133 64413 2145 64416
rect 2179 64413 2191 64447
rect 2133 64407 2191 64413
rect 77481 64447 77539 64453
rect 77481 64413 77493 64447
rect 77527 64444 77539 64447
rect 78122 64444 78128 64456
rect 77527 64416 78128 64444
rect 77527 64413 77539 64416
rect 77481 64407 77539 64413
rect 78122 64404 78128 64416
rect 78180 64404 78186 64456
rect 1486 64268 1492 64320
rect 1544 64308 1550 64320
rect 1581 64311 1639 64317
rect 1581 64308 1593 64311
rect 1544 64280 1593 64308
rect 1544 64268 1550 64280
rect 1581 64277 1593 64280
rect 1627 64277 1639 64311
rect 1581 64271 1639 64277
rect 77478 64268 77484 64320
rect 77536 64308 77542 64320
rect 77941 64311 77999 64317
rect 77941 64308 77953 64311
rect 77536 64280 77953 64308
rect 77536 64268 77542 64280
rect 77941 64277 77953 64280
rect 77987 64277 77999 64311
rect 77941 64271 77999 64277
rect 1104 64218 78844 64240
rect 1104 64166 19574 64218
rect 19626 64166 19638 64218
rect 19690 64166 19702 64218
rect 19754 64166 19766 64218
rect 19818 64166 19830 64218
rect 19882 64166 50294 64218
rect 50346 64166 50358 64218
rect 50410 64166 50422 64218
rect 50474 64166 50486 64218
rect 50538 64166 50550 64218
rect 50602 64166 78844 64218
rect 1104 64144 78844 64166
rect 1394 63968 1400 63980
rect 1355 63940 1400 63968
rect 1394 63928 1400 63940
rect 1452 63968 1458 63980
rect 2133 63971 2191 63977
rect 2133 63968 2145 63971
rect 1452 63940 2145 63968
rect 1452 63928 1458 63940
rect 2133 63937 2145 63940
rect 2179 63937 2191 63971
rect 2133 63931 2191 63937
rect 77297 63971 77355 63977
rect 77297 63937 77309 63971
rect 77343 63968 77355 63971
rect 77938 63968 77944 63980
rect 77343 63940 77944 63968
rect 77343 63937 77355 63940
rect 77297 63931 77355 63937
rect 77938 63928 77944 63940
rect 77996 63928 78002 63980
rect 77757 63835 77815 63841
rect 77757 63832 77769 63835
rect 64846 63804 77769 63832
rect 1581 63767 1639 63773
rect 1581 63733 1593 63767
rect 1627 63764 1639 63767
rect 2222 63764 2228 63776
rect 1627 63736 2228 63764
rect 1627 63733 1639 63736
rect 1581 63727 1639 63733
rect 2222 63724 2228 63736
rect 2280 63724 2286 63776
rect 62666 63724 62672 63776
rect 62724 63764 62730 63776
rect 64846 63764 64874 63804
rect 77757 63801 77769 63804
rect 77803 63801 77815 63835
rect 77757 63795 77815 63801
rect 62724 63736 64874 63764
rect 62724 63724 62730 63736
rect 1104 63674 78844 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 34934 63674
rect 34986 63622 34998 63674
rect 35050 63622 35062 63674
rect 35114 63622 35126 63674
rect 35178 63622 35190 63674
rect 35242 63622 65654 63674
rect 65706 63622 65718 63674
rect 65770 63622 65782 63674
rect 65834 63622 65846 63674
rect 65898 63622 65910 63674
rect 65962 63622 78844 63674
rect 1104 63600 78844 63622
rect 1394 63220 1400 63232
rect 1355 63192 1400 63220
rect 1394 63180 1400 63192
rect 1452 63180 1458 63232
rect 77938 63180 77944 63232
rect 77996 63220 78002 63232
rect 78033 63223 78091 63229
rect 78033 63220 78045 63223
rect 77996 63192 78045 63220
rect 77996 63180 78002 63192
rect 78033 63189 78045 63192
rect 78079 63189 78091 63223
rect 78033 63183 78091 63189
rect 1104 63130 78844 63152
rect 1104 63078 19574 63130
rect 19626 63078 19638 63130
rect 19690 63078 19702 63130
rect 19754 63078 19766 63130
rect 19818 63078 19830 63130
rect 19882 63078 50294 63130
rect 50346 63078 50358 63130
rect 50410 63078 50422 63130
rect 50474 63078 50486 63130
rect 50538 63078 50550 63130
rect 50602 63078 78844 63130
rect 1104 63056 78844 63078
rect 1394 62880 1400 62892
rect 1355 62852 1400 62880
rect 1394 62840 1400 62852
rect 1452 62840 1458 62892
rect 77938 62880 77944 62892
rect 77899 62852 77944 62880
rect 77938 62840 77944 62852
rect 77996 62840 78002 62892
rect 1581 62679 1639 62685
rect 1581 62645 1593 62679
rect 1627 62676 1639 62679
rect 2130 62676 2136 62688
rect 1627 62648 2136 62676
rect 1627 62645 1639 62648
rect 1581 62639 1639 62645
rect 2130 62636 2136 62648
rect 2188 62636 2194 62688
rect 77294 62636 77300 62688
rect 77352 62676 77358 62688
rect 77757 62679 77815 62685
rect 77757 62676 77769 62679
rect 77352 62648 77769 62676
rect 77352 62636 77358 62648
rect 77757 62645 77769 62648
rect 77803 62645 77815 62679
rect 77757 62639 77815 62645
rect 1104 62586 78844 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 34934 62586
rect 34986 62534 34998 62586
rect 35050 62534 35062 62586
rect 35114 62534 35126 62586
rect 35178 62534 35190 62586
rect 35242 62534 65654 62586
rect 65706 62534 65718 62586
rect 65770 62534 65782 62586
rect 65834 62534 65846 62586
rect 65898 62534 65910 62586
rect 65962 62534 78844 62586
rect 1104 62512 78844 62534
rect 65426 62432 65432 62484
rect 65484 62472 65490 62484
rect 65705 62475 65763 62481
rect 65705 62472 65717 62475
rect 65484 62444 65717 62472
rect 65484 62432 65490 62444
rect 65705 62441 65717 62444
rect 65751 62472 65763 62475
rect 65978 62472 65984 62484
rect 65751 62444 65984 62472
rect 65751 62441 65763 62444
rect 65705 62435 65763 62441
rect 65978 62432 65984 62444
rect 66036 62432 66042 62484
rect 1394 62268 1400 62280
rect 1355 62240 1400 62268
rect 1394 62228 1400 62240
rect 1452 62268 1458 62280
rect 2133 62271 2191 62277
rect 2133 62268 2145 62271
rect 1452 62240 2145 62268
rect 1452 62228 1458 62240
rect 2133 62237 2145 62240
rect 2179 62237 2191 62271
rect 2133 62231 2191 62237
rect 77481 62271 77539 62277
rect 77481 62237 77493 62271
rect 77527 62268 77539 62271
rect 78122 62268 78128 62280
rect 77527 62240 78128 62268
rect 77527 62237 77539 62240
rect 77481 62231 77539 62237
rect 78122 62228 78128 62240
rect 78180 62228 78186 62280
rect 1762 62160 1768 62212
rect 1820 62200 1826 62212
rect 1820 62172 6914 62200
rect 1820 62160 1826 62172
rect 1581 62135 1639 62141
rect 1581 62101 1593 62135
rect 1627 62132 1639 62135
rect 1946 62132 1952 62144
rect 1627 62104 1952 62132
rect 1627 62101 1639 62104
rect 1581 62095 1639 62101
rect 1946 62092 1952 62104
rect 2004 62092 2010 62144
rect 6886 62132 6914 62172
rect 64233 62135 64291 62141
rect 64233 62132 64245 62135
rect 6886 62104 64245 62132
rect 64233 62101 64245 62104
rect 64279 62132 64291 62135
rect 64414 62132 64420 62144
rect 64279 62104 64420 62132
rect 64279 62101 64291 62104
rect 64233 62095 64291 62101
rect 64414 62092 64420 62104
rect 64472 62092 64478 62144
rect 77386 62092 77392 62144
rect 77444 62132 77450 62144
rect 77941 62135 77999 62141
rect 77941 62132 77953 62135
rect 77444 62104 77953 62132
rect 77444 62092 77450 62104
rect 77941 62101 77953 62104
rect 77987 62101 77999 62135
rect 77941 62095 77999 62101
rect 1104 62042 78844 62064
rect 1104 61990 19574 62042
rect 19626 61990 19638 62042
rect 19690 61990 19702 62042
rect 19754 61990 19766 62042
rect 19818 61990 19830 62042
rect 19882 61990 50294 62042
rect 50346 61990 50358 62042
rect 50410 61990 50422 62042
rect 50474 61990 50486 62042
rect 50538 61990 50550 62042
rect 50602 61990 78844 62042
rect 1104 61968 78844 61990
rect 64506 61928 64512 61940
rect 64467 61900 64512 61928
rect 64506 61888 64512 61900
rect 64564 61888 64570 61940
rect 65518 61888 65524 61940
rect 65576 61928 65582 61940
rect 66162 61928 66168 61940
rect 65576 61900 66168 61928
rect 65576 61888 65582 61900
rect 66162 61888 66168 61900
rect 66220 61888 66226 61940
rect 65334 61820 65340 61872
rect 65392 61860 65398 61872
rect 65705 61863 65763 61869
rect 65705 61860 65717 61863
rect 65392 61832 65717 61860
rect 65392 61820 65398 61832
rect 65705 61829 65717 61832
rect 65751 61860 65763 61863
rect 66070 61860 66076 61872
rect 65751 61832 66076 61860
rect 65751 61829 65763 61832
rect 65705 61823 65763 61829
rect 66070 61820 66076 61832
rect 66128 61820 66134 61872
rect 1394 61792 1400 61804
rect 1355 61764 1400 61792
rect 1394 61752 1400 61764
rect 1452 61792 1458 61804
rect 2133 61795 2191 61801
rect 2133 61792 2145 61795
rect 1452 61764 2145 61792
rect 1452 61752 1458 61764
rect 2133 61761 2145 61764
rect 2179 61761 2191 61795
rect 64046 61792 64052 61804
rect 64007 61764 64052 61792
rect 2133 61755 2191 61761
rect 64046 61752 64052 61764
rect 64104 61752 64110 61804
rect 77297 61795 77355 61801
rect 77297 61761 77309 61795
rect 77343 61792 77355 61795
rect 77938 61792 77944 61804
rect 77343 61764 77944 61792
rect 77343 61761 77355 61764
rect 77297 61755 77355 61761
rect 77938 61752 77944 61764
rect 77996 61752 78002 61804
rect 61654 61616 61660 61668
rect 61712 61656 61718 61668
rect 64322 61656 64328 61668
rect 61712 61628 64328 61656
rect 61712 61616 61718 61628
rect 64322 61616 64328 61628
rect 64380 61656 64386 61668
rect 65061 61659 65119 61665
rect 65061 61656 65073 61659
rect 64380 61628 65073 61656
rect 64380 61616 64386 61628
rect 65061 61625 65073 61628
rect 65107 61625 65119 61659
rect 65061 61619 65119 61625
rect 1581 61591 1639 61597
rect 1581 61557 1593 61591
rect 1627 61588 1639 61591
rect 2406 61588 2412 61600
rect 1627 61560 2412 61588
rect 1627 61557 1639 61560
rect 1581 61551 1639 61557
rect 2406 61548 2412 61560
rect 2464 61548 2470 61600
rect 2682 61548 2688 61600
rect 2740 61588 2746 61600
rect 63865 61591 63923 61597
rect 63865 61588 63877 61591
rect 2740 61560 63877 61588
rect 2740 61548 2746 61560
rect 63865 61557 63877 61560
rect 63911 61557 63923 61591
rect 63865 61551 63923 61557
rect 66070 61548 66076 61600
rect 66128 61588 66134 61600
rect 66717 61591 66775 61597
rect 66717 61588 66729 61591
rect 66128 61560 66729 61588
rect 66128 61548 66134 61560
rect 66717 61557 66729 61560
rect 66763 61557 66775 61591
rect 77754 61588 77760 61600
rect 77715 61560 77760 61588
rect 66717 61551 66775 61557
rect 77754 61548 77760 61560
rect 77812 61548 77818 61600
rect 1104 61498 78844 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 65654 61498
rect 65706 61446 65718 61498
rect 65770 61446 65782 61498
rect 65834 61446 65846 61498
rect 65898 61446 65910 61498
rect 65962 61446 78844 61498
rect 1104 61424 78844 61446
rect 1578 61344 1584 61396
rect 1636 61384 1642 61396
rect 61654 61384 61660 61396
rect 1636 61356 61660 61384
rect 1636 61344 1642 61356
rect 61654 61344 61660 61356
rect 61712 61344 61718 61396
rect 63126 61384 63132 61396
rect 63087 61356 63132 61384
rect 63126 61344 63132 61356
rect 63184 61344 63190 61396
rect 63218 61344 63224 61396
rect 63276 61384 63282 61396
rect 63276 61356 74534 61384
rect 63276 61344 63282 61356
rect 64966 61316 64972 61328
rect 64927 61288 64972 61316
rect 64966 61276 64972 61288
rect 65024 61276 65030 61328
rect 66162 61316 66168 61328
rect 66123 61288 66168 61316
rect 66162 61276 66168 61288
rect 66220 61276 66226 61328
rect 74506 61248 74534 61356
rect 77754 61248 77760 61260
rect 74506 61220 77760 61248
rect 77754 61208 77760 61220
rect 77812 61208 77818 61260
rect 1394 61180 1400 61192
rect 1355 61152 1400 61180
rect 1394 61140 1400 61152
rect 1452 61180 1458 61192
rect 2133 61183 2191 61189
rect 2133 61180 2145 61183
rect 1452 61152 2145 61180
rect 1452 61140 1458 61152
rect 2133 61149 2145 61152
rect 2179 61149 2191 61183
rect 63954 61180 63960 61192
rect 63915 61152 63960 61180
rect 2133 61143 2191 61149
rect 63954 61140 63960 61152
rect 64012 61140 64018 61192
rect 64414 61180 64420 61192
rect 64375 61152 64420 61180
rect 64414 61140 64420 61152
rect 64472 61140 64478 61192
rect 64837 61183 64895 61189
rect 64837 61149 64849 61183
rect 64883 61180 64895 61183
rect 65242 61180 65248 61192
rect 64883 61152 65248 61180
rect 64883 61149 64895 61152
rect 64837 61143 64895 61149
rect 65242 61140 65248 61152
rect 65300 61140 65306 61192
rect 65518 61140 65524 61192
rect 65576 61180 65582 61192
rect 65613 61183 65671 61189
rect 65613 61180 65625 61183
rect 65576 61152 65625 61180
rect 65576 61140 65582 61152
rect 65613 61149 65625 61152
rect 65659 61149 65671 61183
rect 65613 61143 65671 61149
rect 65978 61140 65984 61192
rect 66036 61189 66042 61192
rect 66036 61180 66044 61189
rect 66714 61180 66720 61192
rect 66036 61152 66081 61180
rect 66675 61152 66720 61180
rect 66036 61143 66044 61152
rect 66036 61140 66042 61143
rect 66714 61140 66720 61152
rect 66772 61140 66778 61192
rect 67453 61183 67511 61189
rect 67453 61180 67465 61183
rect 66824 61152 67465 61180
rect 63678 61072 63684 61124
rect 63736 61112 63742 61124
rect 64601 61115 64659 61121
rect 64601 61112 64613 61115
rect 63736 61084 64613 61112
rect 63736 61072 63742 61084
rect 64601 61081 64613 61084
rect 64647 61081 64659 61115
rect 64601 61075 64659 61081
rect 64693 61115 64751 61121
rect 64693 61081 64705 61115
rect 64739 61112 64751 61115
rect 65426 61112 65432 61124
rect 64739 61084 65432 61112
rect 64739 61081 64751 61084
rect 64693 61075 64751 61081
rect 1581 61047 1639 61053
rect 1581 61013 1593 61047
rect 1627 61044 1639 61047
rect 2038 61044 2044 61056
rect 1627 61016 2044 61044
rect 1627 61013 1639 61016
rect 1581 61007 1639 61013
rect 2038 61004 2044 61016
rect 2096 61004 2102 61056
rect 63770 61044 63776 61056
rect 63731 61016 63776 61044
rect 63770 61004 63776 61016
rect 63828 61004 63834 61056
rect 64616 61044 64644 61075
rect 65426 61072 65432 61084
rect 65484 61072 65490 61124
rect 65797 61115 65855 61121
rect 65797 61081 65809 61115
rect 65843 61081 65855 61115
rect 65797 61075 65855 61081
rect 65889 61115 65947 61121
rect 65889 61081 65901 61115
rect 65935 61112 65947 61115
rect 66824 61112 66852 61152
rect 67453 61149 67465 61152
rect 67499 61180 67511 61183
rect 75178 61180 75184 61192
rect 67499 61152 75184 61180
rect 67499 61149 67511 61152
rect 67453 61143 67511 61149
rect 75178 61140 75184 61152
rect 75236 61140 75242 61192
rect 77481 61183 77539 61189
rect 77481 61149 77493 61183
rect 77527 61180 77539 61183
rect 78122 61180 78128 61192
rect 77527 61152 78128 61180
rect 77527 61149 77539 61152
rect 77481 61143 77539 61149
rect 78122 61140 78128 61152
rect 78180 61140 78186 61192
rect 77018 61112 77024 61124
rect 65935 61084 66852 61112
rect 66916 61084 77024 61112
rect 65935 61081 65947 61084
rect 65889 61075 65947 61081
rect 65812 61044 65840 61075
rect 66916 61053 66944 61084
rect 77018 61072 77024 61084
rect 77076 61072 77082 61124
rect 64616 61016 65840 61044
rect 66901 61047 66959 61053
rect 66901 61013 66913 61047
rect 66947 61013 66959 61047
rect 77938 61044 77944 61056
rect 77899 61016 77944 61044
rect 66901 61007 66959 61013
rect 77938 61004 77944 61016
rect 77996 61004 78002 61056
rect 1104 60954 78844 60976
rect 1104 60902 19574 60954
rect 19626 60902 19638 60954
rect 19690 60902 19702 60954
rect 19754 60902 19766 60954
rect 19818 60902 19830 60954
rect 19882 60902 50294 60954
rect 50346 60902 50358 60954
rect 50410 60902 50422 60954
rect 50474 60902 50486 60954
rect 50538 60902 50550 60954
rect 50602 60902 78844 60954
rect 1104 60880 78844 60902
rect 63957 60843 64015 60849
rect 63957 60809 63969 60843
rect 64003 60840 64015 60843
rect 64046 60840 64052 60852
rect 64003 60812 64052 60840
rect 64003 60809 64015 60812
rect 63957 60803 64015 60809
rect 64046 60800 64052 60812
rect 64104 60800 64110 60852
rect 64156 60812 64874 60840
rect 59998 60732 60004 60784
rect 60056 60772 60062 60784
rect 64156 60772 64184 60812
rect 60056 60744 64184 60772
rect 64846 60772 64874 60812
rect 77938 60772 77944 60784
rect 64846 60744 77944 60772
rect 60056 60732 60062 60744
rect 77938 60732 77944 60744
rect 77996 60732 78002 60784
rect 63678 60664 63684 60716
rect 63736 60704 63742 60716
rect 63773 60707 63831 60713
rect 63773 60704 63785 60707
rect 63736 60676 63785 60704
rect 63736 60664 63742 60676
rect 63773 60673 63785 60676
rect 63819 60673 63831 60707
rect 63773 60667 63831 60673
rect 64322 60664 64328 60716
rect 64380 60704 64386 60716
rect 64417 60707 64475 60713
rect 64417 60704 64429 60707
rect 64380 60676 64429 60704
rect 64380 60664 64386 60676
rect 64417 60673 64429 60676
rect 64463 60673 64475 60707
rect 64598 60704 64604 60716
rect 64559 60676 64604 60704
rect 64417 60667 64475 60673
rect 64598 60664 64604 60676
rect 64656 60664 64662 60716
rect 64693 60707 64751 60713
rect 64693 60673 64705 60707
rect 64739 60673 64751 60707
rect 64693 60667 64751 60673
rect 63589 60639 63647 60645
rect 63589 60605 63601 60639
rect 63635 60605 63647 60639
rect 64708 60636 64736 60667
rect 64782 60664 64788 60716
rect 64840 60713 64846 60716
rect 64840 60704 64848 60713
rect 64840 60676 64885 60704
rect 64840 60667 64848 60676
rect 64840 60664 64846 60667
rect 65242 60664 65248 60716
rect 65300 60704 65306 60716
rect 65426 60704 65432 60716
rect 65300 60676 65432 60704
rect 65300 60664 65306 60676
rect 65426 60664 65432 60676
rect 65484 60704 65490 60716
rect 65705 60707 65763 60713
rect 65705 60704 65717 60707
rect 65484 60676 65717 60704
rect 65484 60664 65490 60676
rect 65705 60673 65717 60676
rect 65751 60704 65763 60707
rect 65978 60704 65984 60716
rect 65751 60676 65984 60704
rect 65751 60673 65763 60676
rect 65705 60667 65763 60673
rect 65978 60664 65984 60676
rect 66036 60664 66042 60716
rect 65334 60636 65340 60648
rect 64708 60608 65340 60636
rect 63589 60599 63647 60605
rect 62485 60571 62543 60577
rect 62485 60537 62497 60571
rect 62531 60568 62543 60571
rect 63604 60568 63632 60599
rect 65334 60596 65340 60608
rect 65392 60596 65398 60648
rect 65518 60636 65524 60648
rect 65479 60608 65524 60636
rect 65518 60596 65524 60608
rect 65576 60596 65582 60648
rect 65889 60639 65947 60645
rect 65889 60605 65901 60639
rect 65935 60636 65947 60639
rect 66349 60639 66407 60645
rect 66349 60636 66361 60639
rect 65935 60608 66361 60636
rect 65935 60605 65947 60608
rect 65889 60599 65947 60605
rect 66349 60605 66361 60608
rect 66395 60605 66407 60639
rect 66349 60599 66407 60605
rect 66625 60639 66683 60645
rect 66625 60605 66637 60639
rect 66671 60636 66683 60639
rect 76558 60636 76564 60648
rect 66671 60608 76564 60636
rect 66671 60605 66683 60608
rect 66625 60599 66683 60605
rect 76558 60596 76564 60608
rect 76616 60596 76622 60648
rect 67358 60568 67364 60580
rect 62531 60540 67364 60568
rect 62531 60537 62543 60540
rect 62485 60531 62543 60537
rect 67358 60528 67364 60540
rect 67416 60528 67422 60580
rect 1394 60500 1400 60512
rect 1355 60472 1400 60500
rect 1394 60460 1400 60472
rect 1452 60460 1458 60512
rect 63034 60500 63040 60512
rect 62995 60472 63040 60500
rect 63034 60460 63040 60472
rect 63092 60460 63098 60512
rect 64969 60503 65027 60509
rect 64969 60469 64981 60503
rect 65015 60500 65027 60503
rect 65150 60500 65156 60512
rect 65015 60472 65156 60500
rect 65015 60469 65027 60472
rect 64969 60463 65027 60469
rect 65150 60460 65156 60472
rect 65208 60460 65214 60512
rect 65518 60460 65524 60512
rect 65576 60500 65582 60512
rect 66070 60500 66076 60512
rect 65576 60472 66076 60500
rect 65576 60460 65582 60472
rect 66070 60460 66076 60472
rect 66128 60460 66134 60512
rect 1104 60410 78844 60432
rect 1104 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 65654 60410
rect 65706 60358 65718 60410
rect 65770 60358 65782 60410
rect 65834 60358 65846 60410
rect 65898 60358 65910 60410
rect 65962 60358 78844 60410
rect 1104 60336 78844 60358
rect 62666 60296 62672 60308
rect 62627 60268 62672 60296
rect 62666 60256 62672 60268
rect 62724 60256 62730 60308
rect 63954 60296 63960 60308
rect 63915 60268 63960 60296
rect 63954 60256 63960 60268
rect 64012 60256 64018 60308
rect 65242 60296 65248 60308
rect 64892 60268 65248 60296
rect 59538 60188 59544 60240
rect 59596 60228 59602 60240
rect 64892 60228 64920 60268
rect 65242 60256 65248 60268
rect 65300 60256 65306 60308
rect 66714 60296 66720 60308
rect 66675 60268 66720 60296
rect 66714 60256 66720 60268
rect 66772 60256 66778 60308
rect 76650 60296 76656 60308
rect 70366 60268 76656 60296
rect 59596 60200 64920 60228
rect 64969 60231 65027 60237
rect 59596 60188 59602 60200
rect 64969 60197 64981 60231
rect 65015 60228 65027 60231
rect 65058 60228 65064 60240
rect 65015 60200 65064 60228
rect 65015 60197 65027 60200
rect 64969 60191 65027 60197
rect 65058 60188 65064 60200
rect 65116 60188 65122 60240
rect 65352 60200 65840 60228
rect 65352 60160 65380 60200
rect 63788 60132 65380 60160
rect 1394 60092 1400 60104
rect 1355 60064 1400 60092
rect 1394 60052 1400 60064
rect 1452 60052 1458 60104
rect 62117 60095 62175 60101
rect 62117 60061 62129 60095
rect 62163 60092 62175 60095
rect 63586 60092 63592 60104
rect 62163 60064 63592 60092
rect 62163 60061 62175 60064
rect 62117 60055 62175 60061
rect 63586 60052 63592 60064
rect 63644 60052 63650 60104
rect 63678 60052 63684 60104
rect 63736 60092 63742 60104
rect 63788 60101 63816 60132
rect 63773 60095 63831 60101
rect 63773 60092 63785 60095
rect 63736 60064 63785 60092
rect 63736 60052 63742 60064
rect 63773 60061 63785 60064
rect 63819 60061 63831 60095
rect 63773 60055 63831 60061
rect 64417 60095 64475 60101
rect 64417 60061 64429 60095
rect 64463 60092 64475 60095
rect 64506 60092 64512 60104
rect 64463 60064 64512 60092
rect 64463 60061 64475 60064
rect 64417 60055 64475 60061
rect 64506 60052 64512 60064
rect 64564 60052 64570 60104
rect 64782 60052 64788 60104
rect 64840 60101 64846 60104
rect 64840 60092 64848 60101
rect 65610 60092 65616 60104
rect 64840 60064 64885 60092
rect 65571 60064 65616 60092
rect 64840 60055 64848 60064
rect 64840 60052 64846 60055
rect 65610 60052 65616 60064
rect 65668 60052 65674 60104
rect 65812 60101 65840 60200
rect 66070 60188 66076 60240
rect 66128 60228 66134 60240
rect 66165 60231 66223 60237
rect 66165 60228 66177 60231
rect 66128 60200 66177 60228
rect 66128 60188 66134 60200
rect 66165 60197 66177 60200
rect 66211 60197 66223 60231
rect 68094 60228 68100 60240
rect 68055 60200 68100 60228
rect 66165 60191 66223 60197
rect 68094 60188 68100 60200
rect 68152 60188 68158 60240
rect 68649 60163 68707 60169
rect 68649 60160 68661 60163
rect 65904 60132 68661 60160
rect 65904 60101 65932 60132
rect 68649 60129 68661 60132
rect 68695 60160 68707 60163
rect 70366 60160 70394 60268
rect 76650 60256 76656 60268
rect 76708 60256 76714 60308
rect 68695 60132 70394 60160
rect 68695 60129 68707 60132
rect 68649 60123 68707 60129
rect 65797 60095 65855 60101
rect 65797 60061 65809 60095
rect 65843 60061 65855 60095
rect 65797 60055 65855 60061
rect 65889 60095 65947 60101
rect 65889 60061 65901 60095
rect 65935 60061 65947 60095
rect 65889 60055 65947 60061
rect 65978 60052 65984 60104
rect 66036 60101 66042 60104
rect 66036 60092 66044 60101
rect 66901 60095 66959 60101
rect 66901 60092 66913 60095
rect 66036 60064 66913 60092
rect 66036 60055 66044 60064
rect 66901 60061 66913 60064
rect 66947 60061 66959 60095
rect 66901 60055 66959 60061
rect 67085 60095 67143 60101
rect 67085 60061 67097 60095
rect 67131 60092 67143 60095
rect 67358 60092 67364 60104
rect 67131 60064 67364 60092
rect 67131 60061 67143 60064
rect 67085 60055 67143 60061
rect 66036 60052 66042 60055
rect 67358 60052 67364 60064
rect 67416 60052 67422 60104
rect 77481 60095 77539 60101
rect 77481 60061 77493 60095
rect 77527 60092 77539 60095
rect 78122 60092 78128 60104
rect 77527 60064 78128 60092
rect 77527 60061 77539 60064
rect 77481 60055 77539 60061
rect 78122 60052 78128 60064
rect 78180 60052 78186 60104
rect 64598 60024 64604 60036
rect 64559 59996 64604 60024
rect 64598 59984 64604 59996
rect 64656 59984 64662 60036
rect 64693 60027 64751 60033
rect 64693 59993 64705 60027
rect 64739 59993 64751 60027
rect 64693 59987 64751 59993
rect 1581 59959 1639 59965
rect 1581 59925 1593 59959
rect 1627 59956 1639 59959
rect 2590 59956 2596 59968
rect 1627 59928 2596 59956
rect 1627 59925 1639 59928
rect 1581 59919 1639 59925
rect 2590 59916 2596 59928
rect 2648 59916 2654 59968
rect 64708 59956 64736 59987
rect 65702 59984 65708 60036
rect 65760 60024 65766 60036
rect 66990 60024 66996 60036
rect 65760 59996 66996 60024
rect 65760 59984 65766 59996
rect 66990 59984 66996 59996
rect 67048 59984 67054 60036
rect 67637 60027 67695 60033
rect 67637 59993 67649 60027
rect 67683 60024 67695 60027
rect 76006 60024 76012 60036
rect 67683 59996 76012 60024
rect 67683 59993 67695 59996
rect 67637 59987 67695 59993
rect 67652 59956 67680 59987
rect 76006 59984 76012 59996
rect 76064 59984 76070 60036
rect 77938 59956 77944 59968
rect 64708 59928 67680 59956
rect 77899 59928 77944 59956
rect 77938 59916 77944 59928
rect 77996 59916 78002 59968
rect 1104 59866 78844 59888
rect 1104 59814 19574 59866
rect 19626 59814 19638 59866
rect 19690 59814 19702 59866
rect 19754 59814 19766 59866
rect 19818 59814 19830 59866
rect 19882 59814 50294 59866
rect 50346 59814 50358 59866
rect 50410 59814 50422 59866
rect 50474 59814 50486 59866
rect 50538 59814 50550 59866
rect 50602 59814 78844 59866
rect 1104 59792 78844 59814
rect 62114 59712 62120 59764
rect 62172 59752 62178 59764
rect 62485 59755 62543 59761
rect 62485 59752 62497 59755
rect 62172 59724 62497 59752
rect 62172 59712 62178 59724
rect 62485 59721 62497 59724
rect 62531 59752 62543 59755
rect 63218 59752 63224 59764
rect 62531 59724 63224 59752
rect 62531 59721 62543 59724
rect 62485 59715 62543 59721
rect 63218 59712 63224 59724
rect 63276 59712 63282 59764
rect 64874 59712 64880 59764
rect 64932 59752 64938 59764
rect 64932 59724 65196 59752
rect 64932 59712 64938 59724
rect 63497 59687 63555 59693
rect 63497 59653 63509 59687
rect 63543 59684 63555 59687
rect 64690 59684 64696 59696
rect 63543 59656 64552 59684
rect 64651 59656 64696 59684
rect 63543 59653 63555 59656
rect 63497 59647 63555 59653
rect 1394 59616 1400 59628
rect 1355 59588 1400 59616
rect 1394 59576 1400 59588
rect 1452 59616 1458 59628
rect 2133 59619 2191 59625
rect 2133 59616 2145 59619
rect 1452 59588 2145 59616
rect 1452 59576 1458 59588
rect 2133 59585 2145 59588
rect 2179 59585 2191 59619
rect 2133 59579 2191 59585
rect 63126 59576 63132 59628
rect 63184 59616 63190 59628
rect 63770 59625 63776 59628
rect 63313 59619 63371 59625
rect 63313 59616 63325 59619
rect 63184 59588 63325 59616
rect 63184 59576 63190 59588
rect 63313 59585 63325 59588
rect 63359 59585 63371 59619
rect 63313 59579 63371 59585
rect 63589 59619 63647 59625
rect 63589 59585 63601 59619
rect 63635 59585 63647 59619
rect 63589 59579 63647 59585
rect 63733 59619 63776 59625
rect 63733 59585 63745 59619
rect 63733 59579 63776 59585
rect 2314 59508 2320 59560
rect 2372 59548 2378 59560
rect 63604 59548 63632 59579
rect 63770 59576 63776 59579
rect 63828 59576 63834 59628
rect 64414 59616 64420 59628
rect 64375 59588 64420 59616
rect 64414 59576 64420 59588
rect 64472 59576 64478 59628
rect 64524 59616 64552 59656
rect 64690 59644 64696 59656
rect 64748 59644 64754 59696
rect 64892 59684 64920 59712
rect 64852 59656 64920 59684
rect 65168 59684 65196 59724
rect 65242 59712 65248 59764
rect 65300 59752 65306 59764
rect 77938 59752 77944 59764
rect 65300 59724 77944 59752
rect 65300 59712 65306 59724
rect 77938 59712 77944 59724
rect 77996 59712 78002 59764
rect 65168 59656 65984 59684
rect 64598 59616 64604 59628
rect 64524 59588 64604 59616
rect 64598 59576 64604 59588
rect 64656 59576 64662 59628
rect 64852 59625 64880 59656
rect 64831 59619 64889 59625
rect 64831 59585 64843 59619
rect 64877 59585 64889 59619
rect 64831 59579 64889 59585
rect 65541 59619 65599 59625
rect 65541 59585 65553 59619
rect 65587 59616 65599 59619
rect 65705 59619 65763 59625
rect 65587 59588 65656 59616
rect 65587 59585 65599 59588
rect 65541 59579 65599 59585
rect 64986 59551 65044 59557
rect 2372 59520 16574 59548
rect 63604 59520 64736 59548
rect 2372 59508 2378 59520
rect 2222 59440 2228 59492
rect 2280 59480 2286 59492
rect 16546 59480 16574 59520
rect 64414 59480 64420 59492
rect 2280 59452 6914 59480
rect 16546 59452 64420 59480
rect 2280 59440 2286 59452
rect 1581 59415 1639 59421
rect 1581 59381 1593 59415
rect 1627 59412 1639 59415
rect 2682 59412 2688 59424
rect 1627 59384 2688 59412
rect 1627 59381 1639 59384
rect 1581 59375 1639 59381
rect 2682 59372 2688 59384
rect 2740 59372 2746 59424
rect 6886 59412 6914 59452
rect 64414 59440 64420 59452
rect 64472 59440 64478 59492
rect 61657 59415 61715 59421
rect 61657 59412 61669 59415
rect 6886 59384 61669 59412
rect 61657 59381 61669 59384
rect 61703 59412 61715 59415
rect 61838 59412 61844 59424
rect 61703 59384 61844 59412
rect 61703 59381 61715 59384
rect 61657 59375 61715 59381
rect 61838 59372 61844 59384
rect 61896 59372 61902 59424
rect 63862 59412 63868 59424
rect 63823 59384 63868 59412
rect 63862 59372 63868 59384
rect 63920 59372 63926 59424
rect 64708 59412 64736 59520
rect 64986 59517 64998 59551
rect 65032 59548 65044 59551
rect 65242 59548 65248 59560
rect 65032 59520 65248 59548
rect 65032 59517 65044 59520
rect 64986 59511 65044 59517
rect 65242 59508 65248 59520
rect 65300 59508 65306 59560
rect 64892 59452 65288 59480
rect 64892 59412 64920 59452
rect 64708 59384 64920 59412
rect 65260 59412 65288 59452
rect 65334 59440 65340 59492
rect 65392 59480 65398 59492
rect 65628 59480 65656 59588
rect 65705 59585 65717 59619
rect 65751 59585 65763 59619
rect 65705 59579 65763 59585
rect 65720 59492 65748 59579
rect 65794 59576 65800 59628
rect 65852 59616 65858 59628
rect 65956 59625 65984 59656
rect 67174 59644 67180 59696
rect 67232 59684 67238 59696
rect 72418 59684 72424 59696
rect 67232 59656 72424 59684
rect 67232 59644 67238 59656
rect 72418 59644 72424 59656
rect 72476 59644 72482 59696
rect 65941 59619 65999 59625
rect 65852 59588 65897 59616
rect 65852 59576 65858 59588
rect 65941 59585 65953 59619
rect 65987 59585 65999 59619
rect 65941 59579 65999 59585
rect 77297 59619 77355 59625
rect 77297 59585 77309 59619
rect 77343 59616 77355 59619
rect 77938 59616 77944 59628
rect 77343 59588 77944 59616
rect 77343 59585 77355 59588
rect 77297 59579 77355 59585
rect 77938 59576 77944 59588
rect 77996 59576 78002 59628
rect 72326 59548 72332 59560
rect 67606 59520 72332 59548
rect 65392 59452 65656 59480
rect 65392 59440 65398 59452
rect 65702 59440 65708 59492
rect 65760 59440 65766 59492
rect 66625 59483 66683 59489
rect 66625 59480 66637 59483
rect 65904 59452 66637 59480
rect 65904 59412 65932 59452
rect 66625 59449 66637 59452
rect 66671 59480 66683 59483
rect 67606 59480 67634 59520
rect 72326 59508 72332 59520
rect 72384 59508 72390 59560
rect 66671 59452 67634 59480
rect 66671 59449 66683 59452
rect 66625 59443 66683 59449
rect 65260 59384 65932 59412
rect 65978 59372 65984 59424
rect 66036 59412 66042 59424
rect 66073 59415 66131 59421
rect 66073 59412 66085 59415
rect 66036 59384 66085 59412
rect 66036 59372 66042 59384
rect 66073 59381 66085 59384
rect 66119 59381 66131 59415
rect 67174 59412 67180 59424
rect 67135 59384 67180 59412
rect 66073 59375 66131 59381
rect 67174 59372 67180 59384
rect 67232 59372 67238 59424
rect 77754 59412 77760 59424
rect 77715 59384 77760 59412
rect 77754 59372 77760 59384
rect 77812 59372 77818 59424
rect 1104 59322 78844 59344
rect 1104 59270 4214 59322
rect 4266 59270 4278 59322
rect 4330 59270 4342 59322
rect 4394 59270 4406 59322
rect 4458 59270 4470 59322
rect 4522 59270 34934 59322
rect 34986 59270 34998 59322
rect 35050 59270 35062 59322
rect 35114 59270 35126 59322
rect 35178 59270 35190 59322
rect 35242 59270 65654 59322
rect 65706 59270 65718 59322
rect 65770 59270 65782 59322
rect 65834 59270 65846 59322
rect 65898 59270 65910 59322
rect 65962 59270 78844 59322
rect 1104 59248 78844 59270
rect 63313 59211 63371 59217
rect 63313 59177 63325 59211
rect 63359 59208 63371 59211
rect 63678 59208 63684 59220
rect 63359 59180 63684 59208
rect 63359 59177 63371 59180
rect 63313 59171 63371 59177
rect 63678 59168 63684 59180
rect 63736 59168 63742 59220
rect 64371 59211 64429 59217
rect 64371 59177 64383 59211
rect 64417 59208 64429 59211
rect 64598 59208 64604 59220
rect 64417 59180 64604 59208
rect 64417 59177 64429 59180
rect 64371 59171 64429 59177
rect 64598 59168 64604 59180
rect 64656 59168 64662 59220
rect 65426 59168 65432 59220
rect 65484 59208 65490 59220
rect 65797 59211 65855 59217
rect 65797 59208 65809 59211
rect 65484 59180 65809 59208
rect 65484 59168 65490 59180
rect 65797 59177 65809 59180
rect 65843 59177 65855 59211
rect 65797 59171 65855 59177
rect 62393 59143 62451 59149
rect 62393 59109 62405 59143
rect 62439 59140 62451 59143
rect 62482 59140 62488 59152
rect 62439 59112 62488 59140
rect 62439 59109 62451 59112
rect 62393 59103 62451 59109
rect 62482 59100 62488 59112
rect 62540 59100 62546 59152
rect 64690 59100 64696 59152
rect 64748 59140 64754 59152
rect 67174 59140 67180 59152
rect 64748 59112 67180 59140
rect 64748 59100 64754 59112
rect 67174 59100 67180 59112
rect 67232 59100 67238 59152
rect 60274 59032 60280 59084
rect 60332 59072 60338 59084
rect 60737 59075 60795 59081
rect 60737 59072 60749 59075
rect 60332 59044 60749 59072
rect 60332 59032 60338 59044
rect 60737 59041 60749 59044
rect 60783 59072 60795 59075
rect 60783 59044 74534 59072
rect 60783 59041 60795 59044
rect 60737 59035 60795 59041
rect 1394 59004 1400 59016
rect 1355 58976 1400 59004
rect 1394 58964 1400 58976
rect 1452 59004 1458 59016
rect 2133 59007 2191 59013
rect 2133 59004 2145 59007
rect 1452 58976 2145 59004
rect 1452 58964 1458 58976
rect 2133 58973 2145 58976
rect 2179 58973 2191 59007
rect 2133 58967 2191 58973
rect 2406 58964 2412 59016
rect 2464 59004 2470 59016
rect 61654 59004 61660 59016
rect 2464 58976 61660 59004
rect 2464 58964 2470 58976
rect 61654 58964 61660 58976
rect 61712 58964 61718 59016
rect 61838 59004 61844 59016
rect 61799 58976 61844 59004
rect 61838 58964 61844 58976
rect 61896 58964 61902 59016
rect 62206 58964 62212 59016
rect 62264 59013 62270 59016
rect 62264 59004 62272 59013
rect 63126 59004 63132 59016
rect 62264 58976 62309 59004
rect 63087 58976 63132 59004
rect 62264 58967 62272 58976
rect 62264 58964 62270 58967
rect 63126 58964 63132 58976
rect 63184 58964 63190 59016
rect 64601 59007 64659 59013
rect 64601 58973 64613 59007
rect 64647 58973 64659 59007
rect 65610 59004 65616 59016
rect 65571 58976 65616 59004
rect 64601 58967 64659 58973
rect 61930 58896 61936 58948
rect 61988 58936 61994 58948
rect 62025 58939 62083 58945
rect 62025 58936 62037 58939
rect 61988 58908 62037 58936
rect 61988 58896 61994 58908
rect 62025 58905 62037 58908
rect 62071 58905 62083 58939
rect 62025 58899 62083 58905
rect 62117 58939 62175 58945
rect 62117 58905 62129 58939
rect 62163 58936 62175 58939
rect 62666 58936 62672 58948
rect 62163 58908 62672 58936
rect 62163 58905 62175 58908
rect 62117 58899 62175 58905
rect 62666 58896 62672 58908
rect 62724 58896 62730 58948
rect 63144 58936 63172 58964
rect 64616 58936 64644 58967
rect 65610 58964 65616 58976
rect 65668 59004 65674 59016
rect 66809 59007 66867 59013
rect 66809 59004 66821 59007
rect 65668 58976 66821 59004
rect 65668 58964 65674 58976
rect 66809 58973 66821 58976
rect 66855 58973 66867 59007
rect 66809 58967 66867 58973
rect 66257 58939 66315 58945
rect 66257 58936 66269 58939
rect 63144 58908 66269 58936
rect 66257 58905 66269 58908
rect 66303 58905 66315 58939
rect 74506 58936 74534 59044
rect 77481 59007 77539 59013
rect 77481 58973 77493 59007
rect 77527 59004 77539 59007
rect 78122 59004 78128 59016
rect 77527 58976 78128 59004
rect 77527 58973 77539 58976
rect 77481 58967 77539 58973
rect 78122 58964 78128 58976
rect 78180 58964 78186 59016
rect 77754 58936 77760 58948
rect 74506 58908 77760 58936
rect 66257 58899 66315 58905
rect 77754 58896 77760 58908
rect 77812 58896 77818 58948
rect 1578 58868 1584 58880
rect 1539 58840 1584 58868
rect 1578 58828 1584 58840
rect 1636 58828 1642 58880
rect 59814 58868 59820 58880
rect 59775 58840 59820 58868
rect 59814 58828 59820 58840
rect 59872 58828 59878 58880
rect 61286 58868 61292 58880
rect 61247 58840 61292 58868
rect 61286 58828 61292 58840
rect 61344 58828 61350 58880
rect 67358 58868 67364 58880
rect 67319 58840 67364 58868
rect 67358 58828 67364 58840
rect 67416 58828 67422 58880
rect 77938 58868 77944 58880
rect 77899 58840 77944 58868
rect 77938 58828 77944 58840
rect 77996 58828 78002 58880
rect 1104 58778 78844 58800
rect 1104 58726 19574 58778
rect 19626 58726 19638 58778
rect 19690 58726 19702 58778
rect 19754 58726 19766 58778
rect 19818 58726 19830 58778
rect 19882 58726 50294 58778
rect 50346 58726 50358 58778
rect 50410 58726 50422 58778
rect 50474 58726 50486 58778
rect 50538 58726 50550 58778
rect 50602 58726 78844 58778
rect 1104 58704 78844 58726
rect 2682 58624 2688 58676
rect 2740 58664 2746 58676
rect 59538 58664 59544 58676
rect 2740 58636 51074 58664
rect 59499 58636 59544 58664
rect 2740 58624 2746 58636
rect 1578 58556 1584 58608
rect 1636 58596 1642 58608
rect 1636 58568 45554 58596
rect 1636 58556 1642 58568
rect 1394 58528 1400 58540
rect 1355 58500 1400 58528
rect 1394 58488 1400 58500
rect 1452 58528 1458 58540
rect 2133 58531 2191 58537
rect 2133 58528 2145 58531
rect 1452 58500 2145 58528
rect 1452 58488 1458 58500
rect 2133 58497 2145 58500
rect 2179 58497 2191 58531
rect 2133 58491 2191 58497
rect 45526 58460 45554 58568
rect 51046 58528 51074 58636
rect 59538 58624 59544 58636
rect 59596 58624 59602 58676
rect 61286 58624 61292 58676
rect 61344 58664 61350 58676
rect 61344 58636 62252 58664
rect 61344 58624 61350 58636
rect 60274 58596 60280 58608
rect 60235 58568 60280 58596
rect 60274 58556 60280 58568
rect 60332 58556 60338 58608
rect 62114 58596 62120 58608
rect 62075 58568 62120 58596
rect 62114 58556 62120 58568
rect 62172 58556 62178 58608
rect 62224 58596 62252 58636
rect 64414 58624 64420 58676
rect 64472 58664 64478 58676
rect 65981 58667 66039 58673
rect 65981 58664 65993 58667
rect 64472 58636 65993 58664
rect 64472 58624 64478 58636
rect 65981 58633 65993 58636
rect 66027 58633 66039 58667
rect 65981 58627 66039 58633
rect 66533 58667 66591 58673
rect 66533 58633 66545 58667
rect 66579 58664 66591 58667
rect 66990 58664 66996 58676
rect 66579 58636 66996 58664
rect 66579 58633 66591 58636
rect 66533 58627 66591 58633
rect 66990 58624 66996 58636
rect 67048 58624 67054 58676
rect 77938 58664 77944 58676
rect 70366 58636 77944 58664
rect 70366 58596 70394 58636
rect 77938 58624 77944 58636
rect 77996 58624 78002 58676
rect 62224 58568 70394 58596
rect 59814 58528 59820 58540
rect 51046 58500 59820 58528
rect 59814 58488 59820 58500
rect 59872 58528 59878 58540
rect 60001 58531 60059 58537
rect 60001 58528 60013 58531
rect 59872 58500 60013 58528
rect 59872 58488 59878 58500
rect 60001 58497 60013 58500
rect 60047 58497 60059 58531
rect 60182 58528 60188 58540
rect 60143 58500 60188 58528
rect 60001 58491 60059 58497
rect 60182 58488 60188 58500
rect 60240 58488 60246 58540
rect 60366 58488 60372 58540
rect 60424 58537 60430 58540
rect 60424 58528 60432 58537
rect 60424 58500 60469 58528
rect 60424 58491 60432 58500
rect 60424 58488 60430 58491
rect 61654 58488 61660 58540
rect 61712 58528 61718 58540
rect 61841 58531 61899 58537
rect 61841 58528 61853 58531
rect 61712 58500 61853 58528
rect 61712 58488 61718 58500
rect 61841 58497 61853 58500
rect 61887 58497 61899 58531
rect 61841 58491 61899 58497
rect 61856 58460 61884 58491
rect 61930 58488 61936 58540
rect 61988 58528 61994 58540
rect 62025 58531 62083 58537
rect 62025 58528 62037 58531
rect 61988 58500 62037 58528
rect 61988 58488 61994 58500
rect 62025 58497 62037 58500
rect 62071 58497 62083 58531
rect 62025 58491 62083 58497
rect 62206 58488 62212 58540
rect 62264 58537 62270 58540
rect 62264 58528 62272 58537
rect 62264 58500 62309 58528
rect 62264 58491 62272 58500
rect 62264 58488 62270 58491
rect 63770 58488 63776 58540
rect 63828 58528 63834 58540
rect 64693 58531 64751 58537
rect 64693 58528 64705 58531
rect 63828 58500 64705 58528
rect 63828 58488 63834 58500
rect 64693 58497 64705 58500
rect 64739 58497 64751 58531
rect 64693 58491 64751 58497
rect 77297 58531 77355 58537
rect 77297 58497 77309 58531
rect 77343 58528 77355 58531
rect 77938 58528 77944 58540
rect 77343 58500 77944 58528
rect 77343 58497 77355 58500
rect 77297 58491 77355 58497
rect 77938 58488 77944 58500
rect 77996 58488 78002 58540
rect 63037 58463 63095 58469
rect 63037 58460 63049 58463
rect 45526 58432 61148 58460
rect 61856 58432 63049 58460
rect 2130 58352 2136 58404
rect 2188 58392 2194 58404
rect 61010 58392 61016 58404
rect 2188 58364 61016 58392
rect 2188 58352 2194 58364
rect 61010 58352 61016 58364
rect 61068 58352 61074 58404
rect 61120 58336 61148 58432
rect 63037 58429 63049 58432
rect 63083 58429 63095 58463
rect 63037 58423 63095 58429
rect 64874 58420 64880 58472
rect 64932 58460 64938 58472
rect 64969 58463 65027 58469
rect 64969 58460 64981 58463
rect 64932 58432 64981 58460
rect 64932 58420 64938 58432
rect 64969 58429 64981 58432
rect 65015 58460 65027 58463
rect 65429 58463 65487 58469
rect 65429 58460 65441 58463
rect 65015 58432 65441 58460
rect 65015 58429 65027 58432
rect 64969 58423 65027 58429
rect 65429 58429 65441 58432
rect 65475 58460 65487 58463
rect 65610 58460 65616 58472
rect 65475 58432 65616 58460
rect 65475 58429 65487 58432
rect 65429 58423 65487 58429
rect 65610 58420 65616 58432
rect 65668 58420 65674 58472
rect 1581 58327 1639 58333
rect 1581 58293 1593 58327
rect 1627 58324 1639 58327
rect 2682 58324 2688 58336
rect 1627 58296 2688 58324
rect 1627 58293 1639 58296
rect 1581 58287 1639 58293
rect 2682 58284 2688 58296
rect 2740 58284 2746 58336
rect 60550 58324 60556 58336
rect 60511 58296 60556 58324
rect 60550 58284 60556 58296
rect 60608 58284 60614 58336
rect 61102 58324 61108 58336
rect 61063 58296 61108 58324
rect 61102 58284 61108 58296
rect 61160 58284 61166 58336
rect 62390 58324 62396 58336
rect 62351 58296 62396 58324
rect 62390 58284 62396 58296
rect 62448 58284 62454 58336
rect 63586 58324 63592 58336
rect 63547 58296 63592 58324
rect 63586 58284 63592 58296
rect 63644 58284 63650 58336
rect 77754 58324 77760 58336
rect 77715 58296 77760 58324
rect 77754 58284 77760 58296
rect 77812 58284 77818 58336
rect 1104 58234 78844 58256
rect 1104 58182 4214 58234
rect 4266 58182 4278 58234
rect 4330 58182 4342 58234
rect 4394 58182 4406 58234
rect 4458 58182 4470 58234
rect 4522 58182 34934 58234
rect 34986 58182 34998 58234
rect 35050 58182 35062 58234
rect 35114 58182 35126 58234
rect 35178 58182 35190 58234
rect 35242 58182 65654 58234
rect 65706 58182 65718 58234
rect 65770 58182 65782 58234
rect 65834 58182 65846 58234
rect 65898 58182 65910 58234
rect 65962 58182 78844 58234
rect 1104 58160 78844 58182
rect 62206 58080 62212 58132
rect 62264 58120 62270 58132
rect 63218 58120 63224 58132
rect 62264 58092 63224 58120
rect 62264 58080 62270 58092
rect 63218 58080 63224 58092
rect 63276 58080 63282 58132
rect 61286 58052 61292 58064
rect 60844 58024 61292 58052
rect 59265 57919 59323 57925
rect 59265 57885 59277 57919
rect 59311 57885 59323 57919
rect 59538 57916 59544 57928
rect 59499 57888 59544 57916
rect 59265 57879 59323 57885
rect 2590 57808 2596 57860
rect 2648 57848 2654 57860
rect 58713 57851 58771 57857
rect 58713 57848 58725 57851
rect 2648 57820 58725 57848
rect 2648 57808 2654 57820
rect 58713 57817 58725 57820
rect 58759 57848 58771 57851
rect 59280 57848 59308 57879
rect 59538 57876 59544 57888
rect 59596 57876 59602 57928
rect 59722 57925 59728 57928
rect 59685 57919 59728 57925
rect 59685 57885 59697 57919
rect 59780 57916 59786 57928
rect 60366 57916 60372 57928
rect 59780 57888 60372 57916
rect 59685 57879 59728 57885
rect 59722 57876 59728 57879
rect 59780 57876 59786 57888
rect 60366 57876 60372 57888
rect 60424 57916 60430 57928
rect 60844 57925 60872 58024
rect 61286 58012 61292 58024
rect 61344 58012 61350 58064
rect 63586 58052 63592 58064
rect 62868 58024 63592 58052
rect 61010 57944 61016 57996
rect 61068 57984 61074 57996
rect 62868 57984 62896 58024
rect 63586 58012 63592 58024
rect 63644 58012 63650 58064
rect 61068 57956 62896 57984
rect 61068 57944 61074 57956
rect 60685 57919 60743 57925
rect 60685 57916 60697 57919
rect 60424 57888 60697 57916
rect 60424 57876 60430 57888
rect 60685 57885 60697 57888
rect 60731 57885 60743 57919
rect 60685 57879 60743 57885
rect 60829 57919 60887 57925
rect 60829 57885 60841 57919
rect 60875 57885 60887 57919
rect 61102 57916 61108 57928
rect 61063 57888 61108 57916
rect 60829 57879 60887 57885
rect 61102 57876 61108 57888
rect 61160 57876 61166 57928
rect 61746 57916 61752 57928
rect 61707 57888 61752 57916
rect 61746 57876 61752 57888
rect 61804 57876 61810 57928
rect 62114 57876 62120 57928
rect 62172 57925 62178 57928
rect 62172 57916 62180 57925
rect 62172 57888 62217 57916
rect 62172 57879 62180 57888
rect 62172 57876 62178 57879
rect 62298 57876 62304 57928
rect 62356 57925 62362 57928
rect 62868 57925 62896 57956
rect 63144 57956 63448 57984
rect 63880 57974 64092 57984
rect 62356 57919 62376 57925
rect 62364 57885 62376 57919
rect 62356 57879 62376 57885
rect 62853 57919 62911 57925
rect 62853 57885 62865 57919
rect 62899 57885 62911 57919
rect 63144 57916 63172 57956
rect 62853 57879 62911 57885
rect 62960 57888 63172 57916
rect 62356 57876 62362 57879
rect 58759 57820 59308 57848
rect 59449 57851 59507 57857
rect 58759 57817 58771 57820
rect 58713 57811 58771 57817
rect 59449 57817 59461 57851
rect 59495 57848 59507 57851
rect 60182 57848 60188 57860
rect 59495 57820 60188 57848
rect 59495 57817 59507 57820
rect 59449 57811 59507 57817
rect 59556 57792 59584 57820
rect 60182 57808 60188 57820
rect 60240 57848 60246 57860
rect 60458 57848 60464 57860
rect 60240 57820 60464 57848
rect 60240 57808 60246 57820
rect 60458 57808 60464 57820
rect 60516 57848 60522 57860
rect 60921 57851 60979 57857
rect 60516 57820 60780 57848
rect 60516 57808 60522 57820
rect 1394 57780 1400 57792
rect 1355 57752 1400 57780
rect 1394 57740 1400 57752
rect 1452 57740 1458 57792
rect 59538 57740 59544 57792
rect 59596 57740 59602 57792
rect 59814 57780 59820 57792
rect 59872 57789 59878 57792
rect 59783 57752 59820 57780
rect 59814 57740 59820 57752
rect 59872 57743 59883 57789
rect 60545 57783 60603 57789
rect 60545 57749 60557 57783
rect 60591 57780 60603 57783
rect 60642 57780 60648 57792
rect 60591 57752 60648 57780
rect 60591 57749 60603 57752
rect 60545 57743 60603 57749
rect 59872 57740 59878 57743
rect 60642 57740 60648 57752
rect 60700 57740 60706 57792
rect 60752 57780 60780 57820
rect 60921 57817 60933 57851
rect 60967 57817 60979 57851
rect 60921 57811 60979 57817
rect 60936 57780 60964 57811
rect 61378 57808 61384 57860
rect 61436 57848 61442 57860
rect 61930 57848 61936 57860
rect 61436 57820 61936 57848
rect 61436 57808 61442 57820
rect 61930 57808 61936 57820
rect 61988 57808 61994 57860
rect 62025 57851 62083 57857
rect 62025 57817 62037 57851
rect 62071 57848 62083 57851
rect 62960 57848 62988 57888
rect 63218 57876 63224 57928
rect 63276 57925 63282 57928
rect 63276 57916 63284 57925
rect 63420 57916 63448 57956
rect 63696 57956 64092 57974
rect 63696 57946 63908 57956
rect 63586 57916 63592 57928
rect 63276 57888 63321 57916
rect 63420 57888 63592 57916
rect 63276 57879 63284 57888
rect 63276 57876 63282 57879
rect 63586 57876 63592 57888
rect 63644 57876 63650 57928
rect 62071 57820 62988 57848
rect 63037 57851 63095 57857
rect 62071 57817 62083 57820
rect 62025 57811 62083 57817
rect 63037 57817 63049 57851
rect 63083 57817 63095 57851
rect 63037 57811 63095 57817
rect 63129 57851 63187 57857
rect 63129 57817 63141 57851
rect 63175 57848 63187 57851
rect 63696 57848 63724 57946
rect 63175 57820 63724 57848
rect 64064 57848 64092 57956
rect 65334 57876 65340 57928
rect 65392 57916 65398 57928
rect 65613 57919 65671 57925
rect 65613 57916 65625 57919
rect 65392 57888 65625 57916
rect 65392 57876 65398 57888
rect 65613 57885 65625 57888
rect 65659 57885 65671 57919
rect 65613 57879 65671 57885
rect 64601 57851 64659 57857
rect 64601 57848 64613 57851
rect 64064 57820 64613 57848
rect 63175 57817 63187 57820
rect 63129 57811 63187 57817
rect 64601 57817 64613 57820
rect 64647 57848 64659 57851
rect 77294 57848 77300 57860
rect 64647 57820 77300 57848
rect 64647 57817 64659 57820
rect 64601 57811 64659 57817
rect 60752 57752 60964 57780
rect 61948 57780 61976 57808
rect 63052 57780 63080 57811
rect 77294 57808 77300 57820
rect 77352 57808 77358 57860
rect 63218 57780 63224 57792
rect 61948 57752 63224 57780
rect 63218 57740 63224 57752
rect 63276 57740 63282 57792
rect 63310 57740 63316 57792
rect 63368 57780 63374 57792
rect 63413 57783 63471 57789
rect 63413 57780 63425 57783
rect 63368 57752 63425 57780
rect 63368 57740 63374 57752
rect 63413 57749 63425 57752
rect 63459 57749 63471 57783
rect 63413 57743 63471 57749
rect 63586 57740 63592 57792
rect 63644 57780 63650 57792
rect 64049 57783 64107 57789
rect 64049 57780 64061 57783
rect 63644 57752 64061 57780
rect 63644 57740 63650 57752
rect 64049 57749 64061 57752
rect 64095 57780 64107 57783
rect 77478 57780 77484 57792
rect 64095 57752 77484 57780
rect 64095 57749 64107 57752
rect 64049 57743 64107 57749
rect 77478 57740 77484 57752
rect 77536 57740 77542 57792
rect 77938 57740 77944 57792
rect 77996 57780 78002 57792
rect 78033 57783 78091 57789
rect 78033 57780 78045 57783
rect 77996 57752 78045 57780
rect 77996 57740 78002 57752
rect 78033 57749 78045 57752
rect 78079 57749 78091 57783
rect 78033 57743 78091 57749
rect 1104 57690 78844 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 78844 57690
rect 1104 57616 78844 57638
rect 1486 57536 1492 57588
rect 1544 57576 1550 57588
rect 1544 57548 59492 57576
rect 1544 57536 1550 57548
rect 1394 57440 1400 57452
rect 1355 57412 1400 57440
rect 1394 57400 1400 57412
rect 1452 57400 1458 57452
rect 59357 57443 59415 57449
rect 59357 57440 59369 57443
rect 58820 57412 59369 57440
rect 58820 57313 58848 57412
rect 59357 57409 59369 57412
rect 59403 57409 59415 57443
rect 59357 57403 59415 57409
rect 59464 57372 59492 57548
rect 59630 57508 59636 57520
rect 59591 57480 59636 57508
rect 59630 57468 59636 57480
rect 59688 57508 59694 57520
rect 77754 57508 77760 57520
rect 59688 57480 77760 57508
rect 59688 57468 59694 57480
rect 77754 57468 77760 57480
rect 77812 57468 77818 57520
rect 59538 57400 59544 57452
rect 59596 57440 59602 57452
rect 59596 57412 59641 57440
rect 59596 57400 59602 57412
rect 59722 57400 59728 57452
rect 59780 57449 59786 57452
rect 59780 57440 59788 57449
rect 61746 57440 61752 57452
rect 59780 57412 59825 57440
rect 60706 57412 61752 57440
rect 59780 57403 59788 57412
rect 59780 57400 59786 57403
rect 60706 57372 60734 57412
rect 61746 57400 61752 57412
rect 61804 57440 61810 57452
rect 62117 57443 62175 57449
rect 62117 57440 62129 57443
rect 61804 57412 62129 57440
rect 61804 57400 61810 57412
rect 62117 57409 62129 57412
rect 62163 57409 62175 57443
rect 63034 57440 63040 57452
rect 62995 57412 63040 57440
rect 62117 57403 62175 57409
rect 63034 57400 63040 57412
rect 63092 57400 63098 57452
rect 63218 57440 63224 57452
rect 63179 57412 63224 57440
rect 63218 57400 63224 57412
rect 63276 57400 63282 57452
rect 63313 57443 63371 57449
rect 63313 57409 63325 57443
rect 63359 57409 63371 57443
rect 63313 57403 63371 57409
rect 61378 57372 61384 57384
rect 59464 57344 60734 57372
rect 61339 57344 61384 57372
rect 61378 57332 61384 57344
rect 61436 57332 61442 57384
rect 61657 57375 61715 57381
rect 61657 57341 61669 57375
rect 61703 57341 61715 57375
rect 63328 57372 63356 57403
rect 63402 57400 63408 57452
rect 63460 57449 63466 57452
rect 63460 57440 63468 57449
rect 77938 57440 77944 57452
rect 63460 57412 63505 57440
rect 77899 57412 77944 57440
rect 63460 57403 63468 57412
rect 63460 57400 63466 57403
rect 77938 57400 77944 57412
rect 77996 57400 78002 57452
rect 64233 57375 64291 57381
rect 64233 57372 64245 57375
rect 63328 57344 64245 57372
rect 61657 57335 61715 57341
rect 64233 57341 64245 57344
rect 64279 57372 64291 57375
rect 64279 57344 70394 57372
rect 64279 57341 64291 57344
rect 64233 57335 64291 57341
rect 58805 57307 58863 57313
rect 58805 57304 58817 57307
rect 51046 57276 58817 57304
rect 1578 57236 1584 57248
rect 1539 57208 1584 57236
rect 1578 57196 1584 57208
rect 1636 57196 1642 57248
rect 2682 57196 2688 57248
rect 2740 57236 2746 57248
rect 51046 57236 51074 57276
rect 58805 57273 58817 57276
rect 58851 57273 58863 57307
rect 58805 57267 58863 57273
rect 60826 57264 60832 57316
rect 60884 57304 60890 57316
rect 61672 57304 61700 57335
rect 60884 57276 61700 57304
rect 63589 57307 63647 57313
rect 60884 57264 60890 57276
rect 63589 57273 63601 57307
rect 63635 57304 63647 57307
rect 64322 57304 64328 57316
rect 63635 57276 64328 57304
rect 63635 57273 63647 57276
rect 63589 57267 63647 57273
rect 64322 57264 64328 57276
rect 64380 57264 64386 57316
rect 70366 57304 70394 57344
rect 77386 57304 77392 57316
rect 70366 57276 77392 57304
rect 77386 57264 77392 57276
rect 77444 57264 77450 57316
rect 2740 57208 51074 57236
rect 58345 57239 58403 57245
rect 2740 57196 2746 57208
rect 58345 57205 58357 57239
rect 58391 57236 58403 57239
rect 59630 57236 59636 57248
rect 58391 57208 59636 57236
rect 58391 57205 58403 57208
rect 58345 57199 58403 57205
rect 59630 57196 59636 57208
rect 59688 57196 59694 57248
rect 59909 57239 59967 57245
rect 59909 57205 59921 57239
rect 59955 57236 59967 57239
rect 60274 57236 60280 57248
rect 59955 57208 60280 57236
rect 59955 57205 59967 57208
rect 59909 57199 59967 57205
rect 60274 57196 60280 57208
rect 60332 57196 60338 57248
rect 77754 57236 77760 57248
rect 77715 57208 77760 57236
rect 77754 57196 77760 57208
rect 77812 57196 77818 57248
rect 1104 57146 78844 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 78844 57146
rect 1104 57072 78844 57094
rect 63034 57032 63040 57044
rect 45526 57004 63040 57032
rect 1946 56856 1952 56908
rect 2004 56896 2010 56908
rect 45526 56896 45554 57004
rect 63034 56992 63040 57004
rect 63092 56992 63098 57044
rect 77754 57032 77760 57044
rect 70366 57004 77760 57032
rect 59814 56964 59820 56976
rect 59775 56936 59820 56964
rect 59814 56924 59820 56936
rect 59872 56924 59878 56976
rect 60458 56924 60464 56976
rect 60516 56964 60522 56976
rect 60516 56936 60780 56964
rect 60516 56924 60522 56936
rect 2004 56868 45554 56896
rect 2004 56856 2010 56868
rect 59078 56856 59084 56908
rect 59136 56896 59142 56908
rect 60752 56905 60780 56936
rect 60737 56899 60795 56905
rect 59136 56868 60596 56896
rect 59136 56856 59142 56868
rect 1394 56828 1400 56840
rect 1355 56800 1400 56828
rect 1394 56788 1400 56800
rect 1452 56828 1458 56840
rect 2133 56831 2191 56837
rect 2133 56828 2145 56831
rect 1452 56800 2145 56828
rect 1452 56788 1458 56800
rect 2133 56797 2145 56800
rect 2179 56797 2191 56831
rect 2133 56791 2191 56797
rect 59265 56831 59323 56837
rect 59265 56797 59277 56831
rect 59311 56797 59323 56831
rect 59446 56828 59452 56840
rect 59407 56800 59452 56828
rect 59265 56791 59323 56797
rect 2038 56720 2044 56772
rect 2096 56760 2102 56772
rect 58713 56763 58771 56769
rect 58713 56760 58725 56763
rect 2096 56732 58725 56760
rect 2096 56720 2102 56732
rect 58713 56729 58725 56732
rect 58759 56760 58771 56763
rect 59280 56760 59308 56791
rect 59446 56788 59452 56800
rect 59504 56788 59510 56840
rect 59722 56837 59728 56840
rect 59685 56831 59728 56837
rect 59685 56797 59697 56831
rect 59685 56791 59728 56797
rect 59722 56788 59728 56791
rect 59780 56788 59786 56840
rect 60461 56831 60519 56837
rect 60461 56797 60473 56831
rect 60507 56797 60519 56831
rect 60568 56828 60596 56868
rect 60737 56865 60749 56899
rect 60783 56865 60795 56899
rect 70366 56896 70394 57004
rect 77754 56992 77760 57004
rect 77812 56992 77818 57044
rect 60737 56859 60795 56865
rect 61672 56868 70394 56896
rect 61672 56828 61700 56868
rect 60568 56800 61700 56828
rect 61749 56831 61807 56837
rect 60461 56791 60519 56797
rect 61749 56797 61761 56831
rect 61795 56797 61807 56831
rect 61749 56791 61807 56797
rect 62025 56831 62083 56837
rect 62025 56797 62037 56831
rect 62071 56828 62083 56831
rect 62114 56828 62120 56840
rect 62071 56800 62120 56828
rect 62071 56797 62083 56800
rect 62025 56791 62083 56797
rect 58759 56732 59308 56760
rect 58759 56729 58771 56732
rect 58713 56723 58771 56729
rect 59538 56720 59544 56772
rect 59596 56760 59602 56772
rect 59998 56760 60004 56772
rect 59596 56732 60004 56760
rect 59596 56720 59602 56732
rect 59998 56720 60004 56732
rect 60056 56720 60062 56772
rect 1581 56695 1639 56701
rect 1581 56661 1593 56695
rect 1627 56692 1639 56695
rect 2682 56692 2688 56704
rect 1627 56664 2688 56692
rect 1627 56661 1639 56664
rect 1581 56655 1639 56661
rect 2682 56652 2688 56664
rect 2740 56652 2746 56704
rect 60476 56692 60504 56791
rect 60734 56720 60740 56772
rect 60792 56760 60798 56772
rect 61764 56760 61792 56791
rect 62114 56788 62120 56800
rect 62172 56788 62178 56840
rect 77481 56831 77539 56837
rect 77481 56797 77493 56831
rect 77527 56828 77539 56831
rect 78122 56828 78128 56840
rect 77527 56800 78128 56828
rect 77527 56797 77539 56800
rect 77481 56791 77539 56797
rect 78122 56788 78128 56800
rect 78180 56788 78186 56840
rect 60792 56732 61792 56760
rect 60792 56720 60798 56732
rect 60826 56692 60832 56704
rect 60476 56664 60832 56692
rect 60826 56652 60832 56664
rect 60884 56652 60890 56704
rect 76190 56652 76196 56704
rect 76248 56692 76254 56704
rect 77941 56695 77999 56701
rect 77941 56692 77953 56695
rect 76248 56664 77953 56692
rect 76248 56652 76254 56664
rect 77941 56661 77953 56664
rect 77987 56661 77999 56695
rect 77941 56655 77999 56661
rect 1104 56602 78844 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 78844 56602
rect 1104 56528 78844 56550
rect 1578 56448 1584 56500
rect 1636 56488 1642 56500
rect 57698 56488 57704 56500
rect 1636 56460 57704 56488
rect 1636 56448 1642 56460
rect 57698 56448 57704 56460
rect 57756 56448 57762 56500
rect 59449 56491 59507 56497
rect 59449 56457 59461 56491
rect 59495 56488 59507 56491
rect 59538 56488 59544 56500
rect 59495 56460 59544 56488
rect 59495 56457 59507 56460
rect 59449 56451 59507 56457
rect 59538 56448 59544 56460
rect 59596 56448 59602 56500
rect 57882 56380 57888 56432
rect 57940 56420 57946 56432
rect 58529 56423 58587 56429
rect 58529 56420 58541 56423
rect 57940 56392 58541 56420
rect 57940 56380 57946 56392
rect 58529 56389 58541 56392
rect 58575 56420 58587 56423
rect 58575 56392 60734 56420
rect 58575 56389 58587 56392
rect 58529 56383 58587 56389
rect 1394 56352 1400 56364
rect 1355 56324 1400 56352
rect 1394 56312 1400 56324
rect 1452 56352 1458 56364
rect 2133 56355 2191 56361
rect 2133 56352 2145 56355
rect 1452 56324 2145 56352
rect 1452 56312 1458 56324
rect 2133 56321 2145 56324
rect 2179 56321 2191 56355
rect 2133 56315 2191 56321
rect 59722 56312 59728 56364
rect 59780 56352 59786 56364
rect 60461 56355 60519 56361
rect 60461 56352 60473 56355
rect 59780 56324 60473 56352
rect 59780 56312 59786 56324
rect 60461 56321 60473 56324
rect 60507 56321 60519 56355
rect 60706 56352 60734 56392
rect 76190 56352 76196 56364
rect 60706 56324 76196 56352
rect 60461 56315 60519 56321
rect 76190 56312 76196 56324
rect 76248 56312 76254 56364
rect 77297 56355 77355 56361
rect 77297 56321 77309 56355
rect 77343 56352 77355 56355
rect 77938 56352 77944 56364
rect 77343 56324 77944 56352
rect 77343 56321 77355 56324
rect 77297 56315 77355 56321
rect 77938 56312 77944 56324
rect 77996 56312 78002 56364
rect 60734 56244 60740 56296
rect 60792 56284 60798 56296
rect 61194 56284 61200 56296
rect 60792 56256 60837 56284
rect 61155 56256 61200 56284
rect 60792 56244 60798 56256
rect 61194 56244 61200 56256
rect 61252 56284 61258 56296
rect 63126 56284 63132 56296
rect 61252 56256 63132 56284
rect 61252 56244 61258 56256
rect 63126 56244 63132 56256
rect 63184 56244 63190 56296
rect 1581 56219 1639 56225
rect 1581 56185 1593 56219
rect 1627 56216 1639 56219
rect 55950 56216 55956 56228
rect 1627 56188 55956 56216
rect 1627 56185 1639 56188
rect 1581 56179 1639 56185
rect 55950 56176 55956 56188
rect 56008 56176 56014 56228
rect 56778 56176 56784 56228
rect 56836 56216 56842 56228
rect 57977 56219 58035 56225
rect 57977 56216 57989 56219
rect 56836 56188 57989 56216
rect 56836 56176 56842 56188
rect 57977 56185 57989 56188
rect 58023 56216 58035 56219
rect 77757 56219 77815 56225
rect 77757 56216 77769 56219
rect 58023 56188 77769 56216
rect 58023 56185 58035 56188
rect 57977 56179 58035 56185
rect 77757 56185 77769 56188
rect 77803 56185 77815 56219
rect 77757 56179 77815 56185
rect 57057 56151 57115 56157
rect 57057 56117 57069 56151
rect 57103 56148 57115 56151
rect 57146 56148 57152 56160
rect 57103 56120 57152 56148
rect 57103 56117 57115 56120
rect 57057 56111 57115 56117
rect 57146 56108 57152 56120
rect 57204 56108 57210 56160
rect 60826 56108 60832 56160
rect 60884 56148 60890 56160
rect 61427 56151 61485 56157
rect 61427 56148 61439 56151
rect 60884 56120 61439 56148
rect 60884 56108 60890 56120
rect 61427 56117 61439 56120
rect 61473 56117 61485 56151
rect 61427 56111 61485 56117
rect 1104 56058 78844 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 78844 56058
rect 1104 55984 78844 56006
rect 55950 55944 55956 55956
rect 55911 55916 55956 55944
rect 55950 55904 55956 55916
rect 56008 55904 56014 55956
rect 57146 55904 57152 55956
rect 57204 55944 57210 55956
rect 77941 55947 77999 55953
rect 77941 55944 77953 55947
rect 57204 55916 77953 55944
rect 57204 55904 57210 55916
rect 77941 55913 77953 55916
rect 77987 55913 77999 55947
rect 77941 55907 77999 55913
rect 45526 55780 51074 55808
rect 2682 55700 2688 55752
rect 2740 55740 2746 55752
rect 45526 55740 45554 55780
rect 2740 55712 45554 55740
rect 2740 55700 2746 55712
rect 1486 55672 1492 55684
rect 1447 55644 1492 55672
rect 1486 55632 1492 55644
rect 1544 55632 1550 55684
rect 1673 55675 1731 55681
rect 1673 55641 1685 55675
rect 1719 55672 1731 55675
rect 51046 55672 51074 55780
rect 55968 55740 55996 55904
rect 57054 55876 57060 55888
rect 57015 55848 57060 55876
rect 57054 55836 57060 55848
rect 57112 55836 57118 55888
rect 58161 55879 58219 55885
rect 58161 55845 58173 55879
rect 58207 55876 58219 55879
rect 58434 55876 58440 55888
rect 58207 55848 58440 55876
rect 58207 55845 58219 55848
rect 58161 55839 58219 55845
rect 58434 55836 58440 55848
rect 58492 55836 58498 55888
rect 60734 55836 60740 55888
rect 60792 55876 60798 55888
rect 60792 55848 61056 55876
rect 60792 55836 60798 55848
rect 61028 55817 61056 55848
rect 58713 55811 58771 55817
rect 58713 55808 58725 55811
rect 56612 55780 58725 55808
rect 56505 55743 56563 55749
rect 56505 55740 56517 55743
rect 55968 55712 56517 55740
rect 56505 55709 56517 55712
rect 56551 55709 56563 55743
rect 56505 55703 56563 55709
rect 56612 55672 56640 55780
rect 56778 55740 56784 55752
rect 56739 55712 56784 55740
rect 56778 55700 56784 55712
rect 56836 55700 56842 55752
rect 56870 55700 56876 55752
rect 56928 55749 56934 55752
rect 57624 55749 57652 55780
rect 58713 55777 58725 55780
rect 58759 55777 58771 55811
rect 58713 55771 58771 55777
rect 61013 55811 61071 55817
rect 61013 55777 61025 55811
rect 61059 55777 61071 55811
rect 61013 55771 61071 55777
rect 56928 55740 56936 55749
rect 57609 55743 57667 55749
rect 56928 55712 56973 55740
rect 56928 55703 56936 55712
rect 57609 55709 57621 55743
rect 57655 55709 57667 55743
rect 57882 55740 57888 55752
rect 57843 55712 57888 55740
rect 57609 55703 57667 55709
rect 56928 55700 56934 55703
rect 57882 55700 57888 55712
rect 57940 55700 57946 55752
rect 57982 55743 58040 55749
rect 57982 55709 57994 55743
rect 58028 55709 58040 55743
rect 57982 55703 58040 55709
rect 1719 55644 6914 55672
rect 51046 55644 56640 55672
rect 56689 55675 56747 55681
rect 1719 55641 1731 55644
rect 1673 55635 1731 55641
rect 1504 55604 1532 55632
rect 2133 55607 2191 55613
rect 2133 55604 2145 55607
rect 1504 55576 2145 55604
rect 2133 55573 2145 55576
rect 2179 55573 2191 55607
rect 6886 55604 6914 55644
rect 56689 55641 56701 55675
rect 56735 55672 56747 55675
rect 57790 55672 57796 55684
rect 56735 55644 57796 55672
rect 56735 55641 56747 55644
rect 56689 55635 56747 55641
rect 55674 55604 55680 55616
rect 6886 55576 55680 55604
rect 2133 55567 2191 55573
rect 55674 55564 55680 55576
rect 55732 55564 55738 55616
rect 56594 55564 56600 55616
rect 56652 55604 56658 55616
rect 56704 55604 56732 55635
rect 57790 55632 57796 55644
rect 57848 55632 57854 55684
rect 56652 55576 56732 55604
rect 56652 55564 56658 55576
rect 56870 55564 56876 55616
rect 56928 55604 56934 55616
rect 57882 55604 57888 55616
rect 56928 55576 57888 55604
rect 56928 55564 56934 55576
rect 57882 55564 57888 55576
rect 57940 55604 57946 55616
rect 57992 55604 58020 55703
rect 60458 55700 60464 55752
rect 60516 55740 60522 55752
rect 60737 55743 60795 55749
rect 60737 55740 60749 55743
rect 60516 55712 60749 55740
rect 60516 55700 60522 55712
rect 60737 55709 60749 55712
rect 60783 55740 60795 55743
rect 64874 55740 64880 55752
rect 60783 55712 64880 55740
rect 60783 55709 60795 55712
rect 60737 55703 60795 55709
rect 64874 55700 64880 55712
rect 64932 55700 64938 55752
rect 77481 55743 77539 55749
rect 77481 55709 77493 55743
rect 77527 55740 77539 55743
rect 78122 55740 78128 55752
rect 77527 55712 78128 55740
rect 77527 55709 77539 55712
rect 77481 55703 77539 55709
rect 78122 55700 78128 55712
rect 78180 55700 78186 55752
rect 57940 55576 58020 55604
rect 57940 55564 57946 55576
rect 1104 55514 78844 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 78844 55514
rect 1104 55440 78844 55462
rect 55674 55400 55680 55412
rect 55635 55372 55680 55400
rect 55674 55360 55680 55372
rect 55732 55360 55738 55412
rect 57882 55360 57888 55412
rect 57940 55400 57946 55412
rect 57940 55372 58296 55400
rect 57940 55360 57946 55372
rect 55692 55264 55720 55360
rect 56505 55335 56563 55341
rect 56505 55301 56517 55335
rect 56551 55332 56563 55335
rect 57146 55332 57152 55344
rect 56551 55304 57152 55332
rect 56551 55301 56563 55304
rect 56505 55295 56563 55301
rect 57146 55292 57152 55304
rect 57204 55292 57210 55344
rect 57790 55292 57796 55344
rect 57848 55332 57854 55344
rect 58069 55335 58127 55341
rect 58069 55332 58081 55335
rect 57848 55304 58081 55332
rect 57848 55292 57854 55304
rect 58069 55301 58081 55304
rect 58115 55301 58127 55335
rect 58069 55295 58127 55301
rect 56686 55273 56692 55276
rect 56229 55267 56287 55273
rect 56229 55264 56241 55267
rect 55692 55236 56241 55264
rect 56229 55233 56241 55236
rect 56275 55233 56287 55267
rect 56229 55227 56287 55233
rect 56413 55267 56471 55273
rect 56413 55233 56425 55267
rect 56459 55233 56471 55267
rect 56413 55227 56471 55233
rect 56649 55267 56692 55273
rect 56649 55233 56661 55267
rect 56649 55227 56692 55233
rect 56428 55196 56456 55227
rect 56686 55224 56692 55227
rect 56744 55224 56750 55276
rect 57698 55224 57704 55276
rect 57756 55264 57762 55276
rect 58268 55273 58296 55372
rect 57885 55267 57943 55273
rect 57885 55264 57897 55267
rect 57756 55236 57897 55264
rect 57756 55224 57762 55236
rect 57885 55233 57897 55236
rect 57931 55264 57943 55267
rect 58161 55267 58219 55273
rect 57931 55236 58112 55264
rect 57931 55233 57943 55236
rect 57885 55227 57943 55233
rect 56428 55168 56640 55196
rect 56612 55140 56640 55168
rect 56594 55088 56600 55140
rect 56652 55088 56658 55140
rect 58084 55128 58112 55236
rect 58161 55233 58173 55267
rect 58207 55233 58219 55267
rect 58161 55227 58219 55233
rect 58258 55267 58316 55273
rect 58258 55233 58270 55267
rect 58304 55233 58316 55267
rect 58258 55227 58316 55233
rect 58454 55267 58512 55273
rect 58454 55233 58466 55267
rect 58500 55264 58512 55267
rect 58986 55264 58992 55276
rect 58500 55236 58992 55264
rect 58500 55233 58512 55236
rect 58454 55227 58512 55233
rect 58176 55196 58204 55227
rect 58986 55224 58992 55236
rect 59044 55224 59050 55276
rect 60458 55224 60464 55276
rect 60516 55264 60522 55276
rect 60553 55267 60611 55273
rect 60553 55264 60565 55267
rect 60516 55236 60565 55264
rect 60516 55224 60522 55236
rect 60553 55233 60565 55236
rect 60599 55233 60611 55267
rect 61194 55264 61200 55276
rect 61155 55236 61200 55264
rect 60553 55227 60611 55233
rect 61194 55224 61200 55236
rect 61252 55224 61258 55276
rect 59078 55196 59084 55208
rect 58176 55168 59084 55196
rect 59078 55156 59084 55168
rect 59136 55156 59142 55208
rect 58989 55131 59047 55137
rect 58989 55128 59001 55131
rect 58084 55100 59001 55128
rect 58989 55097 59001 55100
rect 59035 55097 59047 55131
rect 58989 55091 59047 55097
rect 1486 55060 1492 55072
rect 1447 55032 1492 55060
rect 1486 55020 1492 55032
rect 1544 55020 1550 55072
rect 56781 55063 56839 55069
rect 56781 55029 56793 55063
rect 56827 55060 56839 55063
rect 57146 55060 57152 55072
rect 56827 55032 57152 55060
rect 56827 55029 56839 55032
rect 56781 55023 56839 55029
rect 57146 55020 57152 55032
rect 57204 55020 57210 55072
rect 77941 55063 77999 55069
rect 77941 55029 77953 55063
rect 77987 55060 77999 55063
rect 78122 55060 78128 55072
rect 77987 55032 78128 55060
rect 77987 55029 77999 55032
rect 77941 55023 77999 55029
rect 78122 55020 78128 55032
rect 78180 55020 78186 55072
rect 1104 54970 78844 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 78844 54970
rect 1104 54896 78844 54918
rect 58989 54859 59047 54865
rect 58989 54825 59001 54859
rect 59035 54856 59047 54859
rect 59078 54856 59084 54868
rect 59035 54828 59084 54856
rect 59035 54825 59047 54828
rect 58989 54819 59047 54825
rect 59078 54816 59084 54828
rect 59136 54816 59142 54868
rect 60826 54788 60832 54800
rect 56336 54760 60832 54788
rect 53098 54680 53104 54732
rect 53156 54720 53162 54732
rect 56336 54729 56364 54760
rect 60826 54748 60832 54760
rect 60884 54748 60890 54800
rect 56321 54723 56379 54729
rect 56321 54720 56333 54723
rect 53156 54692 56333 54720
rect 53156 54680 53162 54692
rect 56321 54689 56333 54692
rect 56367 54689 56379 54723
rect 56321 54683 56379 54689
rect 56686 54680 56692 54732
rect 56744 54720 56750 54732
rect 57885 54723 57943 54729
rect 57885 54720 57897 54723
rect 56744 54692 57897 54720
rect 56744 54680 56750 54692
rect 57885 54689 57897 54692
rect 57931 54689 57943 54723
rect 57885 54683 57943 54689
rect 1486 54652 1492 54664
rect 1447 54624 1492 54652
rect 1486 54612 1492 54624
rect 1544 54612 1550 54664
rect 56594 54652 56600 54664
rect 56555 54624 56600 54652
rect 56594 54612 56600 54624
rect 56652 54612 56658 54664
rect 57609 54655 57667 54661
rect 57609 54621 57621 54655
rect 57655 54652 57667 54655
rect 60734 54652 60740 54664
rect 57655 54624 60740 54652
rect 57655 54621 57667 54624
rect 57609 54615 57667 54621
rect 53374 54544 53380 54596
rect 53432 54584 53438 54596
rect 57624 54584 57652 54615
rect 60734 54612 60740 54624
rect 60792 54612 60798 54664
rect 77481 54655 77539 54661
rect 77481 54621 77493 54655
rect 77527 54652 77539 54655
rect 77938 54652 77944 54664
rect 77527 54624 77944 54652
rect 77527 54621 77539 54624
rect 77481 54615 77539 54621
rect 77938 54612 77944 54624
rect 77996 54612 78002 54664
rect 78122 54652 78128 54664
rect 78083 54624 78128 54652
rect 78122 54612 78128 54624
rect 78180 54612 78186 54664
rect 53432 54556 57652 54584
rect 53432 54544 53438 54556
rect 1581 54519 1639 54525
rect 1581 54485 1593 54519
rect 1627 54516 1639 54519
rect 55490 54516 55496 54528
rect 1627 54488 55496 54516
rect 1627 54485 1639 54488
rect 1581 54479 1639 54485
rect 55490 54476 55496 54488
rect 55548 54476 55554 54528
rect 76190 54476 76196 54528
rect 76248 54516 76254 54528
rect 77941 54519 77999 54525
rect 77941 54516 77953 54519
rect 76248 54488 77953 54516
rect 76248 54476 76254 54488
rect 77941 54485 77953 54488
rect 77987 54485 77999 54519
rect 77941 54479 77999 54485
rect 1104 54426 78844 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 78844 54426
rect 1104 54352 78844 54374
rect 55490 54312 55496 54324
rect 55451 54284 55496 54312
rect 55490 54272 55496 54284
rect 55548 54272 55554 54324
rect 1486 54176 1492 54188
rect 1447 54148 1492 54176
rect 1486 54136 1492 54148
rect 1544 54176 1550 54188
rect 2133 54179 2191 54185
rect 2133 54176 2145 54179
rect 1544 54148 2145 54176
rect 1544 54136 1550 54148
rect 2133 54145 2145 54148
rect 2179 54145 2191 54179
rect 55508 54176 55536 54272
rect 56229 54247 56287 54253
rect 56229 54213 56241 54247
rect 56275 54244 56287 54247
rect 56594 54244 56600 54256
rect 56275 54216 56600 54244
rect 56275 54213 56287 54216
rect 56229 54207 56287 54213
rect 56594 54204 56600 54216
rect 56652 54204 56658 54256
rect 56045 54179 56103 54185
rect 56045 54176 56057 54179
rect 55508 54148 56057 54176
rect 2133 54139 2191 54145
rect 56045 54145 56057 54148
rect 56091 54145 56103 54179
rect 56045 54139 56103 54145
rect 56321 54179 56379 54185
rect 56321 54145 56333 54179
rect 56367 54145 56379 54179
rect 56321 54139 56379 54145
rect 56465 54179 56523 54185
rect 56465 54145 56477 54179
rect 56511 54176 56523 54179
rect 56686 54176 56692 54188
rect 56511 54148 56692 54176
rect 56511 54145 56523 54148
rect 56465 54139 56523 54145
rect 56336 54108 56364 54139
rect 56686 54136 56692 54148
rect 56744 54136 56750 54188
rect 56336 54080 57284 54108
rect 1670 54040 1676 54052
rect 1631 54012 1676 54040
rect 1670 54000 1676 54012
rect 1728 54000 1734 54052
rect 56594 53972 56600 53984
rect 56555 53944 56600 53972
rect 56594 53932 56600 53944
rect 56652 53932 56658 53984
rect 57256 53981 57284 54080
rect 77478 54068 77484 54120
rect 77536 54108 77542 54120
rect 77665 54111 77723 54117
rect 77665 54108 77677 54111
rect 77536 54080 77677 54108
rect 77536 54068 77542 54080
rect 77665 54077 77677 54080
rect 77711 54077 77723 54111
rect 77938 54108 77944 54120
rect 77899 54080 77944 54108
rect 77665 54071 77723 54077
rect 77938 54068 77944 54080
rect 77996 54068 78002 54120
rect 57241 53975 57299 53981
rect 57241 53941 57253 53975
rect 57287 53972 57299 53975
rect 76190 53972 76196 53984
rect 57287 53944 76196 53972
rect 57287 53941 57299 53944
rect 57241 53935 57299 53941
rect 76190 53932 76196 53944
rect 76248 53932 76254 53984
rect 1104 53882 78844 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 78844 53882
rect 1104 53808 78844 53830
rect 76837 53567 76895 53573
rect 76837 53533 76849 53567
rect 76883 53564 76895 53567
rect 77294 53564 77300 53576
rect 76883 53536 77300 53564
rect 76883 53533 76895 53536
rect 76837 53527 76895 53533
rect 77294 53524 77300 53536
rect 77352 53524 77358 53576
rect 77386 53524 77392 53576
rect 77444 53564 77450 53576
rect 77573 53567 77631 53573
rect 77573 53564 77585 53567
rect 77444 53536 77585 53564
rect 77444 53524 77450 53536
rect 77573 53533 77585 53536
rect 77619 53533 77631 53567
rect 77573 53527 77631 53533
rect 1486 53496 1492 53508
rect 1447 53468 1492 53496
rect 1486 53456 1492 53468
rect 1544 53496 1550 53508
rect 2133 53499 2191 53505
rect 2133 53496 2145 53499
rect 1544 53468 2145 53496
rect 1544 53456 1550 53468
rect 2133 53465 2145 53468
rect 2179 53465 2191 53499
rect 2133 53459 2191 53465
rect 53282 53456 53288 53508
rect 53340 53496 53346 53508
rect 53837 53499 53895 53505
rect 53837 53496 53849 53499
rect 53340 53468 53849 53496
rect 53340 53456 53346 53468
rect 53837 53465 53849 53468
rect 53883 53496 53895 53499
rect 77662 53496 77668 53508
rect 53883 53468 77668 53496
rect 53883 53465 53895 53468
rect 53837 53459 53895 53465
rect 77662 53456 77668 53468
rect 77720 53456 77726 53508
rect 1581 53431 1639 53437
rect 1581 53397 1593 53431
rect 1627 53428 1639 53431
rect 2682 53428 2688 53440
rect 1627 53400 2688 53428
rect 1627 53397 1639 53400
rect 1581 53391 1639 53397
rect 2682 53388 2688 53400
rect 2740 53388 2746 53440
rect 54110 53388 54116 53440
rect 54168 53428 54174 53440
rect 54297 53431 54355 53437
rect 54297 53428 54309 53431
rect 54168 53400 54309 53428
rect 54168 53388 54174 53400
rect 54297 53397 54309 53400
rect 54343 53397 54355 53431
rect 54297 53391 54355 53397
rect 1104 53338 78844 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 78844 53338
rect 1104 53264 78844 53286
rect 1670 53116 1676 53168
rect 1728 53156 1734 53168
rect 53282 53156 53288 53168
rect 1728 53128 53144 53156
rect 53243 53128 53288 53156
rect 1728 53116 1734 53128
rect 1486 53088 1492 53100
rect 1447 53060 1492 53088
rect 1486 53048 1492 53060
rect 1544 53088 1550 53100
rect 2133 53091 2191 53097
rect 2133 53088 2145 53091
rect 1544 53060 2145 53088
rect 1544 53048 1550 53060
rect 2133 53057 2145 53060
rect 2179 53057 2191 53091
rect 52822 53088 52828 53100
rect 2133 53051 2191 53057
rect 45526 53060 52828 53088
rect 1673 52955 1731 52961
rect 1673 52921 1685 52955
rect 1719 52952 1731 52955
rect 1719 52924 6914 52952
rect 1719 52921 1731 52924
rect 1673 52915 1731 52921
rect 6886 52884 6914 52924
rect 45526 52884 45554 53060
rect 52822 53048 52828 53060
rect 52880 53088 52886 53100
rect 53009 53091 53067 53097
rect 53009 53088 53021 53091
rect 52880 53060 53021 53088
rect 52880 53048 52886 53060
rect 53009 53057 53021 53060
rect 53055 53057 53067 53091
rect 53009 53051 53067 53057
rect 53116 53020 53144 53128
rect 53282 53116 53288 53128
rect 53340 53116 53346 53168
rect 53852 53128 54524 53156
rect 53852 53100 53880 53128
rect 53190 53048 53196 53100
rect 53248 53088 53254 53100
rect 53429 53091 53487 53097
rect 53248 53060 53293 53088
rect 53248 53048 53254 53060
rect 53429 53057 53441 53091
rect 53475 53088 53487 53091
rect 53834 53088 53840 53100
rect 53475 53060 53840 53088
rect 53475 53057 53487 53060
rect 53429 53051 53487 53057
rect 53834 53048 53840 53060
rect 53892 53048 53898 53100
rect 54110 53088 54116 53100
rect 54023 53060 54116 53088
rect 54110 53048 54116 53060
rect 54168 53048 54174 53100
rect 54496 53097 54524 53128
rect 54297 53091 54355 53097
rect 54297 53057 54309 53091
rect 54343 53057 54355 53091
rect 54297 53051 54355 53057
rect 54389 53091 54447 53097
rect 54389 53057 54401 53091
rect 54435 53057 54447 53091
rect 54389 53051 54447 53057
rect 54486 53091 54544 53097
rect 54486 53057 54498 53091
rect 54532 53057 54544 53091
rect 77662 53088 77668 53100
rect 77623 53060 77668 53088
rect 54486 53051 54544 53057
rect 54128 53020 54156 53048
rect 53116 52992 54156 53020
rect 53190 52912 53196 52964
rect 53248 52952 53254 52964
rect 54312 52952 54340 53051
rect 54404 53020 54432 53051
rect 77662 53048 77668 53060
rect 77720 53048 77726 53100
rect 54404 52992 55352 53020
rect 53248 52924 54340 52952
rect 53248 52912 53254 52924
rect 6886 52856 45554 52884
rect 53282 52844 53288 52896
rect 53340 52884 53346 52896
rect 53561 52887 53619 52893
rect 53561 52884 53573 52887
rect 53340 52856 53573 52884
rect 53340 52844 53346 52856
rect 53561 52853 53573 52856
rect 53607 52853 53619 52887
rect 53561 52847 53619 52853
rect 54665 52887 54723 52893
rect 54665 52853 54677 52887
rect 54711 52884 54723 52887
rect 55214 52884 55220 52896
rect 54711 52856 55220 52884
rect 54711 52853 54723 52856
rect 54665 52847 54723 52853
rect 55214 52844 55220 52856
rect 55272 52844 55278 52896
rect 55324 52893 55352 52992
rect 77570 52980 77576 53032
rect 77628 53020 77634 53032
rect 77941 53023 77999 53029
rect 77941 53020 77953 53023
rect 77628 52992 77953 53020
rect 77628 52980 77634 52992
rect 77941 52989 77953 52992
rect 77987 52989 77999 53023
rect 77941 52983 77999 52989
rect 55309 52887 55367 52893
rect 55309 52853 55321 52887
rect 55355 52884 55367 52887
rect 77478 52884 77484 52896
rect 55355 52856 77484 52884
rect 55355 52853 55367 52856
rect 55309 52847 55367 52853
rect 77478 52844 77484 52856
rect 77536 52844 77542 52896
rect 1104 52794 78844 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 78844 52794
rect 1104 52720 78844 52742
rect 52822 52680 52828 52692
rect 52783 52652 52828 52680
rect 52822 52640 52828 52652
rect 52880 52640 52886 52692
rect 77570 52612 77576 52624
rect 77531 52584 77576 52612
rect 77570 52572 77576 52584
rect 77628 52572 77634 52624
rect 51810 52504 51816 52556
rect 51868 52544 51874 52556
rect 52365 52547 52423 52553
rect 52365 52544 52377 52547
rect 51868 52516 52377 52544
rect 51868 52504 51874 52516
rect 52365 52513 52377 52516
rect 52411 52544 52423 52547
rect 77386 52544 77392 52556
rect 52411 52516 77392 52544
rect 52411 52513 52423 52516
rect 52365 52507 52423 52513
rect 77386 52504 77392 52516
rect 77444 52504 77450 52556
rect 53374 52476 53380 52488
rect 53335 52448 53380 52476
rect 53374 52436 53380 52448
rect 53432 52436 53438 52488
rect 53653 52479 53711 52485
rect 53653 52445 53665 52479
rect 53699 52476 53711 52479
rect 53834 52476 53840 52488
rect 53699 52448 53840 52476
rect 53699 52445 53711 52448
rect 53653 52439 53711 52445
rect 52178 52368 52184 52420
rect 52236 52408 52242 52420
rect 53668 52408 53696 52439
rect 53834 52436 53840 52448
rect 53892 52436 53898 52488
rect 52236 52380 53696 52408
rect 52236 52368 52242 52380
rect 1486 52340 1492 52352
rect 1447 52312 1492 52340
rect 1486 52300 1492 52312
rect 1544 52300 1550 52352
rect 54757 52343 54815 52349
rect 54757 52309 54769 52343
rect 54803 52340 54815 52343
rect 55030 52340 55036 52352
rect 54803 52312 55036 52340
rect 54803 52309 54815 52312
rect 54757 52303 54815 52309
rect 55030 52300 55036 52312
rect 55088 52300 55094 52352
rect 77938 52300 77944 52352
rect 77996 52340 78002 52352
rect 78033 52343 78091 52349
rect 78033 52340 78045 52343
rect 77996 52312 78045 52340
rect 77996 52300 78002 52312
rect 78033 52309 78045 52312
rect 78079 52309 78091 52343
rect 78033 52303 78091 52309
rect 1104 52250 78844 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 78844 52250
rect 1104 52176 78844 52198
rect 51810 52068 51816 52080
rect 51771 52040 51816 52068
rect 51810 52028 51816 52040
rect 51868 52028 51874 52080
rect 54849 52071 54907 52077
rect 54849 52068 54861 52071
rect 53392 52040 54861 52068
rect 1486 52000 1492 52012
rect 1447 51972 1492 52000
rect 1486 51960 1492 51972
rect 1544 51960 1550 52012
rect 51537 52003 51595 52009
rect 51537 51969 51549 52003
rect 51583 51969 51595 52003
rect 51718 52000 51724 52012
rect 51679 51972 51724 52000
rect 51537 51963 51595 51969
rect 2682 51824 2688 51876
rect 2740 51864 2746 51876
rect 51077 51867 51135 51873
rect 51077 51864 51089 51867
rect 2740 51836 51089 51864
rect 2740 51824 2746 51836
rect 51077 51833 51089 51836
rect 51123 51864 51135 51867
rect 51552 51864 51580 51963
rect 51718 51960 51724 51972
rect 51776 51960 51782 52012
rect 51957 52003 52015 52009
rect 51957 51969 51969 52003
rect 52003 52000 52015 52003
rect 52178 52000 52184 52012
rect 52003 51972 52184 52000
rect 52003 51969 52015 51972
rect 51957 51963 52015 51969
rect 52178 51960 52184 51972
rect 52236 51960 52242 52012
rect 53190 52000 53196 52012
rect 53024 51972 53196 52000
rect 51736 51932 51764 51960
rect 53024 51932 53052 51972
rect 53190 51960 53196 51972
rect 53248 52000 53254 52012
rect 53392 52009 53420 52040
rect 54849 52037 54861 52040
rect 54895 52037 54907 52071
rect 54849 52031 54907 52037
rect 53377 52003 53435 52009
rect 53377 52000 53389 52003
rect 53248 51972 53389 52000
rect 53248 51960 53254 51972
rect 53377 51969 53389 51972
rect 53423 51969 53435 52003
rect 53377 51963 53435 51969
rect 53834 51960 53840 52012
rect 53892 52000 53898 52012
rect 54613 52003 54671 52009
rect 54613 52000 54625 52003
rect 53892 51972 54625 52000
rect 53892 51960 53898 51972
rect 54613 51969 54625 51972
rect 54659 51969 54671 52003
rect 54613 51963 54671 51969
rect 54757 52003 54815 52009
rect 54757 51969 54769 52003
rect 54803 51969 54815 52003
rect 55030 52000 55036 52012
rect 54991 51972 55036 52000
rect 54757 51963 54815 51969
rect 51736 51904 53052 51932
rect 53098 51892 53104 51944
rect 53156 51932 53162 51944
rect 54772 51932 54800 51963
rect 55030 51960 55036 51972
rect 55088 51960 55094 52012
rect 77665 51935 77723 51941
rect 77665 51932 77677 51935
rect 53156 51904 53201 51932
rect 54772 51904 55628 51932
rect 53156 51892 53162 51904
rect 51123 51836 51580 51864
rect 51123 51833 51135 51836
rect 51077 51827 51135 51833
rect 1578 51796 1584 51808
rect 1539 51768 1584 51796
rect 1578 51756 1584 51768
rect 1636 51756 1642 51808
rect 52086 51796 52092 51808
rect 52047 51768 52092 51796
rect 52086 51756 52092 51768
rect 52144 51756 52150 51808
rect 53834 51756 53840 51808
rect 53892 51796 53898 51808
rect 55600 51805 55628 51904
rect 60706 51904 77677 51932
rect 54481 51799 54539 51805
rect 54481 51796 54493 51799
rect 53892 51768 54493 51796
rect 53892 51756 53898 51768
rect 54481 51765 54493 51768
rect 54527 51765 54539 51799
rect 54481 51759 54539 51765
rect 55585 51799 55643 51805
rect 55585 51765 55597 51799
rect 55631 51796 55643 51799
rect 60706 51796 60734 51904
rect 77665 51901 77677 51904
rect 77711 51901 77723 51935
rect 77938 51932 77944 51944
rect 77899 51904 77944 51932
rect 77665 51895 77723 51901
rect 77938 51892 77944 51904
rect 77996 51892 78002 51944
rect 55631 51768 60734 51796
rect 55631 51765 55643 51768
rect 55585 51759 55643 51765
rect 1104 51706 78844 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 78844 51706
rect 1104 51632 78844 51654
rect 1578 51552 1584 51604
rect 1636 51592 1642 51604
rect 55030 51592 55036 51604
rect 1636 51564 55036 51592
rect 1636 51552 1642 51564
rect 55030 51552 55036 51564
rect 55088 51552 55094 51604
rect 52362 51524 52368 51536
rect 52323 51496 52368 51524
rect 52362 51484 52368 51496
rect 52420 51484 52426 51536
rect 51718 51416 51724 51468
rect 51776 51456 51782 51468
rect 52917 51459 52975 51465
rect 51776 51428 52040 51456
rect 51776 51416 51782 51428
rect 52012 51397 52040 51428
rect 52917 51425 52929 51459
rect 52963 51456 52975 51459
rect 53098 51456 53104 51468
rect 52963 51428 53104 51456
rect 52963 51425 52975 51428
rect 52917 51419 52975 51425
rect 53098 51416 53104 51428
rect 53156 51416 53162 51468
rect 51353 51391 51411 51397
rect 51353 51388 51365 51391
rect 51046 51360 51365 51388
rect 1486 51320 1492 51332
rect 1447 51292 1492 51320
rect 1486 51280 1492 51292
rect 1544 51280 1550 51332
rect 1673 51323 1731 51329
rect 1673 51289 1685 51323
rect 1719 51320 1731 51323
rect 1719 51292 6914 51320
rect 1719 51289 1731 51292
rect 1673 51283 1731 51289
rect 1504 51252 1532 51280
rect 2133 51255 2191 51261
rect 2133 51252 2145 51255
rect 1504 51224 2145 51252
rect 2133 51221 2145 51224
rect 2179 51221 2191 51255
rect 6886 51252 6914 51292
rect 51046 51252 51074 51360
rect 51353 51357 51365 51360
rect 51399 51388 51411 51391
rect 51813 51391 51871 51397
rect 51813 51388 51825 51391
rect 51399 51360 51825 51388
rect 51399 51357 51411 51360
rect 51353 51351 51411 51357
rect 51813 51357 51825 51360
rect 51859 51357 51871 51391
rect 51813 51351 51871 51357
rect 51997 51391 52055 51397
rect 51997 51357 52009 51391
rect 52043 51357 52055 51391
rect 52178 51388 52184 51400
rect 52236 51397 52242 51400
rect 52144 51360 52184 51388
rect 51997 51351 52055 51357
rect 52178 51348 52184 51360
rect 52236 51351 52244 51397
rect 52236 51348 52242 51351
rect 53006 51348 53012 51400
rect 53064 51388 53070 51400
rect 53193 51391 53251 51397
rect 53193 51388 53205 51391
rect 53064 51360 53205 51388
rect 53064 51348 53070 51360
rect 53193 51357 53205 51360
rect 53239 51357 53251 51391
rect 53193 51351 53251 51357
rect 76837 51391 76895 51397
rect 76837 51357 76849 51391
rect 76883 51388 76895 51391
rect 77294 51388 77300 51400
rect 76883 51360 77300 51388
rect 76883 51357 76895 51360
rect 76837 51351 76895 51357
rect 77294 51348 77300 51360
rect 77352 51348 77358 51400
rect 77573 51391 77631 51397
rect 77573 51357 77585 51391
rect 77619 51357 77631 51391
rect 77573 51351 77631 51357
rect 52089 51323 52147 51329
rect 52089 51289 52101 51323
rect 52135 51320 52147 51323
rect 54297 51323 54355 51329
rect 54297 51320 54309 51323
rect 52135 51292 54309 51320
rect 52135 51289 52147 51292
rect 52089 51283 52147 51289
rect 54297 51289 54309 51292
rect 54343 51320 54355 51323
rect 77588 51320 77616 51351
rect 54343 51292 77616 51320
rect 54343 51289 54355 51292
rect 54297 51283 54355 51289
rect 6886 51224 51074 51252
rect 2133 51215 2191 51221
rect 1104 51162 78844 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 78844 51162
rect 1104 51088 78844 51110
rect 1486 50912 1492 50924
rect 1447 50884 1492 50912
rect 1486 50872 1492 50884
rect 1544 50912 1550 50924
rect 2133 50915 2191 50921
rect 2133 50912 2145 50915
rect 1544 50884 2145 50912
rect 1544 50872 1550 50884
rect 2133 50881 2145 50884
rect 2179 50881 2191 50915
rect 2133 50875 2191 50881
rect 53193 50915 53251 50921
rect 53193 50881 53205 50915
rect 53239 50912 53251 50915
rect 53374 50912 53380 50924
rect 53239 50884 53380 50912
rect 53239 50881 53251 50884
rect 53193 50875 53251 50881
rect 53374 50872 53380 50884
rect 53432 50872 53438 50924
rect 53466 50844 53472 50856
rect 53427 50816 53472 50844
rect 53466 50804 53472 50816
rect 53524 50804 53530 50856
rect 76653 50847 76711 50853
rect 76653 50813 76665 50847
rect 76699 50844 76711 50847
rect 77110 50844 77116 50856
rect 76699 50816 77116 50844
rect 76699 50813 76711 50816
rect 76653 50807 76711 50813
rect 77110 50804 77116 50816
rect 77168 50804 77174 50856
rect 77202 50804 77208 50856
rect 77260 50844 77266 50856
rect 77389 50847 77447 50853
rect 77389 50844 77401 50847
rect 77260 50816 77401 50844
rect 77260 50804 77266 50816
rect 77389 50813 77401 50816
rect 77435 50813 77447 50847
rect 77389 50807 77447 50813
rect 1673 50779 1731 50785
rect 1673 50745 1685 50779
rect 1719 50776 1731 50779
rect 1719 50748 6914 50776
rect 1719 50745 1731 50748
rect 1673 50739 1731 50745
rect 6886 50708 6914 50748
rect 50246 50708 50252 50720
rect 6886 50680 50252 50708
rect 50246 50668 50252 50680
rect 50304 50668 50310 50720
rect 1104 50618 78844 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 78844 50618
rect 1104 50544 78844 50566
rect 50246 50504 50252 50516
rect 50207 50476 50252 50504
rect 50246 50464 50252 50476
rect 50304 50464 50310 50516
rect 51997 50507 52055 50513
rect 51997 50473 52009 50507
rect 52043 50504 52055 50507
rect 52043 50476 52408 50504
rect 52043 50473 52055 50476
rect 51997 50467 52055 50473
rect 2498 50328 2504 50380
rect 2556 50368 2562 50380
rect 2556 50340 45554 50368
rect 2556 50328 2562 50340
rect 1486 50232 1492 50244
rect 1447 50204 1492 50232
rect 1486 50192 1492 50204
rect 1544 50192 1550 50244
rect 1673 50235 1731 50241
rect 1673 50201 1685 50235
rect 1719 50232 1731 50235
rect 45526 50232 45554 50340
rect 50264 50300 50292 50464
rect 51353 50439 51411 50445
rect 51353 50405 51365 50439
rect 51399 50436 51411 50439
rect 51810 50436 51816 50448
rect 51399 50408 51816 50436
rect 51399 50405 51411 50408
rect 51353 50399 51411 50405
rect 51810 50396 51816 50408
rect 51868 50396 51874 50448
rect 52012 50368 52040 50467
rect 52380 50436 52408 50476
rect 53374 50436 53380 50448
rect 52380 50408 53236 50436
rect 53335 50408 53380 50436
rect 53208 50368 53236 50408
rect 53374 50396 53380 50408
rect 53432 50396 53438 50448
rect 51092 50340 52040 50368
rect 52564 50340 52960 50368
rect 53208 50340 60734 50368
rect 51092 50309 51120 50340
rect 50801 50303 50859 50309
rect 50801 50300 50813 50303
rect 50264 50272 50813 50300
rect 50801 50269 50813 50272
rect 50847 50269 50859 50303
rect 50801 50263 50859 50269
rect 51077 50303 51135 50309
rect 51077 50269 51089 50303
rect 51123 50269 51135 50303
rect 51077 50263 51135 50269
rect 51166 50260 51172 50312
rect 51224 50309 51230 50312
rect 51224 50303 51279 50309
rect 51224 50269 51233 50303
rect 51267 50300 51279 50303
rect 52564 50300 52592 50340
rect 51267 50272 52592 50300
rect 51267 50269 51279 50272
rect 51224 50263 51279 50269
rect 51224 50260 51230 50263
rect 52730 50260 52736 50312
rect 52788 50300 52794 50312
rect 52825 50303 52883 50309
rect 52825 50300 52837 50303
rect 52788 50272 52837 50300
rect 52788 50260 52794 50272
rect 52825 50269 52837 50272
rect 52871 50269 52883 50303
rect 52932 50300 52960 50340
rect 53245 50303 53303 50309
rect 53245 50300 53257 50303
rect 52932 50272 53257 50300
rect 52825 50263 52883 50269
rect 53245 50269 53257 50272
rect 53291 50300 53303 50303
rect 53466 50300 53472 50312
rect 53291 50272 53472 50300
rect 53291 50269 53303 50272
rect 53245 50263 53303 50269
rect 53466 50260 53472 50272
rect 53524 50260 53530 50312
rect 1719 50204 6914 50232
rect 45526 50204 50936 50232
rect 1719 50201 1731 50204
rect 1673 50195 1731 50201
rect 1504 50164 1532 50192
rect 2133 50167 2191 50173
rect 2133 50164 2145 50167
rect 1504 50136 2145 50164
rect 2133 50133 2145 50136
rect 2179 50133 2191 50167
rect 6886 50164 6914 50204
rect 49786 50164 49792 50176
rect 6886 50136 49792 50164
rect 2133 50127 2191 50133
rect 49786 50124 49792 50136
rect 49844 50124 49850 50176
rect 50908 50164 50936 50204
rect 50982 50192 50988 50244
rect 51040 50232 51046 50244
rect 53006 50232 53012 50244
rect 51040 50204 53012 50232
rect 51040 50192 51046 50204
rect 53006 50192 53012 50204
rect 53064 50192 53070 50244
rect 53101 50235 53159 50241
rect 53101 50201 53113 50235
rect 53147 50201 53159 50235
rect 60706 50232 60734 50340
rect 77297 50303 77355 50309
rect 77297 50269 77309 50303
rect 77343 50300 77355 50303
rect 77386 50300 77392 50312
rect 77343 50272 77392 50300
rect 77343 50269 77355 50272
rect 77297 50263 77355 50269
rect 77386 50260 77392 50272
rect 77444 50260 77450 50312
rect 77570 50300 77576 50312
rect 77531 50272 77576 50300
rect 77570 50260 77576 50272
rect 77628 50260 77634 50312
rect 77202 50232 77208 50244
rect 60706 50204 77208 50232
rect 53101 50195 53159 50201
rect 52730 50164 52736 50176
rect 50908 50136 52736 50164
rect 52730 50124 52736 50136
rect 52788 50124 52794 50176
rect 53116 50164 53144 50195
rect 77202 50192 77208 50204
rect 77260 50192 77266 50244
rect 54021 50167 54079 50173
rect 54021 50164 54033 50167
rect 53116 50136 54033 50164
rect 54021 50133 54033 50136
rect 54067 50164 54079 50167
rect 77754 50164 77760 50176
rect 54067 50136 77760 50164
rect 54067 50133 54079 50136
rect 54021 50127 54079 50133
rect 77754 50124 77760 50136
rect 77812 50124 77818 50176
rect 1104 50074 78844 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 78844 50074
rect 1104 50000 78844 50022
rect 49786 49960 49792 49972
rect 49747 49932 49792 49960
rect 49786 49920 49792 49932
rect 49844 49920 49850 49972
rect 50338 49920 50344 49972
rect 50396 49960 50402 49972
rect 50982 49960 50988 49972
rect 50396 49932 50988 49960
rect 50396 49920 50402 49932
rect 49804 49824 49832 49920
rect 50540 49901 50568 49932
rect 50982 49920 50988 49932
rect 51040 49920 51046 49972
rect 52730 49960 52736 49972
rect 52691 49932 52736 49960
rect 52730 49920 52736 49932
rect 52788 49920 52794 49972
rect 50525 49895 50583 49901
rect 50525 49861 50537 49895
rect 50571 49861 50583 49895
rect 50525 49855 50583 49861
rect 50617 49895 50675 49901
rect 50617 49861 50629 49895
rect 50663 49892 50675 49895
rect 77386 49892 77392 49904
rect 50663 49864 51580 49892
rect 77347 49864 77392 49892
rect 50663 49861 50675 49864
rect 50617 49855 50675 49861
rect 50341 49827 50399 49833
rect 50341 49824 50353 49827
rect 49804 49796 50353 49824
rect 50341 49793 50353 49796
rect 50387 49793 50399 49827
rect 50706 49824 50712 49836
rect 50671 49796 50712 49824
rect 50341 49787 50399 49793
rect 50706 49784 50712 49796
rect 50764 49833 50770 49836
rect 50764 49827 50819 49833
rect 50764 49793 50773 49827
rect 50807 49824 50819 49827
rect 51166 49824 51172 49836
rect 50807 49796 51172 49824
rect 50807 49793 50819 49796
rect 50764 49787 50819 49793
rect 50764 49784 50770 49787
rect 51166 49784 51172 49796
rect 51224 49784 51230 49836
rect 51258 49756 51264 49768
rect 50908 49728 51264 49756
rect 50908 49697 50936 49728
rect 51258 49716 51264 49728
rect 51316 49716 51322 49768
rect 51552 49765 51580 49864
rect 77386 49852 77392 49864
rect 77444 49852 77450 49904
rect 51537 49759 51595 49765
rect 51537 49725 51549 49759
rect 51583 49756 51595 49759
rect 77570 49756 77576 49768
rect 51583 49728 77576 49756
rect 51583 49725 51595 49728
rect 51537 49719 51595 49725
rect 77570 49716 77576 49728
rect 77628 49716 77634 49768
rect 50893 49691 50951 49697
rect 50893 49657 50905 49691
rect 50939 49657 50951 49691
rect 50893 49651 50951 49657
rect 1486 49620 1492 49632
rect 1447 49592 1492 49620
rect 1486 49580 1492 49592
rect 1544 49580 1550 49632
rect 77941 49623 77999 49629
rect 77941 49589 77953 49623
rect 77987 49620 77999 49623
rect 78122 49620 78128 49632
rect 77987 49592 78128 49620
rect 77987 49589 77999 49592
rect 77941 49583 77999 49589
rect 78122 49580 78128 49592
rect 78180 49580 78186 49632
rect 1104 49530 78844 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 78844 49530
rect 1104 49456 78844 49478
rect 50614 49308 50620 49360
rect 50672 49348 50678 49360
rect 50709 49351 50767 49357
rect 50709 49348 50721 49351
rect 50672 49320 50721 49348
rect 50672 49308 50678 49320
rect 50709 49317 50721 49320
rect 50755 49317 50767 49351
rect 50709 49311 50767 49317
rect 1486 49212 1492 49224
rect 1447 49184 1492 49212
rect 1486 49172 1492 49184
rect 1544 49172 1550 49224
rect 50157 49215 50215 49221
rect 50157 49212 50169 49215
rect 49528 49184 50169 49212
rect 49528 49085 49556 49184
rect 50157 49181 50169 49184
rect 50203 49181 50215 49215
rect 50338 49212 50344 49224
rect 50299 49184 50344 49212
rect 50157 49175 50215 49181
rect 50338 49172 50344 49184
rect 50396 49172 50402 49224
rect 50577 49215 50635 49221
rect 50577 49181 50589 49215
rect 50623 49212 50635 49215
rect 50706 49212 50712 49224
rect 50623 49184 50712 49212
rect 50623 49181 50635 49184
rect 50577 49175 50635 49181
rect 50706 49172 50712 49184
rect 50764 49172 50770 49224
rect 77849 49215 77907 49221
rect 77849 49212 77861 49215
rect 64846 49184 77861 49212
rect 50433 49147 50491 49153
rect 50433 49113 50445 49147
rect 50479 49113 50491 49147
rect 50433 49107 50491 49113
rect 1581 49079 1639 49085
rect 1581 49045 1593 49079
rect 1627 49076 1639 49079
rect 49513 49079 49571 49085
rect 49513 49076 49525 49079
rect 1627 49048 49525 49076
rect 1627 49045 1639 49048
rect 1581 49039 1639 49045
rect 49513 49045 49525 49048
rect 49559 49045 49571 49079
rect 50448 49076 50476 49107
rect 51353 49079 51411 49085
rect 51353 49076 51365 49079
rect 50448 49048 51365 49076
rect 49513 49039 49571 49045
rect 51353 49045 51365 49048
rect 51399 49076 51411 49079
rect 64846 49076 64874 49184
rect 77849 49181 77861 49184
rect 77895 49181 77907 49215
rect 78122 49212 78128 49224
rect 78083 49184 78128 49212
rect 77849 49175 77907 49181
rect 78122 49172 78128 49184
rect 78180 49172 78186 49224
rect 51399 49048 64874 49076
rect 51399 49045 51411 49048
rect 51353 49039 51411 49045
rect 1104 48986 78844 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 78844 48986
rect 1104 48912 78844 48934
rect 50154 48832 50160 48884
rect 50212 48832 50218 48884
rect 50172 48804 50200 48832
rect 50341 48807 50399 48813
rect 50341 48804 50353 48807
rect 50172 48776 50353 48804
rect 50341 48773 50353 48776
rect 50387 48773 50399 48807
rect 50341 48767 50399 48773
rect 1486 48736 1492 48748
rect 1447 48708 1492 48736
rect 1486 48696 1492 48708
rect 1544 48736 1550 48748
rect 2133 48739 2191 48745
rect 2133 48736 2145 48739
rect 1544 48708 2145 48736
rect 1544 48696 1550 48708
rect 2133 48705 2145 48708
rect 2179 48705 2191 48739
rect 50157 48739 50215 48745
rect 50157 48736 50169 48739
rect 2133 48699 2191 48705
rect 49712 48708 50169 48736
rect 1673 48603 1731 48609
rect 1673 48569 1685 48603
rect 1719 48600 1731 48603
rect 1719 48572 6914 48600
rect 1719 48569 1731 48572
rect 1673 48563 1731 48569
rect 6886 48532 6914 48572
rect 49712 48541 49740 48708
rect 50157 48705 50169 48708
rect 50203 48705 50215 48739
rect 50157 48699 50215 48705
rect 50433 48739 50491 48745
rect 50433 48705 50445 48739
rect 50479 48705 50491 48739
rect 50433 48699 50491 48705
rect 50577 48739 50635 48745
rect 50577 48705 50589 48739
rect 50623 48736 50635 48739
rect 50706 48736 50712 48748
rect 50623 48708 50712 48736
rect 50623 48705 50635 48708
rect 50577 48699 50635 48705
rect 50448 48668 50476 48699
rect 50706 48696 50712 48708
rect 50764 48696 50770 48748
rect 76653 48671 76711 48677
rect 50448 48640 51074 48668
rect 49697 48535 49755 48541
rect 49697 48532 49709 48535
rect 6886 48504 49709 48532
rect 49697 48501 49709 48504
rect 49743 48501 49755 48535
rect 49697 48495 49755 48501
rect 49970 48492 49976 48544
rect 50028 48532 50034 48544
rect 50709 48535 50767 48541
rect 50709 48532 50721 48535
rect 50028 48504 50721 48532
rect 50028 48492 50034 48504
rect 50709 48501 50721 48504
rect 50755 48501 50767 48535
rect 51046 48532 51074 48640
rect 76653 48637 76665 48671
rect 76699 48668 76711 48671
rect 77110 48668 77116 48680
rect 76699 48640 77116 48668
rect 76699 48637 76711 48640
rect 76653 48631 76711 48637
rect 77110 48628 77116 48640
rect 77168 48628 77174 48680
rect 77389 48671 77447 48677
rect 77389 48637 77401 48671
rect 77435 48637 77447 48671
rect 77389 48631 77447 48637
rect 77404 48600 77432 48631
rect 64846 48572 77432 48600
rect 51353 48535 51411 48541
rect 51353 48532 51365 48535
rect 51046 48504 51365 48532
rect 50709 48495 50767 48501
rect 51353 48501 51365 48504
rect 51399 48532 51411 48535
rect 64846 48532 64874 48572
rect 51399 48504 64874 48532
rect 51399 48501 51411 48504
rect 51353 48495 51411 48501
rect 1104 48442 78844 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 78844 48442
rect 1104 48368 78844 48390
rect 1673 48127 1731 48133
rect 1673 48093 1685 48127
rect 1719 48093 1731 48127
rect 77849 48127 77907 48133
rect 77849 48124 77861 48127
rect 1673 48087 1731 48093
rect 77312 48096 77861 48124
rect 1688 48056 1716 48087
rect 2225 48059 2283 48065
rect 2225 48056 2237 48059
rect 1688 48028 2237 48056
rect 2225 48025 2237 48028
rect 2271 48056 2283 48059
rect 47762 48056 47768 48068
rect 2271 48028 47768 48056
rect 2271 48025 2283 48028
rect 2225 48019 2283 48025
rect 47762 48016 47768 48028
rect 47820 48016 47826 48068
rect 1486 47988 1492 48000
rect 1447 47960 1492 47988
rect 1486 47948 1492 47960
rect 1544 47948 1550 48000
rect 48133 47991 48191 47997
rect 48133 47957 48145 47991
rect 48179 47988 48191 47991
rect 48314 47988 48320 48000
rect 48179 47960 48320 47988
rect 48179 47957 48191 47960
rect 48133 47951 48191 47957
rect 48314 47948 48320 47960
rect 48372 47948 48378 48000
rect 77018 47948 77024 48000
rect 77076 47988 77082 48000
rect 77312 47997 77340 48096
rect 77849 48093 77861 48096
rect 77895 48093 77907 48127
rect 77849 48087 77907 48093
rect 77297 47991 77355 47997
rect 77297 47988 77309 47991
rect 77076 47960 77309 47988
rect 77076 47948 77082 47960
rect 77297 47957 77309 47960
rect 77343 47957 77355 47991
rect 78030 47988 78036 48000
rect 77991 47960 78036 47988
rect 77297 47951 77355 47957
rect 78030 47948 78036 47960
rect 78088 47948 78094 48000
rect 1104 47898 78844 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 78844 47898
rect 1104 47824 78844 47846
rect 47762 47784 47768 47796
rect 47723 47756 47768 47784
rect 47762 47744 47768 47756
rect 47820 47744 47826 47796
rect 1673 47651 1731 47657
rect 1673 47617 1685 47651
rect 1719 47648 1731 47651
rect 2225 47651 2283 47657
rect 2225 47648 2237 47651
rect 1719 47620 2237 47648
rect 1719 47617 1731 47620
rect 1673 47611 1731 47617
rect 2225 47617 2237 47620
rect 2271 47648 2283 47651
rect 47118 47648 47124 47660
rect 2271 47620 47124 47648
rect 2271 47617 2283 47620
rect 2225 47611 2283 47617
rect 47118 47608 47124 47620
rect 47176 47608 47182 47660
rect 47857 47651 47915 47657
rect 47857 47617 47869 47651
rect 47903 47648 47915 47651
rect 48314 47648 48320 47660
rect 47903 47620 48320 47648
rect 47903 47617 47915 47620
rect 47857 47611 47915 47617
rect 48314 47608 48320 47620
rect 48372 47648 48378 47660
rect 48869 47651 48927 47657
rect 48869 47648 48881 47651
rect 48372 47620 48881 47648
rect 48372 47608 48378 47620
rect 48869 47617 48881 47620
rect 48915 47648 48927 47651
rect 49234 47648 49240 47660
rect 48915 47620 49240 47648
rect 48915 47617 48927 47620
rect 48869 47611 48927 47617
rect 49234 47608 49240 47620
rect 49292 47608 49298 47660
rect 77665 47651 77723 47657
rect 77665 47648 77677 47651
rect 77128 47620 77677 47648
rect 49053 47515 49111 47521
rect 49053 47481 49065 47515
rect 49099 47512 49111 47515
rect 77018 47512 77024 47524
rect 49099 47484 77024 47512
rect 49099 47481 49111 47484
rect 49053 47475 49111 47481
rect 77018 47472 77024 47484
rect 77076 47472 77082 47524
rect 1486 47444 1492 47456
rect 1447 47416 1492 47444
rect 1486 47404 1492 47416
rect 1544 47404 1550 47456
rect 49234 47404 49240 47456
rect 49292 47444 49298 47456
rect 49513 47447 49571 47453
rect 49513 47444 49525 47447
rect 49292 47416 49525 47444
rect 49292 47404 49298 47416
rect 49513 47413 49525 47416
rect 49559 47413 49571 47447
rect 49513 47407 49571 47413
rect 69658 47404 69664 47456
rect 69716 47444 69722 47456
rect 77128 47453 77156 47620
rect 77665 47617 77677 47620
rect 77711 47617 77723 47651
rect 77665 47611 77723 47617
rect 77113 47447 77171 47453
rect 77113 47444 77125 47447
rect 69716 47416 77125 47444
rect 69716 47404 69722 47416
rect 77113 47413 77125 47416
rect 77159 47413 77171 47447
rect 77846 47444 77852 47456
rect 77807 47416 77852 47444
rect 77113 47407 77171 47413
rect 77846 47404 77852 47416
rect 77904 47404 77910 47456
rect 1104 47354 78844 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 78844 47354
rect 1104 47280 78844 47302
rect 47118 47240 47124 47252
rect 47079 47212 47124 47240
rect 47118 47200 47124 47212
rect 47176 47200 47182 47252
rect 47213 47039 47271 47045
rect 47213 47005 47225 47039
rect 47259 47036 47271 47039
rect 47670 47036 47676 47048
rect 47259 47008 47676 47036
rect 47259 47005 47271 47008
rect 47213 46999 47271 47005
rect 47670 46996 47676 47008
rect 47728 47036 47734 47048
rect 48133 47039 48191 47045
rect 48133 47036 48145 47039
rect 47728 47008 48145 47036
rect 47728 46996 47734 47008
rect 48133 47005 48145 47008
rect 48179 47036 48191 47039
rect 48777 47039 48835 47045
rect 48777 47036 48789 47039
rect 48179 47008 48789 47036
rect 48179 47005 48191 47008
rect 48133 46999 48191 47005
rect 48777 47005 48789 47008
rect 48823 47005 48835 47039
rect 48777 46999 48835 47005
rect 48317 46971 48375 46977
rect 48317 46937 48329 46971
rect 48363 46968 48375 46971
rect 69658 46968 69664 46980
rect 48363 46940 69664 46968
rect 48363 46937 48375 46940
rect 48317 46931 48375 46937
rect 69658 46928 69664 46940
rect 69716 46928 69722 46980
rect 1104 46810 78844 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 78844 46810
rect 1104 46736 78844 46758
rect 47670 46696 47676 46708
rect 47631 46668 47676 46696
rect 47670 46656 47676 46668
rect 47728 46656 47734 46708
rect 1673 46563 1731 46569
rect 1673 46529 1685 46563
rect 1719 46560 1731 46563
rect 2225 46563 2283 46569
rect 2225 46560 2237 46563
rect 1719 46532 2237 46560
rect 1719 46529 1731 46532
rect 1673 46523 1731 46529
rect 2225 46529 2237 46532
rect 2271 46560 2283 46563
rect 46382 46560 46388 46572
rect 2271 46532 46388 46560
rect 2271 46529 2283 46532
rect 2225 46523 2283 46529
rect 46382 46520 46388 46532
rect 46440 46520 46446 46572
rect 77665 46563 77723 46569
rect 77665 46560 77677 46563
rect 77128 46532 77677 46560
rect 1486 46424 1492 46436
rect 1447 46396 1492 46424
rect 1486 46384 1492 46396
rect 1544 46384 1550 46436
rect 46753 46359 46811 46365
rect 46753 46325 46765 46359
rect 46799 46356 46811 46359
rect 46934 46356 46940 46368
rect 46799 46328 46940 46356
rect 46799 46325 46811 46328
rect 46753 46319 46811 46325
rect 46934 46316 46940 46328
rect 46992 46316 46998 46368
rect 69658 46316 69664 46368
rect 69716 46356 69722 46368
rect 77128 46365 77156 46532
rect 77665 46529 77677 46532
rect 77711 46529 77723 46563
rect 77665 46523 77723 46529
rect 77846 46424 77852 46436
rect 77807 46396 77852 46424
rect 77846 46384 77852 46396
rect 77904 46384 77910 46436
rect 77113 46359 77171 46365
rect 77113 46356 77125 46359
rect 69716 46328 77125 46356
rect 69716 46316 69722 46328
rect 77113 46325 77125 46328
rect 77159 46325 77171 46359
rect 77113 46319 77171 46325
rect 1104 46266 78844 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 78844 46266
rect 1104 46192 78844 46214
rect 46382 46152 46388 46164
rect 46343 46124 46388 46152
rect 46382 46112 46388 46124
rect 46440 46112 46446 46164
rect 46842 45976 46848 46028
rect 46900 46016 46906 46028
rect 46900 45988 51074 46016
rect 46900 45976 46906 45988
rect 1673 45951 1731 45957
rect 1673 45917 1685 45951
rect 1719 45948 1731 45951
rect 46477 45951 46535 45957
rect 1719 45920 2268 45948
rect 1719 45917 1731 45920
rect 1673 45911 1731 45917
rect 2240 45824 2268 45920
rect 46477 45917 46489 45951
rect 46523 45948 46535 45951
rect 46934 45948 46940 45960
rect 46523 45920 46940 45948
rect 46523 45917 46535 45920
rect 46477 45911 46535 45917
rect 46934 45908 46940 45920
rect 46992 45948 46998 45960
rect 47397 45951 47455 45957
rect 47397 45948 47409 45951
rect 46992 45920 47409 45948
rect 46992 45908 46998 45920
rect 47397 45917 47409 45920
rect 47443 45948 47455 45951
rect 47762 45948 47768 45960
rect 47443 45920 47768 45948
rect 47443 45917 47455 45920
rect 47397 45911 47455 45917
rect 47762 45908 47768 45920
rect 47820 45948 47826 45960
rect 48041 45951 48099 45957
rect 48041 45948 48053 45951
rect 47820 45920 48053 45948
rect 47820 45908 47826 45920
rect 48041 45917 48053 45920
rect 48087 45917 48099 45951
rect 51046 45948 51074 45988
rect 77297 45951 77355 45957
rect 77297 45948 77309 45951
rect 51046 45920 77309 45948
rect 48041 45911 48099 45917
rect 77297 45917 77309 45920
rect 77343 45948 77355 45951
rect 77849 45951 77907 45957
rect 77849 45948 77861 45951
rect 77343 45920 77861 45948
rect 77343 45917 77355 45920
rect 77297 45911 77355 45917
rect 77849 45917 77861 45920
rect 77895 45917 77907 45951
rect 77849 45911 77907 45917
rect 47581 45883 47639 45889
rect 47581 45849 47593 45883
rect 47627 45880 47639 45883
rect 47627 45852 51074 45880
rect 47627 45849 47639 45852
rect 47581 45843 47639 45849
rect 1486 45812 1492 45824
rect 1447 45784 1492 45812
rect 1486 45772 1492 45784
rect 1544 45772 1550 45824
rect 2222 45812 2228 45824
rect 2183 45784 2228 45812
rect 2222 45772 2228 45784
rect 2280 45772 2286 45824
rect 51046 45812 51074 45852
rect 69658 45812 69664 45824
rect 51046 45784 69664 45812
rect 69658 45772 69664 45784
rect 69716 45772 69722 45824
rect 78030 45812 78036 45824
rect 77991 45784 78036 45812
rect 78030 45772 78036 45784
rect 78088 45772 78094 45824
rect 1104 45722 78844 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 78844 45722
rect 1104 45648 78844 45670
rect 46842 45540 46848 45552
rect 46803 45512 46848 45540
rect 46842 45500 46848 45512
rect 46900 45500 46906 45552
rect 1673 45475 1731 45481
rect 1673 45441 1685 45475
rect 1719 45472 1731 45475
rect 2225 45475 2283 45481
rect 2225 45472 2237 45475
rect 1719 45444 2237 45472
rect 1719 45441 1731 45444
rect 1673 45435 1731 45441
rect 2225 45441 2237 45444
rect 2271 45472 2283 45475
rect 44910 45472 44916 45484
rect 2271 45444 44916 45472
rect 2271 45441 2283 45444
rect 2225 45435 2283 45441
rect 44910 45432 44916 45444
rect 44968 45432 44974 45484
rect 45741 45475 45799 45481
rect 45741 45472 45753 45475
rect 45526 45444 45753 45472
rect 45097 45407 45155 45413
rect 45097 45373 45109 45407
rect 45143 45404 45155 45407
rect 45526 45404 45554 45444
rect 45741 45441 45753 45444
rect 45787 45472 45799 45475
rect 46658 45472 46664 45484
rect 45787 45444 46664 45472
rect 45787 45441 45799 45444
rect 45741 45435 45799 45441
rect 46658 45432 46664 45444
rect 46716 45472 46722 45484
rect 47581 45475 47639 45481
rect 47581 45472 47593 45475
rect 46716 45444 47593 45472
rect 46716 45432 46722 45444
rect 47581 45441 47593 45444
rect 47627 45441 47639 45475
rect 77665 45475 77723 45481
rect 77665 45472 77677 45475
rect 47581 45435 47639 45441
rect 77128 45444 77677 45472
rect 45143 45376 45554 45404
rect 45143 45373 45155 45376
rect 45097 45367 45155 45373
rect 2222 45296 2228 45348
rect 2280 45336 2286 45348
rect 45557 45339 45615 45345
rect 45557 45336 45569 45339
rect 2280 45308 45569 45336
rect 2280 45296 2286 45308
rect 45557 45305 45569 45308
rect 45603 45305 45615 45339
rect 45557 45299 45615 45305
rect 1486 45268 1492 45280
rect 1447 45240 1492 45268
rect 1486 45228 1492 45240
rect 1544 45228 1550 45280
rect 69658 45228 69664 45280
rect 69716 45268 69722 45280
rect 77128 45277 77156 45444
rect 77665 45441 77677 45444
rect 77711 45441 77723 45475
rect 77665 45435 77723 45441
rect 77113 45271 77171 45277
rect 77113 45268 77125 45271
rect 69716 45240 77125 45268
rect 69716 45228 69722 45240
rect 77113 45237 77125 45240
rect 77159 45237 77171 45271
rect 77846 45268 77852 45280
rect 77807 45240 77852 45268
rect 77113 45231 77171 45237
rect 77846 45228 77852 45240
rect 77904 45228 77910 45280
rect 1104 45178 78844 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 78844 45178
rect 1104 45104 78844 45126
rect 44910 45024 44916 45076
rect 44968 45064 44974 45076
rect 45097 45067 45155 45073
rect 45097 45064 45109 45067
rect 44968 45036 45109 45064
rect 44968 45024 44974 45036
rect 45097 45033 45109 45036
rect 45143 45033 45155 45067
rect 45097 45027 45155 45033
rect 1673 44863 1731 44869
rect 1673 44829 1685 44863
rect 1719 44860 1731 44863
rect 2225 44863 2283 44869
rect 2225 44860 2237 44863
rect 1719 44832 2237 44860
rect 1719 44829 1731 44832
rect 1673 44823 1731 44829
rect 2225 44829 2237 44832
rect 2271 44860 2283 44863
rect 44266 44860 44272 44872
rect 2271 44832 44272 44860
rect 2271 44829 2283 44832
rect 2225 44823 2283 44829
rect 44266 44820 44272 44832
rect 44324 44820 44330 44872
rect 77849 44863 77907 44869
rect 77849 44860 77861 44863
rect 77312 44832 77861 44860
rect 45189 44795 45247 44801
rect 45189 44761 45201 44795
rect 45235 44792 45247 44795
rect 45922 44792 45928 44804
rect 45235 44764 45928 44792
rect 45235 44761 45247 44764
rect 45189 44755 45247 44761
rect 45922 44752 45928 44764
rect 45980 44752 45986 44804
rect 46109 44795 46167 44801
rect 46109 44761 46121 44795
rect 46155 44792 46167 44795
rect 46155 44764 51074 44792
rect 46155 44761 46167 44764
rect 46109 44755 46167 44761
rect 1486 44724 1492 44736
rect 1447 44696 1492 44724
rect 1486 44684 1492 44696
rect 1544 44684 1550 44736
rect 45940 44724 45968 44752
rect 46569 44727 46627 44733
rect 46569 44724 46581 44727
rect 45940 44696 46581 44724
rect 46569 44693 46581 44696
rect 46615 44693 46627 44727
rect 51046 44724 51074 44764
rect 77312 44736 77340 44832
rect 77849 44829 77861 44832
rect 77895 44829 77907 44863
rect 77849 44823 77907 44829
rect 69658 44724 69664 44736
rect 51046 44696 69664 44724
rect 46569 44687 46627 44693
rect 69658 44684 69664 44696
rect 69716 44684 69722 44736
rect 77294 44724 77300 44736
rect 77255 44696 77300 44724
rect 77294 44684 77300 44696
rect 77352 44684 77358 44736
rect 78030 44724 78036 44736
rect 77991 44696 78036 44724
rect 78030 44684 78036 44696
rect 78088 44684 78094 44736
rect 1104 44634 78844 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 78844 44634
rect 1104 44560 78844 44582
rect 44266 44520 44272 44532
rect 44227 44492 44272 44520
rect 44266 44480 44272 44492
rect 44324 44480 44330 44532
rect 43717 44387 43775 44393
rect 43717 44353 43729 44387
rect 43763 44384 43775 44387
rect 44361 44387 44419 44393
rect 44361 44384 44373 44387
rect 43763 44356 44373 44384
rect 43763 44353 43775 44356
rect 43717 44347 43775 44353
rect 44361 44353 44373 44356
rect 44407 44384 44419 44387
rect 45186 44384 45192 44396
rect 44407 44356 45192 44384
rect 44407 44353 44419 44356
rect 44361 44347 44419 44353
rect 45186 44344 45192 44356
rect 45244 44384 45250 44396
rect 45833 44387 45891 44393
rect 45833 44384 45845 44387
rect 45244 44356 45845 44384
rect 45244 44344 45250 44356
rect 45833 44353 45845 44356
rect 45879 44353 45891 44387
rect 45833 44347 45891 44353
rect 45373 44251 45431 44257
rect 45373 44217 45385 44251
rect 45419 44248 45431 44251
rect 45419 44220 51074 44248
rect 45419 44217 45431 44220
rect 45373 44211 45431 44217
rect 45922 44140 45928 44192
rect 45980 44180 45986 44192
rect 46385 44183 46443 44189
rect 46385 44180 46397 44183
rect 45980 44152 46397 44180
rect 45980 44140 45986 44152
rect 46385 44149 46397 44152
rect 46431 44149 46443 44183
rect 51046 44180 51074 44220
rect 77294 44180 77300 44192
rect 51046 44152 77300 44180
rect 46385 44143 46443 44149
rect 77294 44140 77300 44152
rect 77352 44140 77358 44192
rect 1104 44090 78844 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 78844 44090
rect 1104 44016 78844 44038
rect 1673 43775 1731 43781
rect 1673 43741 1685 43775
rect 1719 43772 1731 43775
rect 2225 43775 2283 43781
rect 2225 43772 2237 43775
rect 1719 43744 2237 43772
rect 1719 43741 1731 43744
rect 1673 43735 1731 43741
rect 2225 43741 2237 43744
rect 2271 43772 2283 43775
rect 43530 43772 43536 43784
rect 2271 43744 43536 43772
rect 2271 43741 2283 43744
rect 2225 43735 2283 43741
rect 43530 43732 43536 43744
rect 43588 43732 43594 43784
rect 77849 43775 77907 43781
rect 77849 43772 77861 43775
rect 77312 43744 77861 43772
rect 77312 43648 77340 43744
rect 77849 43741 77861 43744
rect 77895 43741 77907 43775
rect 77849 43735 77907 43741
rect 1486 43636 1492 43648
rect 1447 43608 1492 43636
rect 1486 43596 1492 43608
rect 1544 43596 1550 43648
rect 43901 43639 43959 43645
rect 43901 43605 43913 43639
rect 43947 43636 43959 43639
rect 44266 43636 44272 43648
rect 43947 43608 44272 43636
rect 43947 43605 43959 43608
rect 43901 43599 43959 43605
rect 44266 43596 44272 43608
rect 44324 43636 44330 43648
rect 44361 43639 44419 43645
rect 44361 43636 44373 43639
rect 44324 43608 44373 43636
rect 44324 43596 44330 43608
rect 44361 43605 44373 43608
rect 44407 43605 44419 43639
rect 77294 43636 77300 43648
rect 77255 43608 77300 43636
rect 44361 43599 44419 43605
rect 77294 43596 77300 43608
rect 77352 43596 77358 43648
rect 78030 43636 78036 43648
rect 77991 43608 78036 43636
rect 78030 43596 78036 43608
rect 78088 43596 78094 43648
rect 1104 43546 78844 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 78844 43546
rect 1104 43472 78844 43494
rect 43530 43432 43536 43444
rect 43491 43404 43536 43432
rect 43530 43392 43536 43404
rect 43588 43392 43594 43444
rect 1673 43299 1731 43305
rect 1673 43265 1685 43299
rect 1719 43296 1731 43299
rect 43625 43299 43683 43305
rect 1719 43268 2268 43296
rect 1719 43265 1731 43268
rect 1673 43259 1731 43265
rect 1486 43092 1492 43104
rect 1447 43064 1492 43092
rect 1486 43052 1492 43064
rect 1544 43052 1550 43104
rect 2240 43101 2268 43268
rect 43625 43265 43637 43299
rect 43671 43296 43683 43299
rect 44266 43296 44272 43308
rect 43671 43268 44272 43296
rect 43671 43265 43683 43268
rect 43625 43259 43683 43265
rect 44266 43256 44272 43268
rect 44324 43296 44330 43308
rect 44453 43299 44511 43305
rect 44453 43296 44465 43299
rect 44324 43268 44465 43296
rect 44324 43256 44330 43268
rect 44453 43265 44465 43268
rect 44499 43265 44511 43299
rect 44453 43259 44511 43265
rect 77665 43299 77723 43305
rect 77665 43265 77677 43299
rect 77711 43265 77723 43299
rect 77665 43259 77723 43265
rect 44637 43163 44695 43169
rect 44637 43129 44649 43163
rect 44683 43160 44695 43163
rect 77294 43160 77300 43172
rect 44683 43132 77300 43160
rect 44683 43129 44695 43132
rect 44637 43123 44695 43129
rect 77294 43120 77300 43132
rect 77352 43120 77358 43172
rect 2225 43095 2283 43101
rect 2225 43061 2237 43095
rect 2271 43092 2283 43095
rect 2314 43092 2320 43104
rect 2271 43064 2320 43092
rect 2271 43061 2283 43064
rect 2225 43055 2283 43061
rect 2314 43052 2320 43064
rect 2372 43052 2378 43104
rect 76926 43052 76932 43104
rect 76984 43092 76990 43104
rect 77113 43095 77171 43101
rect 77113 43092 77125 43095
rect 76984 43064 77125 43092
rect 76984 43052 76990 43064
rect 77113 43061 77125 43064
rect 77159 43092 77171 43095
rect 77680 43092 77708 43259
rect 77846 43092 77852 43104
rect 77159 43064 77708 43092
rect 77807 43064 77852 43092
rect 77159 43061 77171 43064
rect 77113 43055 77171 43061
rect 77846 43052 77852 43064
rect 77904 43052 77910 43104
rect 1104 43002 78844 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 78844 43002
rect 1104 42928 78844 42950
rect 1673 42687 1731 42693
rect 1673 42653 1685 42687
rect 1719 42653 1731 42687
rect 1673 42647 1731 42653
rect 1688 42616 1716 42647
rect 2314 42644 2320 42696
rect 2372 42684 2378 42696
rect 42705 42687 42763 42693
rect 42705 42684 42717 42687
rect 2372 42656 42717 42684
rect 2372 42644 2378 42656
rect 42705 42653 42717 42656
rect 42751 42653 42763 42687
rect 77849 42687 77907 42693
rect 77849 42684 77861 42687
rect 42705 42647 42763 42653
rect 77312 42656 77861 42684
rect 2225 42619 2283 42625
rect 2225 42616 2237 42619
rect 1688 42588 2237 42616
rect 2225 42585 2237 42588
rect 2271 42616 2283 42619
rect 42518 42616 42524 42628
rect 2271 42588 42524 42616
rect 2271 42585 2283 42588
rect 2225 42579 2283 42585
rect 42518 42576 42524 42588
rect 42576 42576 42582 42628
rect 42889 42619 42947 42625
rect 42889 42585 42901 42619
rect 42935 42616 42947 42619
rect 43717 42619 43775 42625
rect 43717 42616 43729 42619
rect 42935 42588 43729 42616
rect 42935 42585 42947 42588
rect 42889 42579 42947 42585
rect 43717 42585 43729 42588
rect 43763 42585 43775 42619
rect 43717 42579 43775 42585
rect 43901 42619 43959 42625
rect 43901 42585 43913 42619
rect 43947 42616 43959 42619
rect 43947 42588 45554 42616
rect 43947 42585 43959 42588
rect 43901 42579 43959 42585
rect 1486 42548 1492 42560
rect 1447 42520 1492 42548
rect 1486 42508 1492 42520
rect 1544 42508 1550 42560
rect 42245 42551 42303 42557
rect 42245 42517 42257 42551
rect 42291 42548 42303 42551
rect 42904 42548 42932 42579
rect 42291 42520 42932 42548
rect 43732 42548 43760 42579
rect 44174 42548 44180 42560
rect 43732 42520 44180 42548
rect 42291 42517 42303 42520
rect 42245 42511 42303 42517
rect 44174 42508 44180 42520
rect 44232 42548 44238 42560
rect 44361 42551 44419 42557
rect 44361 42548 44373 42551
rect 44232 42520 44373 42548
rect 44232 42508 44238 42520
rect 44361 42517 44373 42520
rect 44407 42517 44419 42551
rect 45526 42548 45554 42588
rect 76926 42548 76932 42560
rect 45526 42520 76932 42548
rect 44361 42511 44419 42517
rect 76926 42508 76932 42520
rect 76984 42508 76990 42560
rect 77018 42508 77024 42560
rect 77076 42548 77082 42560
rect 77312 42557 77340 42656
rect 77849 42653 77861 42656
rect 77895 42653 77907 42687
rect 77849 42647 77907 42653
rect 77297 42551 77355 42557
rect 77297 42548 77309 42551
rect 77076 42520 77309 42548
rect 77076 42508 77082 42520
rect 77297 42517 77309 42520
rect 77343 42517 77355 42551
rect 78030 42548 78036 42560
rect 77991 42520 78036 42548
rect 77297 42511 77355 42517
rect 78030 42508 78036 42520
rect 78088 42508 78094 42560
rect 1104 42458 78844 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 78844 42458
rect 1104 42384 78844 42406
rect 42518 42344 42524 42356
rect 42479 42316 42524 42344
rect 42518 42304 42524 42316
rect 42576 42304 42582 42356
rect 1673 42211 1731 42217
rect 1673 42177 1685 42211
rect 1719 42208 1731 42211
rect 42613 42211 42671 42217
rect 1719 42180 2268 42208
rect 1719 42177 1731 42180
rect 1673 42171 1731 42177
rect 2240 42081 2268 42180
rect 42613 42177 42625 42211
rect 42659 42208 42671 42211
rect 43257 42211 43315 42217
rect 43257 42208 43269 42211
rect 42659 42180 43269 42208
rect 42659 42177 42671 42180
rect 42613 42171 42671 42177
rect 43257 42177 43269 42180
rect 43303 42208 43315 42211
rect 43346 42208 43352 42220
rect 43303 42180 43352 42208
rect 43303 42177 43315 42180
rect 43257 42171 43315 42177
rect 43346 42168 43352 42180
rect 43404 42208 43410 42220
rect 43901 42211 43959 42217
rect 43901 42208 43913 42211
rect 43404 42180 43913 42208
rect 43404 42168 43410 42180
rect 43901 42177 43913 42180
rect 43947 42177 43959 42211
rect 77665 42211 77723 42217
rect 77665 42208 77677 42211
rect 43901 42171 43959 42177
rect 77128 42180 77677 42208
rect 2225 42075 2283 42081
rect 2225 42041 2237 42075
rect 2271 42072 2283 42075
rect 41322 42072 41328 42084
rect 2271 42044 41328 42072
rect 2271 42041 2283 42044
rect 2225 42035 2283 42041
rect 41322 42032 41328 42044
rect 41380 42032 41386 42084
rect 43441 42075 43499 42081
rect 43441 42041 43453 42075
rect 43487 42072 43499 42075
rect 77018 42072 77024 42084
rect 43487 42044 77024 42072
rect 43487 42041 43499 42044
rect 43441 42035 43499 42041
rect 77018 42032 77024 42044
rect 77076 42032 77082 42084
rect 1486 42004 1492 42016
rect 1447 41976 1492 42004
rect 1486 41964 1492 41976
rect 1544 41964 1550 42016
rect 69658 41964 69664 42016
rect 69716 42004 69722 42016
rect 77128 42013 77156 42180
rect 77665 42177 77677 42180
rect 77711 42177 77723 42211
rect 77665 42171 77723 42177
rect 77113 42007 77171 42013
rect 77113 42004 77125 42007
rect 69716 41976 77125 42004
rect 69716 41964 69722 41976
rect 77113 41973 77125 41976
rect 77159 41973 77171 42007
rect 77846 42004 77852 42016
rect 77807 41976 77852 42004
rect 77113 41967 77171 41973
rect 77846 41964 77852 41976
rect 77904 41964 77910 42016
rect 1104 41914 78844 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 78844 41914
rect 1104 41840 78844 41862
rect 41322 41732 41328 41744
rect 41283 41704 41328 41732
rect 41322 41692 41328 41704
rect 41380 41692 41386 41744
rect 41509 41599 41567 41605
rect 41509 41565 41521 41599
rect 41555 41596 41567 41599
rect 42337 41599 42395 41605
rect 42337 41596 42349 41599
rect 41555 41568 42349 41596
rect 41555 41565 41567 41568
rect 41509 41559 41567 41565
rect 42337 41565 42349 41568
rect 42383 41596 42395 41599
rect 42610 41596 42616 41608
rect 42383 41568 42616 41596
rect 42383 41565 42395 41568
rect 42337 41559 42395 41565
rect 42610 41556 42616 41568
rect 42668 41556 42674 41608
rect 42521 41531 42579 41537
rect 42521 41497 42533 41531
rect 42567 41528 42579 41531
rect 42567 41500 45554 41528
rect 42567 41497 42579 41500
rect 42521 41491 42579 41497
rect 43073 41463 43131 41469
rect 43073 41429 43085 41463
rect 43119 41460 43131 41463
rect 43346 41460 43352 41472
rect 43119 41432 43352 41460
rect 43119 41429 43131 41432
rect 43073 41423 43131 41429
rect 43346 41420 43352 41432
rect 43404 41420 43410 41472
rect 45526 41460 45554 41500
rect 69658 41460 69664 41472
rect 45526 41432 69664 41460
rect 69658 41420 69664 41432
rect 69716 41420 69722 41472
rect 1104 41370 78844 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 78844 41370
rect 1104 41296 78844 41318
rect 1673 41123 1731 41129
rect 1673 41089 1685 41123
rect 1719 41120 1731 41123
rect 77665 41123 77723 41129
rect 77665 41120 77677 41123
rect 1719 41092 2268 41120
rect 1719 41089 1731 41092
rect 1673 41083 1731 41089
rect 1486 40984 1492 40996
rect 1447 40956 1492 40984
rect 1486 40944 1492 40956
rect 1544 40944 1550 40996
rect 2240 40993 2268 41092
rect 77128 41092 77677 41120
rect 2225 40987 2283 40993
rect 2225 40953 2237 40987
rect 2271 40984 2283 40987
rect 40678 40984 40684 40996
rect 2271 40956 40684 40984
rect 2271 40953 2283 40956
rect 2225 40947 2283 40953
rect 40678 40944 40684 40956
rect 40736 40944 40742 40996
rect 77128 40928 77156 41092
rect 77665 41089 77677 41092
rect 77711 41089 77723 41123
rect 77665 41083 77723 41089
rect 77846 40984 77852 40996
rect 77807 40956 77852 40984
rect 77846 40944 77852 40956
rect 77904 40944 77910 40996
rect 41049 40919 41107 40925
rect 41049 40885 41061 40919
rect 41095 40916 41107 40919
rect 41414 40916 41420 40928
rect 41095 40888 41420 40916
rect 41095 40885 41107 40888
rect 41049 40879 41107 40885
rect 41414 40876 41420 40888
rect 41472 40876 41478 40928
rect 41785 40919 41843 40925
rect 41785 40885 41797 40919
rect 41831 40916 41843 40919
rect 42610 40916 42616 40928
rect 41831 40888 42616 40916
rect 41831 40885 41843 40888
rect 41785 40879 41843 40885
rect 42610 40876 42616 40888
rect 42668 40876 42674 40928
rect 77110 40916 77116 40928
rect 77071 40888 77116 40916
rect 77110 40876 77116 40888
rect 77168 40876 77174 40928
rect 1104 40826 78844 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 78844 40826
rect 1104 40752 78844 40774
rect 40678 40712 40684 40724
rect 40639 40684 40684 40712
rect 40678 40672 40684 40684
rect 40736 40672 40742 40724
rect 1673 40511 1731 40517
rect 1673 40477 1685 40511
rect 1719 40508 1731 40511
rect 77849 40511 77907 40517
rect 77849 40508 77861 40511
rect 1719 40480 2268 40508
rect 1719 40477 1731 40480
rect 1673 40471 1731 40477
rect 1486 40372 1492 40384
rect 1447 40344 1492 40372
rect 1486 40332 1492 40344
rect 1544 40332 1550 40384
rect 2240 40381 2268 40480
rect 77312 40480 77861 40508
rect 40773 40443 40831 40449
rect 40773 40409 40785 40443
rect 40819 40440 40831 40443
rect 41414 40440 41420 40452
rect 40819 40412 41420 40440
rect 40819 40409 40831 40412
rect 40773 40403 40831 40409
rect 41414 40400 41420 40412
rect 41472 40440 41478 40452
rect 41601 40443 41659 40449
rect 41601 40440 41613 40443
rect 41472 40412 41613 40440
rect 41472 40400 41478 40412
rect 41601 40409 41613 40412
rect 41647 40409 41659 40443
rect 41601 40403 41659 40409
rect 41785 40443 41843 40449
rect 41785 40409 41797 40443
rect 41831 40440 41843 40443
rect 77110 40440 77116 40452
rect 41831 40412 77116 40440
rect 41831 40409 41843 40412
rect 41785 40403 41843 40409
rect 77110 40400 77116 40412
rect 77168 40400 77174 40452
rect 2225 40375 2283 40381
rect 2225 40341 2237 40375
rect 2271 40372 2283 40375
rect 2314 40372 2320 40384
rect 2271 40344 2320 40372
rect 2271 40341 2283 40344
rect 2225 40335 2283 40341
rect 2314 40332 2320 40344
rect 2372 40332 2378 40384
rect 41046 40332 41052 40384
rect 41104 40372 41110 40384
rect 77312 40381 77340 40480
rect 77849 40477 77861 40480
rect 77895 40477 77907 40511
rect 77849 40471 77907 40477
rect 77297 40375 77355 40381
rect 77297 40372 77309 40375
rect 41104 40344 77309 40372
rect 41104 40332 41110 40344
rect 77297 40341 77309 40344
rect 77343 40341 77355 40375
rect 78030 40372 78036 40384
rect 77991 40344 78036 40372
rect 77297 40335 77355 40341
rect 78030 40332 78036 40344
rect 78088 40332 78094 40384
rect 1104 40282 78844 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 78844 40282
rect 1104 40208 78844 40230
rect 1673 40035 1731 40041
rect 1673 40001 1685 40035
rect 1719 40032 1731 40035
rect 39393 40035 39451 40041
rect 1719 40004 2268 40032
rect 1719 40001 1731 40004
rect 1673 39995 1731 40001
rect 2240 39905 2268 40004
rect 39393 40001 39405 40035
rect 39439 40032 39451 40035
rect 40037 40035 40095 40041
rect 40037 40032 40049 40035
rect 39439 40004 40049 40032
rect 39439 40001 39451 40004
rect 39393 39995 39451 40001
rect 40037 40001 40049 40004
rect 40083 40032 40095 40035
rect 40586 40032 40592 40044
rect 40083 40004 40592 40032
rect 40083 40001 40095 40004
rect 40037 39995 40095 40001
rect 40586 39992 40592 40004
rect 40644 40032 40650 40044
rect 40865 40035 40923 40041
rect 40865 40032 40877 40035
rect 40644 40004 40877 40032
rect 40644 39992 40650 40004
rect 40865 40001 40877 40004
rect 40911 40001 40923 40035
rect 41046 40032 41052 40044
rect 41007 40004 41052 40032
rect 40865 39995 40923 40001
rect 41046 39992 41052 40004
rect 41104 39992 41110 40044
rect 77665 40035 77723 40041
rect 77665 40032 77677 40035
rect 77128 40004 77677 40032
rect 2314 39924 2320 39976
rect 2372 39964 2378 39976
rect 39853 39967 39911 39973
rect 39853 39964 39865 39967
rect 2372 39936 39865 39964
rect 2372 39924 2378 39936
rect 39853 39933 39865 39936
rect 39899 39933 39911 39967
rect 39853 39927 39911 39933
rect 2225 39899 2283 39905
rect 2225 39865 2237 39899
rect 2271 39896 2283 39899
rect 39114 39896 39120 39908
rect 2271 39868 39120 39896
rect 2271 39865 2283 39868
rect 2225 39859 2283 39865
rect 39114 39856 39120 39868
rect 39172 39856 39178 39908
rect 1486 39828 1492 39840
rect 1447 39800 1492 39828
rect 1486 39788 1492 39800
rect 1544 39788 1550 39840
rect 41414 39788 41420 39840
rect 41472 39828 41478 39840
rect 41509 39831 41567 39837
rect 41509 39828 41521 39831
rect 41472 39800 41521 39828
rect 41472 39788 41478 39800
rect 41509 39797 41521 39800
rect 41555 39797 41567 39831
rect 41509 39791 41567 39797
rect 69658 39788 69664 39840
rect 69716 39828 69722 39840
rect 77128 39837 77156 40004
rect 77665 40001 77677 40004
rect 77711 40001 77723 40035
rect 77665 39995 77723 40001
rect 77113 39831 77171 39837
rect 77113 39828 77125 39831
rect 69716 39800 77125 39828
rect 69716 39788 69722 39800
rect 77113 39797 77125 39800
rect 77159 39797 77171 39831
rect 77846 39828 77852 39840
rect 77807 39800 77852 39828
rect 77113 39791 77171 39797
rect 77846 39788 77852 39800
rect 77904 39788 77910 39840
rect 1104 39738 78844 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 78844 39738
rect 1104 39664 78844 39686
rect 39114 39624 39120 39636
rect 39075 39596 39120 39624
rect 39114 39584 39120 39596
rect 39172 39584 39178 39636
rect 1673 39423 1731 39429
rect 1673 39389 1685 39423
rect 1719 39389 1731 39423
rect 77849 39423 77907 39429
rect 77849 39420 77861 39423
rect 1673 39383 1731 39389
rect 77312 39392 77861 39420
rect 1688 39352 1716 39383
rect 2225 39355 2283 39361
rect 2225 39352 2237 39355
rect 1688 39324 2237 39352
rect 2225 39321 2237 39324
rect 2271 39352 2283 39355
rect 38378 39352 38384 39364
rect 2271 39324 38384 39352
rect 2271 39321 2283 39324
rect 2225 39315 2283 39321
rect 38378 39312 38384 39324
rect 38436 39312 38442 39364
rect 38565 39355 38623 39361
rect 38565 39321 38577 39355
rect 38611 39352 38623 39355
rect 39209 39355 39267 39361
rect 39209 39352 39221 39355
rect 38611 39324 39221 39352
rect 38611 39321 38623 39324
rect 38565 39315 38623 39321
rect 39209 39321 39221 39324
rect 39255 39352 39267 39355
rect 39850 39352 39856 39364
rect 39255 39324 39856 39352
rect 39255 39321 39267 39324
rect 39209 39315 39267 39321
rect 39850 39312 39856 39324
rect 39908 39352 39914 39364
rect 40129 39355 40187 39361
rect 40129 39352 40141 39355
rect 39908 39324 40141 39352
rect 39908 39312 39914 39324
rect 40129 39321 40141 39324
rect 40175 39321 40187 39355
rect 40129 39315 40187 39321
rect 40313 39355 40371 39361
rect 40313 39321 40325 39355
rect 40359 39352 40371 39355
rect 40359 39324 45554 39352
rect 40359 39321 40371 39324
rect 40313 39315 40371 39321
rect 1486 39284 1492 39296
rect 1447 39256 1492 39284
rect 1486 39244 1492 39256
rect 1544 39244 1550 39296
rect 40586 39244 40592 39296
rect 40644 39284 40650 39296
rect 40773 39287 40831 39293
rect 40773 39284 40785 39287
rect 40644 39256 40785 39284
rect 40644 39244 40650 39256
rect 40773 39253 40785 39256
rect 40819 39253 40831 39287
rect 45526 39284 45554 39324
rect 77312 39296 77340 39392
rect 77849 39389 77861 39392
rect 77895 39389 77907 39423
rect 77849 39383 77907 39389
rect 69658 39284 69664 39296
rect 45526 39256 69664 39284
rect 40773 39247 40831 39253
rect 69658 39244 69664 39256
rect 69716 39244 69722 39296
rect 77294 39284 77300 39296
rect 77255 39256 77300 39284
rect 77294 39244 77300 39256
rect 77352 39244 77358 39296
rect 78030 39284 78036 39296
rect 77991 39256 78036 39284
rect 78030 39244 78036 39256
rect 78088 39244 78094 39296
rect 1104 39194 78844 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 78844 39194
rect 1104 39120 78844 39142
rect 38378 39040 38384 39092
rect 38436 39080 38442 39092
rect 38473 39083 38531 39089
rect 38473 39080 38485 39083
rect 38436 39052 38485 39080
rect 38436 39040 38442 39052
rect 38473 39049 38485 39052
rect 38519 39049 38531 39083
rect 38473 39043 38531 39049
rect 37921 38947 37979 38953
rect 37921 38913 37933 38947
rect 37967 38944 37979 38947
rect 38565 38947 38623 38953
rect 38565 38944 38577 38947
rect 37967 38916 38577 38944
rect 37967 38913 37979 38916
rect 37921 38907 37979 38913
rect 38565 38913 38577 38916
rect 38611 38944 38623 38947
rect 39114 38944 39120 38956
rect 38611 38916 39120 38944
rect 38611 38913 38623 38916
rect 38565 38907 38623 38913
rect 39114 38904 39120 38916
rect 39172 38944 39178 38956
rect 39393 38947 39451 38953
rect 39393 38944 39405 38947
rect 39172 38916 39405 38944
rect 39172 38904 39178 38916
rect 39393 38913 39405 38916
rect 39439 38913 39451 38947
rect 39393 38907 39451 38913
rect 39577 38811 39635 38817
rect 39577 38777 39589 38811
rect 39623 38808 39635 38811
rect 39623 38780 45554 38808
rect 39623 38777 39635 38780
rect 39577 38771 39635 38777
rect 39850 38700 39856 38752
rect 39908 38740 39914 38752
rect 40037 38743 40095 38749
rect 40037 38740 40049 38743
rect 39908 38712 40049 38740
rect 39908 38700 39914 38712
rect 40037 38709 40049 38712
rect 40083 38709 40095 38743
rect 45526 38740 45554 38780
rect 77294 38740 77300 38752
rect 45526 38712 77300 38740
rect 40037 38703 40095 38709
rect 77294 38700 77300 38712
rect 77352 38700 77358 38752
rect 1104 38650 78844 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 78844 38650
rect 1104 38576 78844 38598
rect 1673 38335 1731 38341
rect 1673 38301 1685 38335
rect 1719 38301 1731 38335
rect 77849 38335 77907 38341
rect 77849 38332 77861 38335
rect 1673 38295 1731 38301
rect 77312 38304 77861 38332
rect 1688 38264 1716 38295
rect 2225 38267 2283 38273
rect 2225 38264 2237 38267
rect 1688 38236 2237 38264
rect 2225 38233 2237 38236
rect 2271 38264 2283 38267
rect 37734 38264 37740 38276
rect 2271 38236 37740 38264
rect 2271 38233 2283 38236
rect 2225 38227 2283 38233
rect 37734 38224 37740 38236
rect 37792 38224 37798 38276
rect 1486 38196 1492 38208
rect 1447 38168 1492 38196
rect 1486 38156 1492 38168
rect 1544 38156 1550 38208
rect 38378 38196 38384 38208
rect 38339 38168 38384 38196
rect 38378 38156 38384 38168
rect 38436 38156 38442 38208
rect 39114 38196 39120 38208
rect 39075 38168 39120 38196
rect 39114 38156 39120 38168
rect 39172 38156 39178 38208
rect 77018 38156 77024 38208
rect 77076 38196 77082 38208
rect 77312 38205 77340 38304
rect 77849 38301 77861 38304
rect 77895 38301 77907 38335
rect 77849 38295 77907 38301
rect 77297 38199 77355 38205
rect 77297 38196 77309 38199
rect 77076 38168 77309 38196
rect 77076 38156 77082 38168
rect 77297 38165 77309 38168
rect 77343 38165 77355 38199
rect 78030 38196 78036 38208
rect 77991 38168 78036 38196
rect 77297 38159 77355 38165
rect 78030 38156 78036 38168
rect 78088 38156 78094 38208
rect 1104 38106 78844 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 78844 38106
rect 1104 38032 78844 38054
rect 37734 37992 37740 38004
rect 37695 37964 37740 37992
rect 37734 37952 37740 37964
rect 37792 37952 37798 38004
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37856 1731 37859
rect 37829 37859 37887 37865
rect 1719 37828 2268 37856
rect 1719 37825 1731 37828
rect 1673 37819 1731 37825
rect 2240 37729 2268 37828
rect 37829 37825 37841 37859
rect 37875 37856 37887 37859
rect 38378 37856 38384 37868
rect 37875 37828 38384 37856
rect 37875 37825 37887 37828
rect 37829 37819 37887 37825
rect 38378 37816 38384 37828
rect 38436 37856 38442 37868
rect 38657 37859 38715 37865
rect 38657 37856 38669 37859
rect 38436 37828 38669 37856
rect 38436 37816 38442 37828
rect 38657 37825 38669 37828
rect 38703 37825 38715 37859
rect 77665 37859 77723 37865
rect 77665 37856 77677 37859
rect 38657 37819 38715 37825
rect 77128 37828 77677 37856
rect 2225 37723 2283 37729
rect 2225 37689 2237 37723
rect 2271 37720 2283 37723
rect 36998 37720 37004 37732
rect 2271 37692 37004 37720
rect 2271 37689 2283 37692
rect 2225 37683 2283 37689
rect 36998 37680 37004 37692
rect 37056 37680 37062 37732
rect 38841 37723 38899 37729
rect 38841 37689 38853 37723
rect 38887 37720 38899 37723
rect 77018 37720 77024 37732
rect 38887 37692 77024 37720
rect 38887 37689 38899 37692
rect 38841 37683 38899 37689
rect 77018 37680 77024 37692
rect 77076 37680 77082 37732
rect 1486 37652 1492 37664
rect 1447 37624 1492 37652
rect 1486 37612 1492 37624
rect 1544 37612 1550 37664
rect 69658 37612 69664 37664
rect 69716 37652 69722 37664
rect 77128 37661 77156 37828
rect 77665 37825 77677 37828
rect 77711 37825 77723 37859
rect 77665 37819 77723 37825
rect 77113 37655 77171 37661
rect 77113 37652 77125 37655
rect 69716 37624 77125 37652
rect 69716 37612 69722 37624
rect 77113 37621 77125 37624
rect 77159 37621 77171 37655
rect 77846 37652 77852 37664
rect 77807 37624 77852 37652
rect 77113 37615 77171 37621
rect 77846 37612 77852 37624
rect 77904 37612 77910 37664
rect 1104 37562 78844 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 78844 37562
rect 1104 37488 78844 37510
rect 36998 37448 37004 37460
rect 36959 37420 37004 37448
rect 36998 37408 37004 37420
rect 37056 37408 37062 37460
rect 38378 37340 38384 37392
rect 38436 37380 38442 37392
rect 38565 37383 38623 37389
rect 38565 37380 38577 37383
rect 38436 37352 38577 37380
rect 38436 37340 38442 37352
rect 38565 37349 38577 37352
rect 38611 37349 38623 37383
rect 38565 37343 38623 37349
rect 38105 37315 38163 37321
rect 38105 37281 38117 37315
rect 38151 37312 38163 37315
rect 69658 37312 69664 37324
rect 38151 37284 69664 37312
rect 38151 37281 38163 37284
rect 38105 37275 38163 37281
rect 69658 37272 69664 37284
rect 69716 37272 69722 37324
rect 1673 37247 1731 37253
rect 1673 37213 1685 37247
rect 1719 37213 1731 37247
rect 77849 37247 77907 37253
rect 77849 37244 77861 37247
rect 1673 37207 1731 37213
rect 77312 37216 77861 37244
rect 1688 37176 1716 37207
rect 2225 37179 2283 37185
rect 2225 37176 2237 37179
rect 1688 37148 2237 37176
rect 2225 37145 2237 37148
rect 2271 37176 2283 37179
rect 36262 37176 36268 37188
rect 2271 37148 36268 37176
rect 2271 37145 2283 37148
rect 2225 37139 2283 37145
rect 36262 37136 36268 37148
rect 36320 37136 36326 37188
rect 36449 37179 36507 37185
rect 36449 37145 36461 37179
rect 36495 37176 36507 37179
rect 37093 37179 37151 37185
rect 37093 37176 37105 37179
rect 36495 37148 37105 37176
rect 36495 37145 36507 37148
rect 36449 37139 36507 37145
rect 37093 37145 37105 37148
rect 37139 37176 37151 37179
rect 37642 37176 37648 37188
rect 37139 37148 37648 37176
rect 37139 37145 37151 37148
rect 37093 37139 37151 37145
rect 37642 37136 37648 37148
rect 37700 37176 37706 37188
rect 37921 37179 37979 37185
rect 37921 37176 37933 37179
rect 37700 37148 37933 37176
rect 37700 37136 37706 37148
rect 37921 37145 37933 37148
rect 37967 37176 37979 37179
rect 38010 37176 38016 37188
rect 37967 37148 38016 37176
rect 37967 37145 37979 37148
rect 37921 37139 37979 37145
rect 38010 37136 38016 37148
rect 38068 37136 38074 37188
rect 77312 37120 77340 37216
rect 77849 37213 77861 37216
rect 77895 37213 77907 37247
rect 77849 37207 77907 37213
rect 1486 37108 1492 37120
rect 1447 37080 1492 37108
rect 1486 37068 1492 37080
rect 1544 37068 1550 37120
rect 77294 37108 77300 37120
rect 77255 37080 77300 37108
rect 77294 37068 77300 37080
rect 77352 37068 77358 37120
rect 78030 37108 78036 37120
rect 77991 37080 78036 37108
rect 78030 37068 78036 37080
rect 78088 37068 78094 37120
rect 1104 37018 78844 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 78844 37018
rect 1104 36944 78844 36966
rect 36262 36904 36268 36916
rect 36223 36876 36268 36904
rect 36262 36864 36268 36876
rect 36320 36864 36326 36916
rect 38010 36904 38016 36916
rect 37971 36876 38016 36904
rect 38010 36864 38016 36876
rect 38068 36864 38074 36916
rect 77294 36836 77300 36848
rect 64846 36808 77300 36836
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36768 1731 36771
rect 2225 36771 2283 36777
rect 2225 36768 2237 36771
rect 1719 36740 2237 36768
rect 1719 36737 1731 36740
rect 1673 36731 1731 36737
rect 2225 36737 2237 36740
rect 2271 36768 2283 36771
rect 35618 36768 35624 36780
rect 2271 36740 35624 36768
rect 2271 36737 2283 36740
rect 2225 36731 2283 36737
rect 35618 36728 35624 36740
rect 35676 36728 35682 36780
rect 35713 36771 35771 36777
rect 35713 36737 35725 36771
rect 35759 36768 35771 36771
rect 36357 36771 36415 36777
rect 36357 36768 36369 36771
rect 35759 36740 36369 36768
rect 35759 36737 35771 36740
rect 35713 36731 35771 36737
rect 36357 36737 36369 36740
rect 36403 36768 36415 36771
rect 36630 36768 36636 36780
rect 36403 36740 36636 36768
rect 36403 36737 36415 36740
rect 36357 36731 36415 36737
rect 36630 36728 36636 36740
rect 36688 36768 36694 36780
rect 37182 36768 37188 36780
rect 36688 36740 37188 36768
rect 36688 36728 36694 36740
rect 37182 36728 37188 36740
rect 37240 36768 37246 36780
rect 37369 36771 37427 36777
rect 37369 36768 37381 36771
rect 37240 36740 37381 36768
rect 37240 36728 37246 36740
rect 37369 36737 37381 36740
rect 37415 36737 37427 36771
rect 37369 36731 37427 36737
rect 37553 36635 37611 36641
rect 37553 36601 37565 36635
rect 37599 36632 37611 36635
rect 64846 36632 64874 36808
rect 77294 36796 77300 36808
rect 77352 36796 77358 36848
rect 77665 36771 77723 36777
rect 77665 36768 77677 36771
rect 37599 36604 64874 36632
rect 77128 36740 77677 36768
rect 37599 36601 37611 36604
rect 37553 36595 37611 36601
rect 1486 36564 1492 36576
rect 1447 36536 1492 36564
rect 1486 36524 1492 36536
rect 1544 36524 1550 36576
rect 69658 36524 69664 36576
rect 69716 36564 69722 36576
rect 77128 36573 77156 36740
rect 77665 36737 77677 36740
rect 77711 36737 77723 36771
rect 77665 36731 77723 36737
rect 77113 36567 77171 36573
rect 77113 36564 77125 36567
rect 69716 36536 77125 36564
rect 69716 36524 69722 36536
rect 77113 36533 77125 36536
rect 77159 36533 77171 36567
rect 77846 36564 77852 36576
rect 77807 36536 77852 36564
rect 77113 36527 77171 36533
rect 77846 36524 77852 36536
rect 77904 36524 77910 36576
rect 1104 36474 78844 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 78844 36474
rect 1104 36400 78844 36422
rect 35618 36360 35624 36372
rect 35579 36332 35624 36360
rect 35618 36320 35624 36332
rect 35676 36320 35682 36372
rect 37182 36360 37188 36372
rect 37143 36332 37188 36360
rect 37182 36320 37188 36332
rect 37240 36320 37246 36372
rect 35069 36091 35127 36097
rect 35069 36057 35081 36091
rect 35115 36088 35127 36091
rect 35713 36091 35771 36097
rect 35713 36088 35725 36091
rect 35115 36060 35725 36088
rect 35115 36057 35127 36060
rect 35069 36051 35127 36057
rect 35713 36057 35725 36060
rect 35759 36088 35771 36091
rect 36262 36088 36268 36100
rect 35759 36060 36268 36088
rect 35759 36057 35771 36060
rect 35713 36051 35771 36057
rect 36262 36048 36268 36060
rect 36320 36088 36326 36100
rect 36541 36091 36599 36097
rect 36541 36088 36553 36091
rect 36320 36060 36553 36088
rect 36320 36048 36326 36060
rect 36541 36057 36553 36060
rect 36587 36057 36599 36091
rect 36541 36051 36599 36057
rect 36725 36091 36783 36097
rect 36725 36057 36737 36091
rect 36771 36088 36783 36091
rect 36771 36060 45554 36088
rect 36771 36057 36783 36060
rect 36725 36051 36783 36057
rect 45526 36020 45554 36060
rect 69658 36020 69664 36032
rect 45526 35992 69664 36020
rect 69658 35980 69664 35992
rect 69716 35980 69722 36032
rect 1104 35930 78844 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 78844 35930
rect 1104 35856 78844 35878
rect 1673 35683 1731 35689
rect 1673 35649 1685 35683
rect 1719 35680 1731 35683
rect 77665 35683 77723 35689
rect 77665 35680 77677 35683
rect 1719 35652 2268 35680
rect 1719 35649 1731 35652
rect 1673 35643 1731 35649
rect 1486 35544 1492 35556
rect 1447 35516 1492 35544
rect 1486 35504 1492 35516
rect 1544 35504 1550 35556
rect 2240 35553 2268 35652
rect 77128 35652 77677 35680
rect 2225 35547 2283 35553
rect 2225 35513 2237 35547
rect 2271 35544 2283 35547
rect 34698 35544 34704 35556
rect 2271 35516 34704 35544
rect 2271 35513 2283 35516
rect 2225 35507 2283 35513
rect 34698 35504 34704 35516
rect 34756 35504 34762 35556
rect 35621 35479 35679 35485
rect 35621 35445 35633 35479
rect 35667 35476 35679 35479
rect 35710 35476 35716 35488
rect 35667 35448 35716 35476
rect 35667 35445 35679 35448
rect 35621 35439 35679 35445
rect 35710 35436 35716 35448
rect 35768 35436 35774 35488
rect 36262 35476 36268 35488
rect 36223 35448 36268 35476
rect 36262 35436 36268 35448
rect 36320 35436 36326 35488
rect 68002 35436 68008 35488
rect 68060 35476 68066 35488
rect 77128 35485 77156 35652
rect 77665 35649 77677 35652
rect 77711 35649 77723 35683
rect 77665 35643 77723 35649
rect 77846 35544 77852 35556
rect 77807 35516 77852 35544
rect 77846 35504 77852 35516
rect 77904 35504 77910 35556
rect 77113 35479 77171 35485
rect 77113 35476 77125 35479
rect 68060 35448 77125 35476
rect 68060 35436 68066 35448
rect 77113 35445 77125 35448
rect 77159 35445 77171 35479
rect 77113 35439 77171 35445
rect 1104 35386 78844 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 78844 35386
rect 1104 35312 78844 35334
rect 34698 35232 34704 35284
rect 34756 35272 34762 35284
rect 34885 35275 34943 35281
rect 34885 35272 34897 35275
rect 34756 35244 34897 35272
rect 34756 35232 34762 35244
rect 34885 35241 34897 35244
rect 34931 35241 34943 35275
rect 34885 35235 34943 35241
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35068 1731 35071
rect 2225 35071 2283 35077
rect 2225 35068 2237 35071
rect 1719 35040 2237 35068
rect 1719 35037 1731 35040
rect 1673 35031 1731 35037
rect 2225 35037 2237 35040
rect 2271 35068 2283 35071
rect 34146 35068 34152 35080
rect 2271 35040 34152 35068
rect 2271 35037 2283 35040
rect 2225 35031 2283 35037
rect 34146 35028 34152 35040
rect 34204 35028 34210 35080
rect 77849 35071 77907 35077
rect 77849 35068 77861 35071
rect 77312 35040 77861 35068
rect 34790 34960 34796 35012
rect 34848 35000 34854 35012
rect 34977 35003 35035 35009
rect 34977 35000 34989 35003
rect 34848 34972 34989 35000
rect 34848 34960 34854 34972
rect 34977 34969 34989 34972
rect 35023 35000 35035 35003
rect 35710 35000 35716 35012
rect 35023 34972 35716 35000
rect 35023 34969 35035 34972
rect 34977 34963 35035 34969
rect 35710 34960 35716 34972
rect 35768 35000 35774 35012
rect 35805 35003 35863 35009
rect 35805 35000 35817 35003
rect 35768 34972 35817 35000
rect 35768 34960 35774 34972
rect 35805 34969 35817 34972
rect 35851 34969 35863 35003
rect 35805 34963 35863 34969
rect 77312 34944 77340 35040
rect 77849 35037 77861 35040
rect 77895 35037 77907 35071
rect 77849 35031 77907 35037
rect 1486 34932 1492 34944
rect 1447 34904 1492 34932
rect 1486 34892 1492 34904
rect 1544 34892 1550 34944
rect 35897 34935 35955 34941
rect 35897 34901 35909 34935
rect 35943 34932 35955 34935
rect 68002 34932 68008 34944
rect 35943 34904 68008 34932
rect 35943 34901 35955 34904
rect 35897 34895 35955 34901
rect 68002 34892 68008 34904
rect 68060 34892 68066 34944
rect 77294 34932 77300 34944
rect 77255 34904 77300 34932
rect 77294 34892 77300 34904
rect 77352 34892 77358 34944
rect 78030 34932 78036 34944
rect 77991 34904 78036 34932
rect 78030 34892 78036 34904
rect 78088 34892 78094 34944
rect 1104 34842 78844 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 78844 34842
rect 1104 34768 78844 34790
rect 34146 34728 34152 34740
rect 34107 34700 34152 34728
rect 34146 34688 34152 34700
rect 34204 34688 34210 34740
rect 35710 34728 35716 34740
rect 35671 34700 35716 34728
rect 35710 34688 35716 34700
rect 35768 34688 35774 34740
rect 35253 34663 35311 34669
rect 35253 34629 35265 34663
rect 35299 34660 35311 34663
rect 77294 34660 77300 34672
rect 35299 34632 77300 34660
rect 35299 34629 35311 34632
rect 35253 34623 35311 34629
rect 77294 34620 77300 34632
rect 77352 34620 77358 34672
rect 1673 34595 1731 34601
rect 1673 34561 1685 34595
rect 1719 34561 1731 34595
rect 1673 34555 1731 34561
rect 33597 34595 33655 34601
rect 33597 34561 33609 34595
rect 33643 34592 33655 34595
rect 34241 34595 34299 34601
rect 34241 34592 34253 34595
rect 33643 34564 34253 34592
rect 33643 34561 33655 34564
rect 33597 34555 33655 34561
rect 34241 34561 34253 34564
rect 34287 34592 34299 34595
rect 34698 34592 34704 34604
rect 34287 34564 34704 34592
rect 34287 34561 34299 34564
rect 34241 34555 34299 34561
rect 1688 34524 1716 34555
rect 34698 34552 34704 34564
rect 34756 34592 34762 34604
rect 35069 34595 35127 34601
rect 35069 34592 35081 34595
rect 34756 34564 35081 34592
rect 34756 34552 34762 34564
rect 35069 34561 35081 34564
rect 35115 34561 35127 34595
rect 77665 34595 77723 34601
rect 77665 34592 77677 34595
rect 35069 34555 35127 34561
rect 77128 34564 77677 34592
rect 77128 34536 77156 34564
rect 77665 34561 77677 34564
rect 77711 34561 77723 34595
rect 77665 34555 77723 34561
rect 2225 34527 2283 34533
rect 2225 34524 2237 34527
rect 1688 34496 2237 34524
rect 2225 34493 2237 34496
rect 2271 34524 2283 34527
rect 2314 34524 2320 34536
rect 2271 34496 2320 34524
rect 2271 34493 2283 34496
rect 2225 34487 2283 34493
rect 2314 34484 2320 34496
rect 2372 34484 2378 34536
rect 77110 34524 77116 34536
rect 77071 34496 77116 34524
rect 77110 34484 77116 34496
rect 77168 34484 77174 34536
rect 1486 34388 1492 34400
rect 1447 34360 1492 34388
rect 1486 34348 1492 34360
rect 1544 34348 1550 34400
rect 77846 34388 77852 34400
rect 77807 34360 77852 34388
rect 77846 34348 77852 34360
rect 77904 34348 77910 34400
rect 1104 34298 78844 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 78844 34298
rect 1104 34224 78844 34246
rect 1673 33983 1731 33989
rect 1673 33949 1685 33983
rect 1719 33949 1731 33983
rect 1673 33943 1731 33949
rect 1688 33912 1716 33943
rect 2314 33940 2320 33992
rect 2372 33980 2378 33992
rect 33321 33983 33379 33989
rect 33321 33980 33333 33983
rect 2372 33952 33333 33980
rect 2372 33940 2378 33952
rect 33321 33949 33333 33952
rect 33367 33949 33379 33983
rect 77849 33983 77907 33989
rect 77849 33980 77861 33983
rect 33321 33943 33379 33949
rect 77312 33952 77861 33980
rect 2225 33915 2283 33921
rect 2225 33912 2237 33915
rect 1688 33884 2237 33912
rect 2225 33881 2237 33884
rect 2271 33912 2283 33915
rect 32674 33912 32680 33924
rect 2271 33884 32680 33912
rect 2271 33881 2283 33884
rect 2225 33875 2283 33881
rect 32674 33872 32680 33884
rect 32732 33872 32738 33924
rect 33505 33915 33563 33921
rect 33505 33881 33517 33915
rect 33551 33881 33563 33915
rect 34793 33915 34851 33921
rect 34793 33912 34805 33915
rect 33505 33875 33563 33881
rect 34072 33884 34805 33912
rect 1486 33844 1492 33856
rect 1447 33816 1492 33844
rect 1486 33804 1492 33816
rect 1544 33804 1550 33856
rect 32861 33847 32919 33853
rect 32861 33813 32873 33847
rect 32907 33844 32919 33847
rect 33520 33844 33548 33875
rect 33962 33844 33968 33856
rect 32907 33816 33968 33844
rect 32907 33813 32919 33816
rect 32861 33807 32919 33813
rect 33962 33804 33968 33816
rect 34020 33844 34026 33856
rect 34072 33853 34100 33884
rect 34793 33881 34805 33884
rect 34839 33881 34851 33915
rect 34793 33875 34851 33881
rect 34977 33915 35035 33921
rect 34977 33881 34989 33915
rect 35023 33912 35035 33915
rect 35023 33884 35894 33912
rect 35023 33881 35035 33884
rect 34977 33875 35035 33881
rect 34057 33847 34115 33853
rect 34057 33844 34069 33847
rect 34020 33816 34069 33844
rect 34020 33804 34026 33816
rect 34057 33813 34069 33816
rect 34103 33813 34115 33847
rect 34057 33807 34115 33813
rect 34698 33804 34704 33856
rect 34756 33844 34762 33856
rect 35437 33847 35495 33853
rect 35437 33844 35449 33847
rect 34756 33816 35449 33844
rect 34756 33804 34762 33816
rect 35437 33813 35449 33816
rect 35483 33813 35495 33847
rect 35866 33844 35894 33884
rect 77312 33856 77340 33952
rect 77849 33949 77861 33952
rect 77895 33949 77907 33983
rect 77849 33943 77907 33949
rect 77110 33844 77116 33856
rect 35866 33816 77116 33844
rect 35437 33807 35495 33813
rect 77110 33804 77116 33816
rect 77168 33804 77174 33856
rect 77294 33844 77300 33856
rect 77255 33816 77300 33844
rect 77294 33804 77300 33816
rect 77352 33804 77358 33856
rect 78030 33844 78036 33856
rect 77991 33816 78036 33844
rect 78030 33804 78036 33816
rect 78088 33804 78094 33856
rect 1104 33754 78844 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 78844 33754
rect 1104 33680 78844 33702
rect 32674 33640 32680 33652
rect 32635 33612 32680 33640
rect 32674 33600 32680 33612
rect 32732 33600 32738 33652
rect 32769 33507 32827 33513
rect 32769 33473 32781 33507
rect 32815 33504 32827 33507
rect 33226 33504 33232 33516
rect 32815 33476 33232 33504
rect 32815 33473 32827 33476
rect 32769 33467 32827 33473
rect 33226 33464 33232 33476
rect 33284 33504 33290 33516
rect 33689 33507 33747 33513
rect 33689 33504 33701 33507
rect 33284 33476 33701 33504
rect 33284 33464 33290 33476
rect 33689 33473 33701 33476
rect 33735 33504 33747 33507
rect 34333 33507 34391 33513
rect 34333 33504 34345 33507
rect 33735 33476 34345 33504
rect 33735 33473 33747 33476
rect 33689 33467 33747 33473
rect 34333 33473 34345 33476
rect 34379 33473 34391 33507
rect 34333 33467 34391 33473
rect 33873 33371 33931 33377
rect 33873 33337 33885 33371
rect 33919 33368 33931 33371
rect 33919 33340 35894 33368
rect 33919 33337 33931 33340
rect 33873 33331 33931 33337
rect 35866 33300 35894 33340
rect 77294 33300 77300 33312
rect 35866 33272 77300 33300
rect 77294 33260 77300 33272
rect 77352 33260 77358 33312
rect 1104 33210 78844 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 78844 33210
rect 1104 33136 78844 33158
rect 1673 32895 1731 32901
rect 1673 32861 1685 32895
rect 1719 32861 1731 32895
rect 77849 32895 77907 32901
rect 77849 32892 77861 32895
rect 1673 32855 1731 32861
rect 77312 32864 77861 32892
rect 1688 32824 1716 32855
rect 2225 32827 2283 32833
rect 2225 32824 2237 32827
rect 1688 32796 2237 32824
rect 2225 32793 2237 32796
rect 2271 32824 2283 32827
rect 32214 32824 32220 32836
rect 2271 32796 32220 32824
rect 2271 32793 2283 32796
rect 2225 32787 2283 32793
rect 32214 32784 32220 32796
rect 32272 32784 32278 32836
rect 1486 32756 1492 32768
rect 1447 32728 1492 32756
rect 1486 32716 1492 32728
rect 1544 32716 1550 32768
rect 32769 32759 32827 32765
rect 32769 32725 32781 32759
rect 32815 32756 32827 32759
rect 32950 32756 32956 32768
rect 32815 32728 32956 32756
rect 32815 32725 32827 32728
rect 32769 32719 32827 32725
rect 32950 32716 32956 32728
rect 33008 32716 33014 32768
rect 33226 32716 33232 32768
rect 33284 32756 33290 32768
rect 33413 32759 33471 32765
rect 33413 32756 33425 32759
rect 33284 32728 33425 32756
rect 33284 32716 33290 32728
rect 33413 32725 33425 32728
rect 33459 32725 33471 32759
rect 33413 32719 33471 32725
rect 77018 32716 77024 32768
rect 77076 32756 77082 32768
rect 77312 32765 77340 32864
rect 77849 32861 77861 32864
rect 77895 32861 77907 32895
rect 77849 32855 77907 32861
rect 77297 32759 77355 32765
rect 77297 32756 77309 32759
rect 77076 32728 77309 32756
rect 77076 32716 77082 32728
rect 77297 32725 77309 32728
rect 77343 32725 77355 32759
rect 78030 32756 78036 32768
rect 77991 32728 78036 32756
rect 77297 32719 77355 32725
rect 78030 32716 78036 32728
rect 78088 32716 78094 32768
rect 1104 32666 78844 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 78844 32666
rect 1104 32592 78844 32614
rect 32214 32552 32220 32564
rect 32175 32524 32220 32552
rect 32214 32512 32220 32524
rect 32272 32512 32278 32564
rect 1673 32419 1731 32425
rect 1673 32385 1685 32419
rect 1719 32416 1731 32419
rect 2225 32419 2283 32425
rect 2225 32416 2237 32419
rect 1719 32388 2237 32416
rect 1719 32385 1731 32388
rect 1673 32379 1731 32385
rect 2225 32385 2237 32388
rect 2271 32416 2283 32419
rect 31202 32416 31208 32428
rect 2271 32388 31208 32416
rect 2271 32385 2283 32388
rect 2225 32379 2283 32385
rect 31202 32376 31208 32388
rect 31260 32376 31266 32428
rect 32309 32419 32367 32425
rect 32309 32385 32321 32419
rect 32355 32416 32367 32419
rect 32950 32416 32956 32428
rect 32355 32388 32956 32416
rect 32355 32385 32367 32388
rect 32309 32379 32367 32385
rect 32950 32376 32956 32388
rect 33008 32376 33014 32428
rect 77665 32419 77723 32425
rect 77665 32416 77677 32419
rect 77128 32388 77677 32416
rect 33137 32283 33195 32289
rect 33137 32249 33149 32283
rect 33183 32280 33195 32283
rect 77018 32280 77024 32292
rect 33183 32252 77024 32280
rect 33183 32249 33195 32252
rect 33137 32243 33195 32249
rect 77018 32240 77024 32252
rect 77076 32240 77082 32292
rect 1486 32212 1492 32224
rect 1447 32184 1492 32212
rect 1486 32172 1492 32184
rect 1544 32172 1550 32224
rect 69658 32172 69664 32224
rect 69716 32212 69722 32224
rect 77128 32221 77156 32388
rect 77665 32385 77677 32388
rect 77711 32385 77723 32419
rect 77665 32379 77723 32385
rect 77113 32215 77171 32221
rect 77113 32212 77125 32215
rect 69716 32184 77125 32212
rect 69716 32172 69722 32184
rect 77113 32181 77125 32184
rect 77159 32181 77171 32215
rect 77846 32212 77852 32224
rect 77807 32184 77852 32212
rect 77113 32175 77171 32181
rect 77846 32172 77852 32184
rect 77904 32172 77910 32224
rect 1104 32122 78844 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 78844 32122
rect 1104 32048 78844 32070
rect 31202 32008 31208 32020
rect 31163 31980 31208 32008
rect 31202 31968 31208 31980
rect 31260 31968 31266 32020
rect 32398 31900 32404 31952
rect 32456 31940 32462 31952
rect 77297 31943 77355 31949
rect 77297 31940 77309 31943
rect 32456 31912 77309 31940
rect 32456 31900 32462 31912
rect 77297 31909 77309 31912
rect 77343 31909 77355 31943
rect 78030 31940 78036 31952
rect 77991 31912 78036 31940
rect 77297 31903 77355 31909
rect 32493 31875 32551 31881
rect 32493 31841 32505 31875
rect 32539 31872 32551 31875
rect 69658 31872 69664 31884
rect 32539 31844 69664 31872
rect 32539 31841 32551 31844
rect 32493 31835 32551 31841
rect 69658 31832 69664 31844
rect 69716 31832 69722 31884
rect 1673 31807 1731 31813
rect 1673 31773 1685 31807
rect 1719 31804 1731 31807
rect 2225 31807 2283 31813
rect 2225 31804 2237 31807
rect 1719 31776 2237 31804
rect 1719 31773 1731 31776
rect 1673 31767 1731 31773
rect 2225 31773 2237 31776
rect 2271 31804 2283 31807
rect 2314 31804 2320 31816
rect 2271 31776 2320 31804
rect 2271 31773 2283 31776
rect 2225 31767 2283 31773
rect 2314 31764 2320 31776
rect 2372 31764 2378 31816
rect 32582 31764 32588 31816
rect 32640 31804 32646 31816
rect 32950 31804 32956 31816
rect 32640 31776 32956 31804
rect 32640 31764 32646 31776
rect 32950 31764 32956 31776
rect 33008 31764 33014 31816
rect 77312 31804 77340 31903
rect 78030 31900 78036 31912
rect 78088 31900 78094 31952
rect 77849 31807 77907 31813
rect 77849 31804 77861 31807
rect 77312 31776 77861 31804
rect 77849 31773 77861 31776
rect 77895 31773 77907 31807
rect 77849 31767 77907 31773
rect 31297 31739 31355 31745
rect 31297 31705 31309 31739
rect 31343 31736 31355 31739
rect 31938 31736 31944 31748
rect 31343 31708 31944 31736
rect 31343 31705 31355 31708
rect 31297 31699 31355 31705
rect 31938 31696 31944 31708
rect 31996 31736 32002 31748
rect 32309 31739 32367 31745
rect 32309 31736 32321 31739
rect 31996 31708 32321 31736
rect 31996 31696 32002 31708
rect 32309 31705 32321 31708
rect 32355 31705 32367 31739
rect 32309 31699 32367 31705
rect 1486 31668 1492 31680
rect 1447 31640 1492 31668
rect 1486 31628 1492 31640
rect 1544 31628 1550 31680
rect 1104 31578 78844 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 78844 31578
rect 1104 31504 78844 31526
rect 32398 31396 32404 31408
rect 32359 31368 32404 31396
rect 32398 31356 32404 31368
rect 32456 31356 32462 31408
rect 1673 31331 1731 31337
rect 1673 31297 1685 31331
rect 1719 31328 1731 31331
rect 29917 31331 29975 31337
rect 1719 31300 2268 31328
rect 1719 31297 1731 31300
rect 1673 31291 1731 31297
rect 2240 31201 2268 31300
rect 29917 31297 29929 31331
rect 29963 31328 29975 31331
rect 30561 31331 30619 31337
rect 30561 31328 30573 31331
rect 29963 31300 30573 31328
rect 29963 31297 29975 31300
rect 29917 31291 29975 31297
rect 30561 31297 30573 31300
rect 30607 31328 30619 31331
rect 31662 31328 31668 31340
rect 30607 31300 31668 31328
rect 30607 31297 30619 31300
rect 30561 31291 30619 31297
rect 31662 31288 31668 31300
rect 31720 31328 31726 31340
rect 32217 31331 32275 31337
rect 32217 31328 32229 31331
rect 31720 31300 32229 31328
rect 31720 31288 31726 31300
rect 32217 31297 32229 31300
rect 32263 31297 32275 31331
rect 77665 31331 77723 31337
rect 77665 31328 77677 31331
rect 32217 31291 32275 31297
rect 77128 31300 77677 31328
rect 2314 31220 2320 31272
rect 2372 31260 2378 31272
rect 30377 31263 30435 31269
rect 30377 31260 30389 31263
rect 2372 31232 30389 31260
rect 2372 31220 2378 31232
rect 30377 31229 30389 31232
rect 30423 31229 30435 31263
rect 30377 31223 30435 31229
rect 2225 31195 2283 31201
rect 2225 31161 2237 31195
rect 2271 31192 2283 31195
rect 29730 31192 29736 31204
rect 2271 31164 29736 31192
rect 2271 31161 2283 31164
rect 2225 31155 2283 31161
rect 29730 31152 29736 31164
rect 29788 31152 29794 31204
rect 1486 31124 1492 31136
rect 1447 31096 1492 31124
rect 1486 31084 1492 31096
rect 1544 31084 1550 31136
rect 31573 31127 31631 31133
rect 31573 31093 31585 31127
rect 31619 31124 31631 31127
rect 31938 31124 31944 31136
rect 31619 31096 31944 31124
rect 31619 31093 31631 31096
rect 31573 31087 31631 31093
rect 31938 31084 31944 31096
rect 31996 31124 32002 31136
rect 32861 31127 32919 31133
rect 32861 31124 32873 31127
rect 31996 31096 32873 31124
rect 31996 31084 32002 31096
rect 32861 31093 32873 31096
rect 32907 31093 32919 31127
rect 32861 31087 32919 31093
rect 68002 31084 68008 31136
rect 68060 31124 68066 31136
rect 77128 31133 77156 31300
rect 77665 31297 77677 31300
rect 77711 31297 77723 31331
rect 77665 31291 77723 31297
rect 77113 31127 77171 31133
rect 77113 31124 77125 31127
rect 68060 31096 77125 31124
rect 68060 31084 68066 31096
rect 77113 31093 77125 31096
rect 77159 31093 77171 31127
rect 77846 31124 77852 31136
rect 77807 31096 77852 31124
rect 77113 31087 77171 31093
rect 77846 31084 77852 31096
rect 77904 31084 77910 31136
rect 1104 31034 78844 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 78844 31034
rect 1104 30960 78844 30982
rect 29730 30920 29736 30932
rect 29691 30892 29736 30920
rect 29730 30880 29736 30892
rect 29788 30880 29794 30932
rect 29825 30651 29883 30657
rect 29825 30617 29837 30651
rect 29871 30648 29883 30651
rect 30374 30648 30380 30660
rect 29871 30620 30380 30648
rect 29871 30617 29883 30620
rect 29825 30611 29883 30617
rect 30374 30608 30380 30620
rect 30432 30648 30438 30660
rect 30929 30651 30987 30657
rect 30929 30648 30941 30651
rect 30432 30620 30941 30648
rect 30432 30608 30438 30620
rect 30929 30617 30941 30620
rect 30975 30617 30987 30651
rect 30929 30611 30987 30617
rect 31113 30651 31171 30657
rect 31113 30617 31125 30651
rect 31159 30648 31171 30651
rect 31159 30620 35894 30648
rect 31159 30617 31171 30620
rect 31113 30611 31171 30617
rect 31018 30540 31024 30592
rect 31076 30580 31082 30592
rect 31662 30580 31668 30592
rect 31076 30552 31668 30580
rect 31076 30540 31082 30552
rect 31662 30540 31668 30552
rect 31720 30580 31726 30592
rect 31941 30583 31999 30589
rect 31941 30580 31953 30583
rect 31720 30552 31953 30580
rect 31720 30540 31726 30552
rect 31941 30549 31953 30552
rect 31987 30549 31999 30583
rect 35866 30580 35894 30620
rect 68002 30580 68008 30592
rect 35866 30552 68008 30580
rect 31941 30543 31999 30549
rect 68002 30540 68008 30552
rect 68060 30540 68066 30592
rect 1104 30490 78844 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 78844 30490
rect 1104 30416 78844 30438
rect 1673 30243 1731 30249
rect 1673 30209 1685 30243
rect 1719 30240 1731 30243
rect 77665 30243 77723 30249
rect 77665 30240 77677 30243
rect 1719 30212 2268 30240
rect 1719 30209 1731 30212
rect 1673 30203 1731 30209
rect 1486 30104 1492 30116
rect 1447 30076 1492 30104
rect 1486 30064 1492 30076
rect 1544 30064 1550 30116
rect 2240 30113 2268 30212
rect 77128 30212 77677 30240
rect 2225 30107 2283 30113
rect 2225 30073 2237 30107
rect 2271 30104 2283 30107
rect 28810 30104 28816 30116
rect 2271 30076 28816 30104
rect 2271 30073 2283 30076
rect 2225 30067 2283 30073
rect 28810 30064 28816 30076
rect 28868 30064 28874 30116
rect 29181 30039 29239 30045
rect 29181 30005 29193 30039
rect 29227 30036 29239 30039
rect 29362 30036 29368 30048
rect 29227 30008 29368 30036
rect 29227 30005 29239 30008
rect 29181 29999 29239 30005
rect 29362 29996 29368 30008
rect 29420 29996 29426 30048
rect 30101 30039 30159 30045
rect 30101 30005 30113 30039
rect 30147 30036 30159 30039
rect 30374 30036 30380 30048
rect 30147 30008 30380 30036
rect 30147 30005 30159 30008
rect 30101 29999 30159 30005
rect 30374 29996 30380 30008
rect 30432 30036 30438 30048
rect 30653 30039 30711 30045
rect 30653 30036 30665 30039
rect 30432 30008 30665 30036
rect 30432 29996 30438 30008
rect 30653 30005 30665 30008
rect 30699 30005 30711 30039
rect 30653 29999 30711 30005
rect 69658 29996 69664 30048
rect 69716 30036 69722 30048
rect 77128 30045 77156 30212
rect 77665 30209 77677 30212
rect 77711 30209 77723 30243
rect 77665 30203 77723 30209
rect 77846 30104 77852 30116
rect 77807 30076 77852 30104
rect 77846 30064 77852 30076
rect 77904 30064 77910 30116
rect 77113 30039 77171 30045
rect 77113 30036 77125 30039
rect 69716 30008 77125 30036
rect 69716 29996 69722 30008
rect 77113 30005 77125 30008
rect 77159 30005 77171 30039
rect 77113 29999 77171 30005
rect 1104 29946 78844 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 78844 29946
rect 1104 29872 78844 29894
rect 28810 29832 28816 29844
rect 28771 29804 28816 29832
rect 28810 29792 28816 29804
rect 28868 29792 28874 29844
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29628 1731 29631
rect 2225 29631 2283 29637
rect 2225 29628 2237 29631
rect 1719 29600 2237 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 2225 29597 2237 29600
rect 2271 29628 2283 29631
rect 28258 29628 28264 29640
rect 2271 29600 28264 29628
rect 2271 29597 2283 29600
rect 2225 29591 2283 29597
rect 28258 29588 28264 29600
rect 28316 29588 28322 29640
rect 77849 29631 77907 29637
rect 77849 29628 77861 29631
rect 77312 29600 77861 29628
rect 28905 29563 28963 29569
rect 28905 29529 28917 29563
rect 28951 29529 28963 29563
rect 28905 29523 28963 29529
rect 30193 29563 30251 29569
rect 30193 29529 30205 29563
rect 30239 29529 30251 29563
rect 30193 29523 30251 29529
rect 30377 29563 30435 29569
rect 30377 29529 30389 29563
rect 30423 29560 30435 29563
rect 30423 29532 35894 29560
rect 30423 29529 30435 29532
rect 30377 29523 30435 29529
rect 1486 29492 1492 29504
rect 1447 29464 1492 29492
rect 1486 29452 1492 29464
rect 1544 29452 1550 29504
rect 28920 29492 28948 29523
rect 29362 29492 29368 29504
rect 28920 29464 29368 29492
rect 29362 29452 29368 29464
rect 29420 29492 29426 29504
rect 29549 29495 29607 29501
rect 29549 29492 29561 29495
rect 29420 29464 29561 29492
rect 29420 29452 29426 29464
rect 29549 29461 29561 29464
rect 29595 29492 29607 29495
rect 30208 29492 30236 29523
rect 29595 29464 30236 29492
rect 35866 29492 35894 29532
rect 77312 29504 77340 29600
rect 77849 29597 77861 29600
rect 77895 29597 77907 29631
rect 77849 29591 77907 29597
rect 69658 29492 69664 29504
rect 35866 29464 69664 29492
rect 29595 29461 29607 29464
rect 29549 29455 29607 29461
rect 69658 29452 69664 29464
rect 69716 29452 69722 29504
rect 77294 29492 77300 29504
rect 77255 29464 77300 29492
rect 77294 29452 77300 29464
rect 77352 29452 77358 29504
rect 78030 29492 78036 29504
rect 77991 29464 78036 29492
rect 78030 29452 78036 29464
rect 78088 29452 78094 29504
rect 1104 29402 78844 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 78844 29402
rect 1104 29328 78844 29350
rect 28258 29288 28264 29300
rect 28219 29260 28264 29288
rect 28258 29248 28264 29260
rect 28316 29248 28322 29300
rect 1673 29155 1731 29161
rect 1673 29121 1685 29155
rect 1719 29152 1731 29155
rect 27709 29155 27767 29161
rect 1719 29124 2268 29152
rect 1719 29121 1731 29124
rect 1673 29115 1731 29121
rect 2240 29093 2268 29124
rect 27709 29121 27721 29155
rect 27755 29152 27767 29155
rect 28353 29155 28411 29161
rect 28353 29152 28365 29155
rect 27755 29124 28365 29152
rect 27755 29121 27767 29124
rect 27709 29115 27767 29121
rect 28353 29121 28365 29124
rect 28399 29152 28411 29155
rect 29549 29155 29607 29161
rect 29549 29152 29561 29155
rect 28399 29124 29561 29152
rect 28399 29121 28411 29124
rect 28353 29115 28411 29121
rect 2225 29087 2283 29093
rect 2225 29053 2237 29087
rect 2271 29084 2283 29087
rect 26142 29084 26148 29096
rect 2271 29056 26148 29084
rect 2271 29053 2283 29056
rect 2225 29047 2283 29053
rect 26142 29044 26148 29056
rect 26200 29044 26206 29096
rect 28736 29028 28764 29124
rect 29549 29121 29561 29124
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 29733 29155 29791 29161
rect 29733 29121 29745 29155
rect 29779 29152 29791 29155
rect 77294 29152 77300 29164
rect 29779 29124 77300 29152
rect 29779 29121 29791 29124
rect 29733 29115 29791 29121
rect 77294 29112 77300 29124
rect 77352 29112 77358 29164
rect 77665 29155 77723 29161
rect 77665 29121 77677 29155
rect 77711 29121 77723 29155
rect 77665 29115 77723 29121
rect 77680 29084 77708 29115
rect 77128 29056 77708 29084
rect 77128 29028 77156 29056
rect 1486 29016 1492 29028
rect 1447 28988 1492 29016
rect 1486 28976 1492 28988
rect 1544 28976 1550 29028
rect 28718 28976 28724 29028
rect 28776 29016 28782 29028
rect 28905 29019 28963 29025
rect 28905 29016 28917 29019
rect 28776 28988 28917 29016
rect 28776 28976 28782 28988
rect 28905 28985 28917 28988
rect 28951 28985 28963 29019
rect 77110 29016 77116 29028
rect 77071 28988 77116 29016
rect 28905 28979 28963 28985
rect 77110 28976 77116 28988
rect 77168 28976 77174 29028
rect 77846 29016 77852 29028
rect 77807 28988 77852 29016
rect 77846 28976 77852 28988
rect 77904 28976 77910 29028
rect 1104 28858 78844 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 78844 28858
rect 1104 28784 78844 28806
rect 26142 28636 26148 28688
rect 26200 28676 26206 28688
rect 27433 28679 27491 28685
rect 27433 28676 27445 28679
rect 26200 28648 27445 28676
rect 26200 28636 26206 28648
rect 27433 28645 27445 28648
rect 27479 28645 27491 28679
rect 27433 28639 27491 28645
rect 1673 28543 1731 28549
rect 1673 28509 1685 28543
rect 1719 28540 1731 28543
rect 2225 28543 2283 28549
rect 2225 28540 2237 28543
rect 1719 28512 2237 28540
rect 1719 28509 1731 28512
rect 1673 28503 1731 28509
rect 2225 28509 2237 28512
rect 2271 28540 2283 28543
rect 27062 28540 27068 28552
rect 2271 28512 27068 28540
rect 2271 28509 2283 28512
rect 2225 28503 2283 28509
rect 27062 28500 27068 28512
rect 27120 28500 27126 28552
rect 77849 28543 77907 28549
rect 77849 28540 77861 28543
rect 77312 28512 77861 28540
rect 26973 28475 27031 28481
rect 26973 28441 26985 28475
rect 27019 28472 27031 28475
rect 27617 28475 27675 28481
rect 27617 28472 27629 28475
rect 27019 28444 27629 28472
rect 27019 28441 27031 28444
rect 26973 28435 27031 28441
rect 27617 28441 27629 28444
rect 27663 28472 27675 28475
rect 28813 28475 28871 28481
rect 28813 28472 28825 28475
rect 27663 28444 28825 28472
rect 27663 28441 27675 28444
rect 27617 28435 27675 28441
rect 28000 28416 28028 28444
rect 28813 28441 28825 28444
rect 28859 28441 28871 28475
rect 28813 28435 28871 28441
rect 28997 28475 29055 28481
rect 28997 28441 29009 28475
rect 29043 28472 29055 28475
rect 29043 28444 35894 28472
rect 29043 28441 29055 28444
rect 28997 28435 29055 28441
rect 1486 28404 1492 28416
rect 1447 28376 1492 28404
rect 1486 28364 1492 28376
rect 1544 28364 1550 28416
rect 27982 28364 27988 28416
rect 28040 28404 28046 28416
rect 28169 28407 28227 28413
rect 28169 28404 28181 28407
rect 28040 28376 28181 28404
rect 28040 28364 28046 28376
rect 28169 28373 28181 28376
rect 28215 28373 28227 28407
rect 35866 28404 35894 28444
rect 77312 28416 77340 28512
rect 77849 28509 77861 28512
rect 77895 28509 77907 28543
rect 77849 28503 77907 28509
rect 77110 28404 77116 28416
rect 35866 28376 77116 28404
rect 28169 28367 28227 28373
rect 77110 28364 77116 28376
rect 77168 28364 77174 28416
rect 77294 28404 77300 28416
rect 77255 28376 77300 28404
rect 77294 28364 77300 28376
rect 77352 28364 77358 28416
rect 78030 28404 78036 28416
rect 77991 28376 78036 28404
rect 78030 28364 78036 28376
rect 78088 28364 78094 28416
rect 1104 28314 78844 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 78844 28314
rect 1104 28240 78844 28262
rect 27062 28200 27068 28212
rect 27023 28172 27068 28200
rect 27062 28160 27068 28172
rect 27120 28160 27126 28212
rect 27157 28067 27215 28073
rect 27157 28033 27169 28067
rect 27203 28064 27215 28067
rect 27430 28064 27436 28076
rect 27203 28036 27436 28064
rect 27203 28033 27215 28036
rect 27157 28027 27215 28033
rect 27430 28024 27436 28036
rect 27488 28064 27494 28076
rect 28169 28067 28227 28073
rect 28169 28064 28181 28067
rect 27488 28036 28181 28064
rect 27488 28024 27494 28036
rect 28169 28033 28181 28036
rect 28215 28033 28227 28067
rect 28169 28027 28227 28033
rect 28261 27863 28319 27869
rect 28261 27829 28273 27863
rect 28307 27860 28319 27863
rect 77294 27860 77300 27872
rect 28307 27832 77300 27860
rect 28307 27829 28319 27832
rect 28261 27823 28319 27829
rect 77294 27820 77300 27832
rect 77352 27820 77358 27872
rect 1104 27770 78844 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 78844 27770
rect 1104 27696 78844 27718
rect 1673 27455 1731 27461
rect 1673 27421 1685 27455
rect 1719 27452 1731 27455
rect 2225 27455 2283 27461
rect 2225 27452 2237 27455
rect 1719 27424 2237 27452
rect 1719 27421 1731 27424
rect 1673 27415 1731 27421
rect 2225 27421 2237 27424
rect 2271 27452 2283 27455
rect 26050 27452 26056 27464
rect 2271 27424 26056 27452
rect 2271 27421 2283 27424
rect 2225 27415 2283 27421
rect 26050 27412 26056 27424
rect 26108 27412 26114 27464
rect 77849 27455 77907 27461
rect 77849 27452 77861 27455
rect 77312 27424 77861 27452
rect 1486 27316 1492 27328
rect 1447 27288 1492 27316
rect 1486 27276 1492 27288
rect 1544 27276 1550 27328
rect 26142 27276 26148 27328
rect 26200 27316 26206 27328
rect 26329 27319 26387 27325
rect 26329 27316 26341 27319
rect 26200 27288 26341 27316
rect 26200 27276 26206 27288
rect 26329 27285 26341 27288
rect 26375 27285 26387 27319
rect 27430 27316 27436 27328
rect 27391 27288 27436 27316
rect 26329 27279 26387 27285
rect 27430 27276 27436 27288
rect 27488 27316 27494 27328
rect 27893 27319 27951 27325
rect 27893 27316 27905 27319
rect 27488 27288 27905 27316
rect 27488 27276 27494 27288
rect 27893 27285 27905 27288
rect 27939 27285 27951 27319
rect 27893 27279 27951 27285
rect 77018 27276 77024 27328
rect 77076 27316 77082 27328
rect 77312 27325 77340 27424
rect 77849 27421 77861 27424
rect 77895 27421 77907 27455
rect 77849 27415 77907 27421
rect 77297 27319 77355 27325
rect 77297 27316 77309 27319
rect 77076 27288 77309 27316
rect 77076 27276 77082 27288
rect 77297 27285 77309 27288
rect 77343 27285 77355 27319
rect 78030 27316 78036 27328
rect 77991 27288 78036 27316
rect 77297 27279 77355 27285
rect 78030 27276 78036 27288
rect 78088 27276 78094 27328
rect 1104 27226 78844 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 78844 27226
rect 1104 27152 78844 27174
rect 26050 27112 26056 27124
rect 26011 27084 26056 27112
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 1673 26979 1731 26985
rect 1673 26945 1685 26979
rect 1719 26976 1731 26979
rect 2225 26979 2283 26985
rect 2225 26976 2237 26979
rect 1719 26948 2237 26976
rect 1719 26945 1731 26948
rect 1673 26939 1731 26945
rect 2225 26945 2237 26948
rect 2271 26976 2283 26979
rect 25222 26976 25228 26988
rect 2271 26948 25228 26976
rect 2271 26945 2283 26948
rect 2225 26939 2283 26945
rect 25222 26936 25228 26948
rect 25280 26936 25286 26988
rect 26142 26976 26148 26988
rect 26103 26948 26148 26976
rect 26142 26936 26148 26948
rect 26200 26976 26206 26988
rect 27433 26979 27491 26985
rect 27433 26976 27445 26979
rect 26200 26948 27445 26976
rect 26200 26936 26206 26948
rect 27433 26945 27445 26948
rect 27479 26945 27491 26979
rect 77665 26979 77723 26985
rect 77665 26976 77677 26979
rect 27433 26939 27491 26945
rect 77128 26948 77677 26976
rect 27617 26843 27675 26849
rect 27617 26809 27629 26843
rect 27663 26840 27675 26843
rect 77018 26840 77024 26852
rect 27663 26812 77024 26840
rect 27663 26809 27675 26812
rect 27617 26803 27675 26809
rect 77018 26800 77024 26812
rect 77076 26800 77082 26852
rect 1486 26772 1492 26784
rect 1447 26744 1492 26772
rect 1486 26732 1492 26744
rect 1544 26732 1550 26784
rect 69658 26732 69664 26784
rect 69716 26772 69722 26784
rect 77128 26781 77156 26948
rect 77665 26945 77677 26948
rect 77711 26945 77723 26979
rect 77665 26939 77723 26945
rect 77113 26775 77171 26781
rect 77113 26772 77125 26775
rect 69716 26744 77125 26772
rect 69716 26732 69722 26744
rect 77113 26741 77125 26744
rect 77159 26741 77171 26775
rect 77846 26772 77852 26784
rect 77807 26744 77852 26772
rect 77113 26735 77171 26741
rect 77846 26732 77852 26744
rect 77904 26732 77910 26784
rect 1104 26682 78844 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 78844 26682
rect 1104 26608 78844 26630
rect 25222 26568 25228 26580
rect 25183 26540 25228 26568
rect 25222 26528 25228 26540
rect 25280 26528 25286 26580
rect 78030 26500 78036 26512
rect 77991 26472 78036 26500
rect 78030 26460 78036 26472
rect 78088 26460 78094 26512
rect 26142 26392 26148 26444
rect 26200 26432 26206 26444
rect 27341 26435 27399 26441
rect 27341 26432 27353 26435
rect 26200 26404 27353 26432
rect 26200 26392 26206 26404
rect 27341 26401 27353 26404
rect 27387 26401 27399 26435
rect 27341 26395 27399 26401
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26364 1731 26367
rect 2225 26367 2283 26373
rect 2225 26364 2237 26367
rect 1719 26336 2237 26364
rect 1719 26333 1731 26336
rect 1673 26327 1731 26333
rect 2225 26333 2237 26336
rect 2271 26364 2283 26367
rect 22830 26364 22836 26376
rect 2271 26336 22836 26364
rect 2271 26333 2283 26336
rect 2225 26327 2283 26333
rect 22830 26324 22836 26336
rect 22888 26324 22894 26376
rect 26881 26367 26939 26373
rect 26881 26333 26893 26367
rect 26927 26364 26939 26367
rect 77386 26364 77392 26376
rect 26927 26336 35894 26364
rect 77299 26336 77392 26364
rect 26927 26333 26939 26336
rect 26881 26327 26939 26333
rect 25317 26299 25375 26305
rect 25317 26265 25329 26299
rect 25363 26265 25375 26299
rect 26697 26299 26755 26305
rect 26697 26296 26709 26299
rect 25317 26259 25375 26265
rect 26068 26268 26709 26296
rect 1486 26228 1492 26240
rect 1447 26200 1492 26228
rect 1486 26188 1492 26200
rect 1544 26188 1550 26240
rect 25332 26228 25360 26259
rect 26068 26240 26096 26268
rect 26697 26265 26709 26268
rect 26743 26265 26755 26299
rect 35866 26296 35894 26336
rect 77386 26324 77392 26336
rect 77444 26364 77450 26376
rect 77849 26367 77907 26373
rect 77849 26364 77861 26367
rect 77444 26336 77861 26364
rect 77444 26324 77450 26336
rect 77849 26333 77861 26336
rect 77895 26333 77907 26367
rect 77849 26327 77907 26333
rect 69658 26296 69664 26308
rect 35866 26268 69664 26296
rect 26697 26259 26755 26265
rect 69658 26256 69664 26268
rect 69716 26256 69722 26308
rect 26050 26228 26056 26240
rect 25332 26200 26056 26228
rect 26050 26188 26056 26200
rect 26108 26188 26114 26240
rect 32493 26231 32551 26237
rect 32493 26197 32505 26231
rect 32539 26228 32551 26231
rect 32674 26228 32680 26240
rect 32539 26200 32680 26228
rect 32539 26197 32551 26200
rect 32493 26191 32551 26197
rect 32674 26188 32680 26200
rect 32732 26188 32738 26240
rect 1104 26138 78844 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 78844 26138
rect 1104 26064 78844 26086
rect 22830 25956 22836 25968
rect 22791 25928 22836 25956
rect 22830 25916 22836 25928
rect 22888 25916 22894 25968
rect 31662 25916 31668 25968
rect 31720 25956 31726 25968
rect 32674 25956 32680 25968
rect 31720 25928 32680 25956
rect 31720 25916 31726 25928
rect 32674 25916 32680 25928
rect 32732 25916 32738 25968
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25888 1731 25891
rect 23017 25891 23075 25897
rect 1719 25860 2268 25888
rect 1719 25857 1731 25860
rect 1673 25851 1731 25857
rect 2240 25761 2268 25860
rect 23017 25857 23029 25891
rect 23063 25888 23075 25891
rect 23569 25891 23627 25897
rect 23569 25888 23581 25891
rect 23063 25860 23581 25888
rect 23063 25857 23075 25860
rect 23017 25851 23075 25857
rect 23569 25857 23581 25860
rect 23615 25888 23627 25891
rect 24946 25888 24952 25900
rect 23615 25860 24952 25888
rect 23615 25857 23627 25860
rect 23569 25851 23627 25857
rect 24946 25848 24952 25860
rect 25004 25848 25010 25900
rect 77665 25891 77723 25897
rect 77665 25888 77677 25891
rect 77128 25860 77677 25888
rect 2225 25755 2283 25761
rect 2225 25721 2237 25755
rect 2271 25752 2283 25755
rect 22278 25752 22284 25764
rect 2271 25724 22284 25752
rect 2271 25721 2283 25724
rect 2225 25715 2283 25721
rect 22278 25712 22284 25724
rect 22336 25712 22342 25764
rect 69658 25712 69664 25764
rect 69716 25752 69722 25764
rect 77128 25761 77156 25860
rect 77665 25857 77677 25860
rect 77711 25857 77723 25891
rect 77665 25851 77723 25857
rect 77113 25755 77171 25761
rect 77113 25752 77125 25755
rect 69716 25724 77125 25752
rect 69716 25712 69722 25724
rect 77113 25721 77125 25724
rect 77159 25721 77171 25755
rect 77113 25715 77171 25721
rect 1486 25684 1492 25696
rect 1447 25656 1492 25684
rect 1486 25644 1492 25656
rect 1544 25644 1550 25696
rect 25593 25687 25651 25693
rect 25593 25653 25605 25687
rect 25639 25684 25651 25687
rect 26050 25684 26056 25696
rect 25639 25656 26056 25684
rect 25639 25653 25651 25656
rect 25593 25647 25651 25653
rect 26050 25644 26056 25656
rect 26108 25644 26114 25696
rect 32769 25687 32827 25693
rect 32769 25653 32781 25687
rect 32815 25684 32827 25687
rect 77386 25684 77392 25696
rect 32815 25656 77392 25684
rect 32815 25653 32827 25656
rect 32769 25647 32827 25653
rect 77386 25644 77392 25656
rect 77444 25644 77450 25696
rect 77846 25684 77852 25696
rect 77807 25656 77852 25684
rect 77846 25644 77852 25656
rect 77904 25644 77910 25696
rect 1104 25594 78844 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 78844 25594
rect 1104 25520 78844 25542
rect 22278 25480 22284 25492
rect 22239 25452 22284 25480
rect 22278 25440 22284 25452
rect 22336 25440 22342 25492
rect 22465 25279 22523 25285
rect 22465 25245 22477 25279
rect 22511 25276 22523 25279
rect 22925 25279 22983 25285
rect 22925 25276 22937 25279
rect 22511 25248 22937 25276
rect 22511 25245 22523 25248
rect 22465 25239 22523 25245
rect 22925 25245 22937 25248
rect 22971 25276 22983 25279
rect 24394 25276 24400 25288
rect 22971 25248 24400 25276
rect 22971 25245 22983 25248
rect 22925 25239 22983 25245
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 32585 25211 32643 25217
rect 32585 25208 32597 25211
rect 31956 25180 32597 25208
rect 30834 25100 30840 25152
rect 30892 25140 30898 25152
rect 31956 25149 31984 25180
rect 32585 25177 32597 25180
rect 32631 25177 32643 25211
rect 32585 25171 32643 25177
rect 31941 25143 31999 25149
rect 31941 25140 31953 25143
rect 30892 25112 31953 25140
rect 30892 25100 30898 25112
rect 31941 25109 31953 25112
rect 31987 25109 31999 25143
rect 31941 25103 31999 25109
rect 32677 25143 32735 25149
rect 32677 25109 32689 25143
rect 32723 25140 32735 25143
rect 69658 25140 69664 25152
rect 32723 25112 69664 25140
rect 32723 25109 32735 25112
rect 32677 25103 32735 25109
rect 69658 25100 69664 25112
rect 69716 25100 69722 25152
rect 1104 25050 78844 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 78844 25050
rect 1104 24976 78844 24998
rect 24394 24828 24400 24880
rect 24452 24868 24458 24880
rect 30834 24868 30840 24880
rect 24452 24840 30840 24868
rect 24452 24828 24458 24840
rect 30834 24828 30840 24840
rect 30892 24828 30898 24880
rect 41610 24871 41668 24877
rect 41610 24837 41622 24871
rect 41656 24837 41668 24871
rect 41610 24831 41668 24837
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24800 1731 24803
rect 2225 24803 2283 24809
rect 2225 24800 2237 24803
rect 1719 24772 2237 24800
rect 1719 24769 1731 24772
rect 1673 24763 1731 24769
rect 2225 24769 2237 24772
rect 2271 24800 2283 24803
rect 22278 24800 22284 24812
rect 2271 24772 22284 24800
rect 2271 24769 2283 24772
rect 2225 24763 2283 24769
rect 22278 24760 22284 24772
rect 22336 24760 22342 24812
rect 41233 24803 41291 24809
rect 41233 24769 41245 24803
rect 41279 24800 41291 24803
rect 41506 24800 41512 24812
rect 41279 24772 41512 24800
rect 41279 24769 41291 24772
rect 41233 24763 41291 24769
rect 41506 24760 41512 24772
rect 41564 24760 41570 24812
rect 1486 24664 1492 24676
rect 1447 24636 1492 24664
rect 1486 24624 1492 24636
rect 1544 24624 1550 24676
rect 40773 24667 40831 24673
rect 40773 24633 40785 24667
rect 40819 24664 40831 24667
rect 41616 24664 41644 24831
rect 77665 24803 77723 24809
rect 77665 24800 77677 24803
rect 77128 24772 77677 24800
rect 41690 24664 41696 24676
rect 40819 24636 41696 24664
rect 40819 24633 40831 24636
rect 40773 24627 40831 24633
rect 41690 24624 41696 24636
rect 41748 24624 41754 24676
rect 41785 24667 41843 24673
rect 41785 24633 41797 24667
rect 41831 24664 41843 24667
rect 60458 24664 60464 24676
rect 41831 24636 60464 24664
rect 41831 24633 41843 24636
rect 41785 24627 41843 24633
rect 60458 24624 60464 24636
rect 60516 24624 60522 24676
rect 41598 24596 41604 24608
rect 41559 24568 41604 24596
rect 41598 24556 41604 24568
rect 41656 24556 41662 24608
rect 69658 24556 69664 24608
rect 69716 24596 69722 24608
rect 77128 24605 77156 24772
rect 77665 24769 77677 24772
rect 77711 24769 77723 24803
rect 77665 24763 77723 24769
rect 77846 24664 77852 24676
rect 77807 24636 77852 24664
rect 77846 24624 77852 24636
rect 77904 24624 77910 24676
rect 77113 24599 77171 24605
rect 77113 24596 77125 24599
rect 69716 24568 77125 24596
rect 69716 24556 69722 24568
rect 77113 24565 77125 24568
rect 77159 24565 77171 24599
rect 77113 24559 77171 24565
rect 1104 24506 78844 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 78844 24506
rect 1104 24432 78844 24454
rect 22278 24392 22284 24404
rect 22239 24364 22284 24392
rect 22278 24352 22284 24364
rect 22336 24352 22342 24404
rect 41598 24352 41604 24404
rect 41656 24392 41662 24404
rect 41693 24395 41751 24401
rect 41693 24392 41705 24395
rect 41656 24364 41705 24392
rect 41656 24352 41662 24364
rect 41693 24361 41705 24364
rect 41739 24361 41751 24395
rect 41693 24355 41751 24361
rect 1673 24191 1731 24197
rect 1673 24157 1685 24191
rect 1719 24188 1731 24191
rect 2225 24191 2283 24197
rect 2225 24188 2237 24191
rect 1719 24160 2237 24188
rect 1719 24157 1731 24160
rect 1673 24151 1731 24157
rect 2225 24157 2237 24160
rect 2271 24188 2283 24191
rect 21818 24188 21824 24200
rect 2271 24160 21824 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 22465 24191 22523 24197
rect 22465 24157 22477 24191
rect 22511 24188 22523 24191
rect 32217 24191 32275 24197
rect 22511 24160 23060 24188
rect 22511 24157 22523 24160
rect 22465 24151 22523 24157
rect 23032 24129 23060 24160
rect 32217 24157 32229 24191
rect 32263 24188 32275 24191
rect 41969 24191 42027 24197
rect 32263 24160 41644 24188
rect 32263 24157 32275 24160
rect 32217 24151 32275 24157
rect 23017 24123 23075 24129
rect 23017 24089 23029 24123
rect 23063 24120 23075 24123
rect 23658 24120 23664 24132
rect 23063 24092 23664 24120
rect 23063 24089 23075 24092
rect 23017 24083 23075 24089
rect 23658 24080 23664 24092
rect 23716 24120 23722 24132
rect 31481 24123 31539 24129
rect 31481 24120 31493 24123
rect 23716 24092 31493 24120
rect 23716 24080 23722 24092
rect 31481 24089 31493 24092
rect 31527 24120 31539 24123
rect 32030 24120 32036 24132
rect 31527 24092 32036 24120
rect 31527 24089 31539 24092
rect 31481 24083 31539 24089
rect 32030 24080 32036 24092
rect 32088 24080 32094 24132
rect 40957 24123 41015 24129
rect 40957 24089 40969 24123
rect 41003 24120 41015 24123
rect 41506 24120 41512 24132
rect 41003 24092 41512 24120
rect 41003 24089 41015 24092
rect 40957 24083 41015 24089
rect 41506 24080 41512 24092
rect 41564 24080 41570 24132
rect 41616 24120 41644 24160
rect 41969 24157 41981 24191
rect 42015 24188 42027 24191
rect 77849 24191 77907 24197
rect 77849 24188 77861 24191
rect 42015 24160 55214 24188
rect 42015 24157 42027 24160
rect 41969 24151 42027 24157
rect 55186 24120 55214 24160
rect 77312 24160 77861 24188
rect 61194 24120 61200 24132
rect 41616 24092 45554 24120
rect 55186 24092 61200 24120
rect 1486 24052 1492 24064
rect 1447 24024 1492 24052
rect 1486 24012 1492 24024
rect 1544 24012 1550 24064
rect 41690 24052 41696 24064
rect 41651 24024 41696 24052
rect 41690 24012 41696 24024
rect 41748 24012 41754 24064
rect 45526 24052 45554 24092
rect 61194 24080 61200 24092
rect 61252 24080 61258 24132
rect 77312 24064 77340 24160
rect 77849 24157 77861 24160
rect 77895 24157 77907 24191
rect 77849 24151 77907 24157
rect 69658 24052 69664 24064
rect 45526 24024 69664 24052
rect 69658 24012 69664 24024
rect 69716 24012 69722 24064
rect 77294 24052 77300 24064
rect 77255 24024 77300 24052
rect 77294 24012 77300 24024
rect 77352 24012 77358 24064
rect 78030 24052 78036 24064
rect 77991 24024 78036 24052
rect 78030 24012 78036 24024
rect 78088 24012 78094 24064
rect 1104 23962 78844 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 78844 23962
rect 1104 23888 78844 23910
rect 21818 23848 21824 23860
rect 21779 23820 21824 23848
rect 21818 23808 21824 23820
rect 21876 23808 21882 23860
rect 30834 23848 30840 23860
rect 30795 23820 30840 23848
rect 30834 23808 30840 23820
rect 30892 23848 30898 23860
rect 31570 23848 31576 23860
rect 30892 23820 31576 23848
rect 30892 23808 30898 23820
rect 31570 23808 31576 23820
rect 31628 23808 31634 23860
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 22005 23715 22063 23721
rect 1719 23684 2268 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 2240 23585 2268 23684
rect 22005 23681 22017 23715
rect 22051 23712 22063 23715
rect 22554 23712 22560 23724
rect 22051 23684 22560 23712
rect 22051 23681 22063 23684
rect 22005 23675 22063 23681
rect 22554 23672 22560 23684
rect 22612 23672 22618 23724
rect 31386 23712 31392 23724
rect 31347 23684 31392 23712
rect 31386 23672 31392 23684
rect 31444 23672 31450 23724
rect 31478 23672 31484 23724
rect 31536 23712 31542 23724
rect 31573 23715 31631 23721
rect 31573 23712 31585 23715
rect 31536 23684 31585 23712
rect 31536 23672 31542 23684
rect 31573 23681 31585 23684
rect 31619 23681 31631 23715
rect 32214 23712 32220 23724
rect 32175 23684 32220 23712
rect 31573 23675 31631 23681
rect 32214 23672 32220 23684
rect 32272 23712 32278 23724
rect 32861 23715 32919 23721
rect 32861 23712 32873 23715
rect 32272 23684 32873 23712
rect 32272 23672 32278 23684
rect 32861 23681 32873 23684
rect 32907 23681 32919 23715
rect 32861 23675 32919 23681
rect 37182 23672 37188 23724
rect 37240 23712 37246 23724
rect 41690 23712 41696 23724
rect 37240 23684 41696 23712
rect 37240 23672 37246 23684
rect 41690 23672 41696 23684
rect 41748 23672 41754 23724
rect 77110 23672 77116 23724
rect 77168 23712 77174 23724
rect 77665 23715 77723 23721
rect 77665 23712 77677 23715
rect 77168 23684 77677 23712
rect 77168 23672 77174 23684
rect 77665 23681 77677 23684
rect 77711 23681 77723 23715
rect 77665 23675 77723 23681
rect 32401 23647 32459 23653
rect 32401 23613 32413 23647
rect 32447 23644 32459 23647
rect 77294 23644 77300 23656
rect 32447 23616 77300 23644
rect 32447 23613 32459 23616
rect 32401 23607 32459 23613
rect 77294 23604 77300 23616
rect 77352 23604 77358 23656
rect 2225 23579 2283 23585
rect 2225 23545 2237 23579
rect 2271 23576 2283 23579
rect 19702 23576 19708 23588
rect 2271 23548 19708 23576
rect 2271 23545 2283 23548
rect 2225 23539 2283 23545
rect 19702 23536 19708 23548
rect 19760 23536 19766 23588
rect 31573 23579 31631 23585
rect 31573 23545 31585 23579
rect 31619 23576 31631 23579
rect 41598 23576 41604 23588
rect 31619 23548 41604 23576
rect 31619 23545 31631 23548
rect 31573 23539 31631 23545
rect 41598 23536 41604 23548
rect 41656 23536 41662 23588
rect 1486 23508 1492 23520
rect 1447 23480 1492 23508
rect 1486 23468 1492 23480
rect 1544 23468 1550 23520
rect 22554 23508 22560 23520
rect 22515 23480 22560 23508
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 41233 23511 41291 23517
rect 41233 23477 41245 23511
rect 41279 23508 41291 23511
rect 41506 23508 41512 23520
rect 41279 23480 41512 23508
rect 41279 23477 41291 23480
rect 41233 23471 41291 23477
rect 41506 23468 41512 23480
rect 41564 23468 41570 23520
rect 77110 23508 77116 23520
rect 77071 23480 77116 23508
rect 77110 23468 77116 23480
rect 77168 23468 77174 23520
rect 77846 23508 77852 23520
rect 77807 23480 77852 23508
rect 77846 23468 77852 23480
rect 77904 23468 77910 23520
rect 1104 23418 78844 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 78844 23418
rect 1104 23344 78844 23366
rect 19702 23304 19708 23316
rect 19663 23276 19708 23304
rect 19702 23264 19708 23276
rect 19760 23264 19766 23316
rect 24946 23264 24952 23316
rect 25004 23304 25010 23316
rect 30282 23304 30288 23316
rect 25004 23276 30288 23304
rect 25004 23264 25010 23276
rect 30282 23264 30288 23276
rect 30340 23264 30346 23316
rect 31389 23307 31447 23313
rect 31389 23273 31401 23307
rect 31435 23304 31447 23307
rect 31478 23304 31484 23316
rect 31435 23276 31484 23304
rect 31435 23273 31447 23276
rect 31389 23267 31447 23273
rect 31478 23264 31484 23276
rect 31536 23264 31542 23316
rect 31570 23264 31576 23316
rect 31628 23304 31634 23316
rect 31628 23276 31673 23304
rect 31628 23264 31634 23276
rect 27985 23171 28043 23177
rect 27985 23137 27997 23171
rect 28031 23168 28043 23171
rect 77110 23168 77116 23180
rect 28031 23140 77116 23168
rect 28031 23137 28043 23140
rect 27985 23131 28043 23137
rect 77110 23128 77116 23140
rect 77168 23128 77174 23180
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23069 1731 23103
rect 1673 23063 1731 23069
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23100 19947 23103
rect 19935 23072 20484 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 1688 23032 1716 23063
rect 2225 23035 2283 23041
rect 2225 23032 2237 23035
rect 1688 23004 2237 23032
rect 2225 23001 2237 23004
rect 2271 23032 2283 23035
rect 19978 23032 19984 23044
rect 2271 23004 19984 23032
rect 2271 23001 2283 23004
rect 2225 22995 2283 23001
rect 19978 22992 19984 23004
rect 20036 22992 20042 23044
rect 1486 22964 1492 22976
rect 1447 22936 1492 22964
rect 1486 22924 1492 22936
rect 1544 22924 1550 22976
rect 20456 22973 20484 23072
rect 22554 23060 22560 23112
rect 22612 23100 22618 23112
rect 22922 23100 22928 23112
rect 22612 23072 22928 23100
rect 22612 23060 22618 23072
rect 22922 23060 22928 23072
rect 22980 23100 22986 23112
rect 31573 23103 31631 23109
rect 22980 23072 30972 23100
rect 22980 23060 22986 23072
rect 30944 23041 30972 23072
rect 31573 23069 31585 23103
rect 31619 23100 31631 23103
rect 31662 23100 31668 23112
rect 31619 23072 31668 23100
rect 31619 23069 31631 23072
rect 31573 23063 31631 23069
rect 31662 23060 31668 23072
rect 31720 23060 31726 23112
rect 31941 23103 31999 23109
rect 31941 23069 31953 23103
rect 31987 23069 31999 23103
rect 31941 23063 31999 23069
rect 27801 23035 27859 23041
rect 27801 23001 27813 23035
rect 27847 23001 27859 23035
rect 27801 22995 27859 23001
rect 30929 23035 30987 23041
rect 30929 23001 30941 23035
rect 30975 23032 30987 23035
rect 31956 23032 31984 23063
rect 32030 23060 32036 23112
rect 32088 23100 32094 23112
rect 77849 23103 77907 23109
rect 77849 23100 77861 23103
rect 32088 23072 32133 23100
rect 77312 23072 77861 23100
rect 32088 23060 32094 23072
rect 32214 23032 32220 23044
rect 30975 23004 32220 23032
rect 30975 23001 30987 23004
rect 30929 22995 30987 23001
rect 20441 22967 20499 22973
rect 20441 22933 20453 22967
rect 20487 22964 20499 22967
rect 27154 22964 27160 22976
rect 20487 22936 27160 22964
rect 20487 22933 20499 22936
rect 20441 22927 20499 22933
rect 27154 22924 27160 22936
rect 27212 22964 27218 22976
rect 27816 22964 27844 22995
rect 32214 22992 32220 23004
rect 32272 22992 32278 23044
rect 77312 22976 77340 23072
rect 77849 23069 77861 23072
rect 77895 23069 77907 23103
rect 77849 23063 77907 23069
rect 27212 22936 27844 22964
rect 27212 22924 27218 22936
rect 30282 22924 30288 22976
rect 30340 22964 30346 22976
rect 30377 22967 30435 22973
rect 30377 22964 30389 22967
rect 30340 22936 30389 22964
rect 30340 22924 30346 22936
rect 30377 22933 30389 22936
rect 30423 22964 30435 22967
rect 31662 22964 31668 22976
rect 30423 22936 31668 22964
rect 30423 22933 30435 22936
rect 30377 22927 30435 22933
rect 31662 22924 31668 22936
rect 31720 22924 31726 22976
rect 77294 22964 77300 22976
rect 77255 22936 77300 22964
rect 77294 22924 77300 22936
rect 77352 22924 77358 22976
rect 78030 22964 78036 22976
rect 77991 22936 78036 22964
rect 78030 22924 78036 22936
rect 78088 22924 78094 22976
rect 1104 22874 78844 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 78844 22874
rect 1104 22800 78844 22822
rect 19978 22760 19984 22772
rect 19939 22732 19984 22760
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 31113 22763 31171 22769
rect 31113 22729 31125 22763
rect 31159 22760 31171 22763
rect 32030 22760 32036 22772
rect 31159 22732 32036 22760
rect 31159 22729 31171 22732
rect 31113 22723 31171 22729
rect 32030 22720 32036 22732
rect 32088 22720 32094 22772
rect 20165 22627 20223 22633
rect 20165 22593 20177 22627
rect 20211 22624 20223 22627
rect 27801 22627 27859 22633
rect 27801 22624 27813 22627
rect 20211 22596 20760 22624
rect 20211 22593 20223 22596
rect 20165 22587 20223 22593
rect 20732 22429 20760 22596
rect 27172 22596 27813 22624
rect 20717 22423 20775 22429
rect 20717 22389 20729 22423
rect 20763 22420 20775 22423
rect 26970 22420 26976 22432
rect 20763 22392 26976 22420
rect 20763 22389 20775 22392
rect 20717 22383 20775 22389
rect 26970 22380 26976 22392
rect 27028 22420 27034 22432
rect 27172 22429 27200 22596
rect 27801 22593 27813 22596
rect 27847 22593 27859 22627
rect 27801 22587 27859 22593
rect 27985 22491 28043 22497
rect 27985 22457 27997 22491
rect 28031 22488 28043 22491
rect 77294 22488 77300 22500
rect 28031 22460 77300 22488
rect 28031 22457 28043 22460
rect 27985 22451 28043 22457
rect 77294 22448 77300 22460
rect 77352 22448 77358 22500
rect 27157 22423 27215 22429
rect 27157 22420 27169 22423
rect 27028 22392 27169 22420
rect 27028 22380 27034 22392
rect 27157 22389 27169 22392
rect 27203 22389 27215 22423
rect 27157 22383 27215 22389
rect 1104 22330 78844 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 78844 22330
rect 1104 22256 78844 22278
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 22012 1731 22015
rect 19058 22012 19064 22024
rect 1719 21984 19064 22012
rect 1719 21981 1731 21984
rect 1673 21975 1731 21981
rect 19058 21972 19064 21984
rect 19116 21972 19122 22024
rect 77849 22015 77907 22021
rect 77849 22012 77861 22015
rect 77312 21984 77861 22012
rect 27338 21904 27344 21956
rect 27396 21944 27402 21956
rect 27433 21947 27491 21953
rect 27433 21944 27445 21947
rect 27396 21916 27445 21944
rect 27396 21904 27402 21916
rect 27433 21913 27445 21916
rect 27479 21944 27491 21947
rect 27985 21947 28043 21953
rect 27985 21944 27997 21947
rect 27479 21916 27997 21944
rect 27479 21913 27491 21916
rect 27433 21907 27491 21913
rect 27985 21913 27997 21916
rect 28031 21913 28043 21947
rect 27985 21907 28043 21913
rect 1486 21876 1492 21888
rect 1447 21848 1492 21876
rect 1486 21836 1492 21848
rect 1544 21836 1550 21888
rect 77312 21885 77340 21984
rect 77849 21981 77861 21984
rect 77895 21981 77907 22015
rect 77849 21975 77907 21981
rect 28077 21879 28135 21885
rect 28077 21845 28089 21879
rect 28123 21876 28135 21879
rect 77297 21879 77355 21885
rect 77297 21876 77309 21879
rect 28123 21848 77309 21876
rect 28123 21845 28135 21848
rect 28077 21839 28135 21845
rect 77297 21845 77309 21848
rect 77343 21845 77355 21879
rect 78030 21876 78036 21888
rect 77991 21848 78036 21876
rect 77297 21839 77355 21845
rect 78030 21836 78036 21848
rect 78088 21836 78094 21888
rect 1104 21786 78844 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 78844 21786
rect 1104 21712 78844 21734
rect 19058 21672 19064 21684
rect 19019 21644 19064 21672
rect 19058 21632 19064 21644
rect 19116 21632 19122 21684
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 17862 21536 17868 21548
rect 1719 21508 17868 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 17862 21496 17868 21508
rect 17920 21496 17926 21548
rect 19245 21539 19303 21545
rect 19245 21505 19257 21539
rect 19291 21536 19303 21539
rect 77665 21539 77723 21545
rect 77665 21536 77677 21539
rect 19291 21508 19840 21536
rect 19291 21505 19303 21508
rect 19245 21499 19303 21505
rect 1486 21332 1492 21344
rect 1447 21304 1492 21332
rect 1486 21292 1492 21304
rect 1544 21292 1550 21344
rect 19812 21341 19840 21508
rect 77128 21508 77677 21536
rect 77128 21344 77156 21508
rect 77665 21505 77677 21508
rect 77711 21505 77723 21539
rect 77665 21499 77723 21505
rect 19797 21335 19855 21341
rect 19797 21301 19809 21335
rect 19843 21332 19855 21335
rect 20346 21332 20352 21344
rect 19843 21304 20352 21332
rect 19843 21301 19855 21304
rect 19797 21295 19855 21301
rect 20346 21292 20352 21304
rect 20404 21292 20410 21344
rect 77110 21332 77116 21344
rect 77071 21304 77116 21332
rect 77110 21292 77116 21304
rect 77168 21292 77174 21344
rect 77846 21332 77852 21344
rect 77807 21304 77852 21332
rect 77846 21292 77852 21304
rect 77904 21292 77910 21344
rect 1104 21242 78844 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 78844 21242
rect 1104 21168 78844 21190
rect 17862 21128 17868 21140
rect 17823 21100 17868 21128
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 17954 20924 17960 20936
rect 1719 20896 17960 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20924 18107 20927
rect 18601 20927 18659 20933
rect 18601 20924 18613 20927
rect 18095 20896 18613 20924
rect 18095 20893 18107 20896
rect 18049 20887 18107 20893
rect 18601 20893 18613 20896
rect 18647 20924 18659 20927
rect 19426 20924 19432 20936
rect 18647 20896 19432 20924
rect 18647 20893 18659 20896
rect 18601 20887 18659 20893
rect 19426 20884 19432 20896
rect 19484 20924 19490 20936
rect 19484 20896 26234 20924
rect 19484 20884 19490 20896
rect 1486 20788 1492 20800
rect 1447 20760 1492 20788
rect 1486 20748 1492 20760
rect 1544 20748 1550 20800
rect 26206 20788 26234 20896
rect 32398 20884 32404 20936
rect 32456 20924 32462 20936
rect 77297 20927 77355 20933
rect 77297 20924 77309 20927
rect 32456 20896 77309 20924
rect 32456 20884 32462 20896
rect 77297 20893 77309 20896
rect 77343 20924 77355 20927
rect 77849 20927 77907 20933
rect 77849 20924 77861 20927
rect 77343 20896 77861 20924
rect 77343 20893 77355 20896
rect 77297 20887 77355 20893
rect 77849 20893 77861 20896
rect 77895 20893 77907 20927
rect 77849 20887 77907 20893
rect 27801 20859 27859 20865
rect 27801 20825 27813 20859
rect 27847 20825 27859 20859
rect 27801 20819 27859 20825
rect 27062 20788 27068 20800
rect 26206 20760 27068 20788
rect 27062 20748 27068 20760
rect 27120 20788 27126 20800
rect 27157 20791 27215 20797
rect 27157 20788 27169 20791
rect 27120 20760 27169 20788
rect 27120 20748 27126 20760
rect 27157 20757 27169 20760
rect 27203 20788 27215 20791
rect 27816 20788 27844 20819
rect 27203 20760 27844 20788
rect 27893 20791 27951 20797
rect 27203 20757 27215 20760
rect 27157 20751 27215 20757
rect 27893 20757 27905 20791
rect 27939 20788 27951 20791
rect 77110 20788 77116 20800
rect 27939 20760 77116 20788
rect 27939 20757 27951 20760
rect 27893 20751 27951 20757
rect 77110 20748 77116 20760
rect 77168 20748 77174 20800
rect 78030 20788 78036 20800
rect 77991 20760 78036 20788
rect 78030 20748 78036 20760
rect 78088 20748 78094 20800
rect 1104 20698 78844 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 78844 20698
rect 1104 20624 78844 20646
rect 17954 20544 17960 20596
rect 18012 20584 18018 20596
rect 18509 20587 18567 20593
rect 18509 20584 18521 20587
rect 18012 20556 18521 20584
rect 18012 20544 18018 20556
rect 18509 20553 18521 20556
rect 18555 20553 18567 20587
rect 18509 20547 18567 20553
rect 32398 20516 32404 20528
rect 32359 20488 32404 20516
rect 32398 20476 32404 20488
rect 32456 20476 32462 20528
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 17034 20448 17040 20460
rect 1719 20420 17040 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20448 18751 20451
rect 18739 20420 19288 20448
rect 18739 20417 18751 20420
rect 18693 20411 18751 20417
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 19260 20253 19288 20420
rect 31478 20408 31484 20460
rect 31536 20448 31542 20460
rect 32217 20451 32275 20457
rect 32217 20448 32229 20451
rect 31536 20420 32229 20448
rect 31536 20408 31542 20420
rect 32217 20417 32229 20420
rect 32263 20417 32275 20451
rect 77665 20451 77723 20457
rect 77665 20448 77677 20451
rect 32217 20411 32275 20417
rect 77128 20420 77677 20448
rect 19245 20247 19303 20253
rect 19245 20213 19257 20247
rect 19291 20244 19303 20247
rect 19334 20244 19340 20256
rect 19291 20216 19340 20244
rect 19291 20213 19303 20216
rect 19245 20207 19303 20213
rect 19334 20204 19340 20216
rect 19392 20204 19398 20256
rect 31478 20244 31484 20256
rect 31439 20216 31484 20244
rect 31478 20204 31484 20216
rect 31536 20204 31542 20256
rect 68002 20204 68008 20256
rect 68060 20244 68066 20256
rect 77128 20253 77156 20420
rect 77665 20417 77677 20420
rect 77711 20417 77723 20451
rect 77665 20411 77723 20417
rect 77113 20247 77171 20253
rect 77113 20244 77125 20247
rect 68060 20216 77125 20244
rect 68060 20204 68066 20216
rect 77113 20213 77125 20216
rect 77159 20213 77171 20247
rect 77846 20244 77852 20256
rect 77807 20216 77852 20244
rect 77113 20207 77171 20213
rect 77846 20204 77852 20216
rect 77904 20204 77910 20256
rect 1104 20154 78844 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 78844 20154
rect 1104 20080 78844 20102
rect 17034 20040 17040 20052
rect 16995 20012 17040 20040
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 17221 19839 17279 19845
rect 17221 19805 17233 19839
rect 17267 19836 17279 19839
rect 17267 19808 17816 19836
rect 17267 19805 17279 19808
rect 17221 19799 17279 19805
rect 17788 19709 17816 19808
rect 31573 19771 31631 19777
rect 31573 19737 31585 19771
rect 31619 19737 31631 19771
rect 31573 19731 31631 19737
rect 31757 19771 31815 19777
rect 31757 19737 31769 19771
rect 31803 19768 31815 19771
rect 31803 19740 35894 19768
rect 31803 19737 31815 19740
rect 31757 19731 31815 19737
rect 17773 19703 17831 19709
rect 17773 19669 17785 19703
rect 17819 19700 17831 19703
rect 17954 19700 17960 19712
rect 17819 19672 17960 19700
rect 17819 19669 17831 19672
rect 17773 19663 17831 19669
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 30926 19700 30932 19712
rect 30887 19672 30932 19700
rect 30926 19660 30932 19672
rect 30984 19700 30990 19712
rect 31588 19700 31616 19731
rect 30984 19672 31616 19700
rect 35866 19700 35894 19740
rect 68002 19700 68008 19712
rect 35866 19672 68008 19700
rect 30984 19660 30990 19672
rect 68002 19660 68008 19672
rect 68060 19660 68066 19712
rect 1104 19610 78844 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 78844 19610
rect 1104 19536 78844 19558
rect 16669 19499 16727 19505
rect 16669 19496 16681 19499
rect 6886 19468 16681 19496
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 6886 19360 6914 19468
rect 16669 19465 16681 19468
rect 16715 19465 16727 19499
rect 77846 19496 77852 19508
rect 77807 19468 77852 19496
rect 16669 19459 16727 19465
rect 77846 19456 77852 19468
rect 77904 19456 77910 19508
rect 1719 19332 6914 19360
rect 16853 19363 16911 19369
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 16853 19329 16865 19363
rect 16899 19360 16911 19363
rect 16899 19332 17448 19360
rect 16899 19329 16911 19332
rect 16853 19323 16911 19329
rect 1486 19224 1492 19236
rect 1447 19196 1492 19224
rect 1486 19184 1492 19196
rect 1544 19184 1550 19236
rect 17420 19165 17448 19332
rect 17954 19320 17960 19372
rect 18012 19360 18018 19372
rect 18506 19360 18512 19372
rect 18012 19332 18512 19360
rect 18012 19320 18018 19332
rect 18506 19320 18512 19332
rect 18564 19360 18570 19372
rect 30561 19363 30619 19369
rect 30561 19360 30573 19363
rect 18564 19332 30573 19360
rect 18564 19320 18570 19332
rect 30561 19329 30573 19332
rect 30607 19360 30619 19363
rect 30926 19360 30932 19372
rect 30607 19332 30932 19360
rect 30607 19329 30619 19332
rect 30561 19323 30619 19329
rect 30926 19320 30932 19332
rect 30984 19320 30990 19372
rect 31754 19320 31760 19372
rect 31812 19360 31818 19372
rect 32217 19363 32275 19369
rect 32217 19360 32229 19363
rect 31812 19332 32229 19360
rect 31812 19320 31818 19332
rect 32217 19329 32229 19332
rect 32263 19329 32275 19363
rect 32217 19323 32275 19329
rect 77665 19363 77723 19369
rect 77665 19329 77677 19363
rect 77711 19329 77723 19363
rect 77665 19323 77723 19329
rect 77680 19292 77708 19323
rect 77128 19264 77708 19292
rect 17405 19159 17463 19165
rect 17405 19125 17417 19159
rect 17451 19156 17463 19159
rect 17770 19156 17776 19168
rect 17451 19128 17776 19156
rect 17451 19125 17463 19128
rect 17405 19119 17463 19125
rect 17770 19116 17776 19128
rect 17828 19156 17834 19168
rect 31481 19159 31539 19165
rect 31481 19156 31493 19159
rect 17828 19128 31493 19156
rect 17828 19116 17834 19128
rect 31481 19125 31493 19128
rect 31527 19156 31539 19159
rect 31754 19156 31760 19168
rect 31527 19128 31760 19156
rect 31527 19125 31539 19128
rect 31481 19119 31539 19125
rect 31754 19116 31760 19128
rect 31812 19116 31818 19168
rect 77128 19165 77156 19264
rect 32309 19159 32367 19165
rect 32309 19125 32321 19159
rect 32355 19156 32367 19159
rect 77113 19159 77171 19165
rect 77113 19156 77125 19159
rect 32355 19128 77125 19156
rect 32355 19125 32367 19128
rect 32309 19119 32367 19125
rect 77113 19125 77125 19128
rect 77159 19125 77171 19159
rect 77113 19119 77171 19125
rect 1104 19066 78844 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 78844 19066
rect 1104 18992 78844 19014
rect 31113 18955 31171 18961
rect 31113 18952 31125 18955
rect 30576 18924 31125 18952
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 16301 18751 16359 18757
rect 1719 18720 6914 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 6886 18612 6914 18720
rect 16301 18717 16313 18751
rect 16347 18748 16359 18751
rect 16347 18720 16574 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 6886 18584 16129 18612
rect 16117 18581 16129 18584
rect 16163 18581 16175 18615
rect 16546 18612 16574 18720
rect 19334 18640 19340 18692
rect 19392 18680 19398 18692
rect 30009 18683 30067 18689
rect 30009 18680 30021 18683
rect 19392 18652 30021 18680
rect 19392 18640 19398 18652
rect 30009 18649 30021 18652
rect 30055 18680 30067 18683
rect 30466 18680 30472 18692
rect 30055 18652 30472 18680
rect 30055 18649 30067 18652
rect 30009 18643 30067 18649
rect 30466 18640 30472 18652
rect 30524 18640 30530 18692
rect 30576 18680 30604 18924
rect 31113 18921 31125 18924
rect 31159 18921 31171 18955
rect 31113 18915 31171 18921
rect 31386 18912 31392 18964
rect 31444 18952 31450 18964
rect 31573 18955 31631 18961
rect 31573 18952 31585 18955
rect 31444 18924 31585 18952
rect 31444 18912 31450 18924
rect 31573 18921 31585 18924
rect 31619 18921 31631 18955
rect 31573 18915 31631 18921
rect 30650 18776 30656 18828
rect 30708 18816 30714 18828
rect 31205 18819 31263 18825
rect 31205 18816 31217 18819
rect 30708 18788 31217 18816
rect 30708 18776 30714 18788
rect 31205 18785 31217 18788
rect 31251 18816 31263 18819
rect 31478 18816 31484 18828
rect 31251 18788 31484 18816
rect 31251 18785 31263 18788
rect 31205 18779 31263 18785
rect 31478 18776 31484 18788
rect 31536 18776 31542 18828
rect 30926 18708 30932 18760
rect 30984 18748 30990 18760
rect 31113 18751 31171 18757
rect 31113 18748 31125 18751
rect 30984 18720 31125 18748
rect 30984 18708 30990 18720
rect 31113 18717 31125 18720
rect 31159 18717 31171 18751
rect 31113 18711 31171 18717
rect 31389 18751 31447 18757
rect 31389 18717 31401 18751
rect 31435 18748 31447 18751
rect 31754 18748 31760 18760
rect 31435 18720 31760 18748
rect 31435 18717 31447 18720
rect 31389 18711 31447 18717
rect 31754 18708 31760 18720
rect 31812 18708 31818 18760
rect 77849 18751 77907 18757
rect 77849 18748 77861 18751
rect 77312 18720 77861 18748
rect 32125 18683 32183 18689
rect 32125 18680 32137 18683
rect 30576 18652 32137 18680
rect 30576 18624 30604 18652
rect 32125 18649 32137 18652
rect 32171 18649 32183 18683
rect 32125 18643 32183 18649
rect 16850 18612 16856 18624
rect 16546 18584 16856 18612
rect 16117 18575 16175 18581
rect 16850 18572 16856 18584
rect 16908 18572 16914 18624
rect 26326 18612 26332 18624
rect 26287 18584 26332 18612
rect 26326 18572 26332 18584
rect 26384 18572 26390 18624
rect 26973 18615 27031 18621
rect 26973 18581 26985 18615
rect 27019 18612 27031 18615
rect 27062 18612 27068 18624
rect 27019 18584 27068 18612
rect 27019 18581 27031 18584
rect 26973 18575 27031 18581
rect 27062 18572 27068 18584
rect 27120 18572 27126 18624
rect 30558 18612 30564 18624
rect 30519 18584 30564 18612
rect 30558 18572 30564 18584
rect 30616 18572 30622 18624
rect 77312 18621 77340 18720
rect 77849 18717 77861 18720
rect 77895 18717 77907 18751
rect 77849 18711 77907 18717
rect 32217 18615 32275 18621
rect 32217 18581 32229 18615
rect 32263 18612 32275 18615
rect 77297 18615 77355 18621
rect 77297 18612 77309 18615
rect 32263 18584 77309 18612
rect 32263 18581 32275 18584
rect 32217 18575 32275 18581
rect 77297 18581 77309 18584
rect 77343 18581 77355 18615
rect 78030 18612 78036 18624
rect 77991 18584 78036 18612
rect 77297 18575 77355 18581
rect 78030 18572 78036 18584
rect 78088 18572 78094 18624
rect 1104 18522 78844 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 78844 18522
rect 1104 18448 78844 18470
rect 16850 18368 16856 18420
rect 16908 18408 16914 18420
rect 17034 18408 17040 18420
rect 16908 18380 17040 18408
rect 16908 18368 16914 18380
rect 17034 18368 17040 18380
rect 17092 18408 17098 18420
rect 30558 18408 30564 18420
rect 17092 18380 30564 18408
rect 17092 18368 17098 18380
rect 30558 18368 30564 18380
rect 30616 18408 30622 18420
rect 32125 18411 32183 18417
rect 32125 18408 32137 18411
rect 30616 18380 32137 18408
rect 30616 18368 30622 18380
rect 32125 18377 32137 18380
rect 32171 18377 32183 18411
rect 32125 18371 32183 18377
rect 26421 18343 26479 18349
rect 26421 18340 26433 18343
rect 26206 18312 26433 18340
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 12342 18272 12348 18284
rect 1719 18244 12348 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 20346 18028 20352 18080
rect 20404 18068 20410 18080
rect 26206 18068 26234 18312
rect 26421 18309 26433 18312
rect 26467 18340 26479 18343
rect 30837 18343 30895 18349
rect 26467 18312 27384 18340
rect 26467 18309 26479 18312
rect 26421 18303 26479 18309
rect 27356 18284 27384 18312
rect 30837 18309 30849 18343
rect 30883 18340 30895 18343
rect 31754 18340 31760 18352
rect 30883 18312 31760 18340
rect 30883 18309 30895 18312
rect 30837 18303 30895 18309
rect 31754 18300 31760 18312
rect 31812 18300 31818 18352
rect 26510 18232 26516 18284
rect 26568 18272 26574 18284
rect 26970 18272 26976 18284
rect 26568 18244 26976 18272
rect 26568 18232 26574 18244
rect 26970 18232 26976 18244
rect 27028 18272 27034 18284
rect 27065 18275 27123 18281
rect 27065 18272 27077 18275
rect 27028 18244 27077 18272
rect 27028 18232 27034 18244
rect 27065 18241 27077 18244
rect 27111 18241 27123 18275
rect 27338 18272 27344 18284
rect 27299 18244 27344 18272
rect 27065 18235 27123 18241
rect 27338 18232 27344 18244
rect 27396 18232 27402 18284
rect 77110 18232 77116 18284
rect 77168 18272 77174 18284
rect 77665 18275 77723 18281
rect 77665 18272 77677 18275
rect 77168 18244 77677 18272
rect 77168 18232 77174 18244
rect 77665 18241 77677 18244
rect 77711 18241 77723 18275
rect 77665 18235 77723 18241
rect 27154 18204 27160 18216
rect 27067 18176 27160 18204
rect 27154 18164 27160 18176
rect 27212 18164 27218 18216
rect 26326 18096 26332 18148
rect 26384 18136 26390 18148
rect 27172 18136 27200 18164
rect 26384 18108 27200 18136
rect 26384 18096 26390 18108
rect 27062 18068 27068 18080
rect 20404 18040 26234 18068
rect 27023 18040 27068 18068
rect 20404 18028 20410 18040
rect 27062 18028 27068 18040
rect 27120 18028 27126 18080
rect 27525 18071 27583 18077
rect 27525 18037 27537 18071
rect 27571 18068 27583 18071
rect 27706 18068 27712 18080
rect 27571 18040 27712 18068
rect 27571 18037 27583 18040
rect 27525 18031 27583 18037
rect 27706 18028 27712 18040
rect 27764 18028 27770 18080
rect 77110 18068 77116 18080
rect 77071 18040 77116 18068
rect 77110 18028 77116 18040
rect 77168 18028 77174 18080
rect 77846 18068 77852 18080
rect 77807 18040 77852 18068
rect 77846 18028 77852 18040
rect 77904 18028 77910 18080
rect 1104 17978 78844 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 78844 17978
rect 1104 17904 78844 17926
rect 12342 17824 12348 17876
rect 12400 17864 12406 17876
rect 14829 17867 14887 17873
rect 14829 17864 14841 17867
rect 12400 17836 14841 17864
rect 12400 17824 12406 17836
rect 14829 17833 14841 17836
rect 14875 17833 14887 17867
rect 14829 17827 14887 17833
rect 27706 17728 27712 17740
rect 27667 17700 27712 17728
rect 27706 17688 27712 17700
rect 27764 17688 27770 17740
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 14458 17660 14464 17672
rect 1719 17632 14464 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 14458 17620 14464 17632
rect 14516 17620 14522 17672
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17660 15071 17663
rect 27338 17660 27344 17672
rect 15059 17632 15608 17660
rect 27299 17632 27344 17660
rect 15059 17629 15071 17632
rect 15013 17623 15071 17629
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 15580 17533 15608 17632
rect 27338 17620 27344 17632
rect 27396 17620 27402 17672
rect 27522 17660 27528 17672
rect 27483 17632 27528 17660
rect 27522 17620 27528 17632
rect 27580 17620 27586 17672
rect 77849 17663 77907 17669
rect 77849 17660 77861 17663
rect 77312 17632 77861 17660
rect 15565 17527 15623 17533
rect 15565 17493 15577 17527
rect 15611 17524 15623 17527
rect 15930 17524 15936 17536
rect 15611 17496 15936 17524
rect 15611 17493 15623 17496
rect 15565 17487 15623 17493
rect 15930 17484 15936 17496
rect 15988 17524 15994 17536
rect 26418 17524 26424 17536
rect 15988 17496 26424 17524
rect 15988 17484 15994 17496
rect 26418 17484 26424 17496
rect 26476 17484 26482 17536
rect 26510 17484 26516 17536
rect 26568 17524 26574 17536
rect 27801 17527 27859 17533
rect 26568 17496 26613 17524
rect 26568 17484 26574 17496
rect 27801 17493 27813 17527
rect 27847 17524 27859 17527
rect 37182 17524 37188 17536
rect 27847 17496 37188 17524
rect 27847 17493 27859 17496
rect 27801 17487 27859 17493
rect 37182 17484 37188 17496
rect 37240 17484 37246 17536
rect 77018 17484 77024 17536
rect 77076 17524 77082 17536
rect 77312 17533 77340 17632
rect 77849 17629 77861 17632
rect 77895 17629 77907 17663
rect 77849 17623 77907 17629
rect 77297 17527 77355 17533
rect 77297 17524 77309 17527
rect 77076 17496 77309 17524
rect 77076 17484 77082 17496
rect 77297 17493 77309 17496
rect 77343 17493 77355 17527
rect 78030 17524 78036 17536
rect 77991 17496 78036 17524
rect 77297 17487 77355 17493
rect 78030 17484 78036 17496
rect 78088 17484 78094 17536
rect 1104 17434 78844 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 78844 17434
rect 1104 17360 78844 17382
rect 14458 17320 14464 17332
rect 14419 17292 14464 17320
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 14645 17187 14703 17193
rect 14645 17153 14657 17187
rect 14691 17184 14703 17187
rect 26418 17184 26424 17196
rect 14691 17156 15240 17184
rect 26331 17156 26424 17184
rect 14691 17153 14703 17156
rect 14645 17147 14703 17153
rect 15102 16940 15108 16992
rect 15160 16980 15166 16992
rect 15212 16989 15240 17156
rect 26418 17144 26424 17156
rect 26476 17184 26482 17196
rect 27525 17187 27583 17193
rect 27525 17184 27537 17187
rect 26476 17156 27537 17184
rect 26476 17144 26482 17156
rect 27525 17153 27537 17156
rect 27571 17153 27583 17187
rect 27525 17147 27583 17153
rect 27709 17051 27767 17057
rect 27709 17017 27721 17051
rect 27755 17048 27767 17051
rect 27755 17020 35894 17048
rect 27755 17017 27767 17020
rect 27709 17011 27767 17017
rect 15197 16983 15255 16989
rect 15197 16980 15209 16983
rect 15160 16952 15209 16980
rect 15160 16940 15166 16952
rect 15197 16949 15209 16952
rect 15243 16980 15255 16983
rect 26234 16980 26240 16992
rect 15243 16952 26240 16980
rect 15243 16949 15255 16952
rect 15197 16943 15255 16949
rect 26234 16940 26240 16952
rect 26292 16940 26298 16992
rect 28166 16980 28172 16992
rect 28127 16952 28172 16980
rect 28166 16940 28172 16952
rect 28224 16940 28230 16992
rect 35866 16980 35894 17020
rect 77110 16980 77116 16992
rect 35866 16952 77116 16980
rect 77110 16940 77116 16952
rect 77168 16940 77174 16992
rect 1104 16890 78844 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 78844 16890
rect 1104 16816 78844 16838
rect 26237 16779 26295 16785
rect 26237 16745 26249 16779
rect 26283 16776 26295 16779
rect 26418 16776 26424 16788
rect 26283 16748 26424 16776
rect 26283 16745 26295 16748
rect 26237 16739 26295 16745
rect 26418 16736 26424 16748
rect 26476 16736 26482 16788
rect 28169 16779 28227 16785
rect 28169 16745 28181 16779
rect 28215 16776 28227 16779
rect 28215 16748 35894 16776
rect 28215 16745 28227 16748
rect 28169 16739 28227 16745
rect 27525 16711 27583 16717
rect 27525 16677 27537 16711
rect 27571 16708 27583 16711
rect 35866 16708 35894 16748
rect 77297 16711 77355 16717
rect 77297 16708 77309 16711
rect 27571 16680 31708 16708
rect 35866 16680 77309 16708
rect 27571 16677 27583 16680
rect 27525 16671 27583 16677
rect 31680 16640 31708 16680
rect 77297 16677 77309 16680
rect 77343 16708 77355 16711
rect 77343 16680 77892 16708
rect 77343 16677 77355 16680
rect 77297 16671 77355 16677
rect 77018 16640 77024 16652
rect 31680 16612 77024 16640
rect 77018 16600 77024 16612
rect 77076 16600 77082 16652
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 12710 16572 12716 16584
rect 1719 16544 12716 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 12710 16532 12716 16544
rect 12768 16532 12774 16584
rect 28077 16575 28135 16581
rect 28077 16541 28089 16575
rect 28123 16572 28135 16575
rect 28166 16572 28172 16584
rect 28123 16544 28172 16572
rect 28123 16541 28135 16544
rect 28077 16535 28135 16541
rect 28166 16532 28172 16544
rect 28224 16532 28230 16584
rect 77864 16581 77892 16680
rect 77849 16575 77907 16581
rect 77849 16541 77861 16575
rect 77895 16541 77907 16575
rect 77849 16535 77907 16541
rect 27341 16507 27399 16513
rect 27341 16473 27353 16507
rect 27387 16473 27399 16507
rect 27341 16467 27399 16473
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 26234 16396 26240 16448
rect 26292 16436 26298 16448
rect 26697 16439 26755 16445
rect 26697 16436 26709 16439
rect 26292 16408 26709 16436
rect 26292 16396 26298 16408
rect 26697 16405 26709 16408
rect 26743 16436 26755 16439
rect 27356 16436 27384 16467
rect 78030 16436 78036 16448
rect 26743 16408 27384 16436
rect 77991 16408 78036 16436
rect 26743 16405 26755 16408
rect 26697 16399 26755 16405
rect 78030 16396 78036 16408
rect 78088 16396 78094 16448
rect 1104 16346 78844 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 78844 16346
rect 1104 16272 78844 16294
rect 12710 16232 12716 16244
rect 12671 16204 12716 16232
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 25869 16235 25927 16241
rect 25869 16201 25881 16235
rect 25915 16232 25927 16235
rect 26234 16232 26240 16244
rect 25915 16204 26240 16232
rect 25915 16201 25927 16204
rect 25869 16195 25927 16201
rect 26234 16192 26240 16204
rect 26292 16232 26298 16244
rect 27433 16235 27491 16241
rect 26292 16204 27016 16232
rect 26292 16192 26298 16204
rect 26988 16173 27016 16204
rect 27433 16201 27445 16235
rect 27479 16232 27491 16235
rect 27522 16232 27528 16244
rect 27479 16204 27528 16232
rect 27479 16201 27491 16204
rect 27433 16195 27491 16201
rect 27522 16192 27528 16204
rect 27580 16192 27586 16244
rect 26973 16167 27031 16173
rect 26973 16133 26985 16167
rect 27019 16133 27031 16167
rect 27614 16164 27620 16176
rect 26973 16127 27031 16133
rect 27264 16136 27620 16164
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 12897 16099 12955 16105
rect 1719 16068 6914 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 6886 15960 6914 16068
rect 12897 16065 12909 16099
rect 12943 16065 12955 16099
rect 12897 16059 12955 16065
rect 13633 16099 13691 16105
rect 13633 16065 13645 16099
rect 13679 16096 13691 16099
rect 14090 16096 14096 16108
rect 13679 16068 14096 16096
rect 13679 16065 13691 16068
rect 13633 16059 13691 16065
rect 12912 16028 12940 16059
rect 14090 16056 14096 16068
rect 14148 16056 14154 16108
rect 27264 16105 27292 16136
rect 27614 16124 27620 16136
rect 27672 16164 27678 16176
rect 28166 16164 28172 16176
rect 27672 16136 28172 16164
rect 27672 16124 27678 16136
rect 28166 16124 28172 16136
rect 28224 16124 28230 16176
rect 27249 16099 27307 16105
rect 27249 16065 27261 16099
rect 27295 16065 27307 16099
rect 27249 16059 27307 16065
rect 27985 16099 28043 16105
rect 27985 16065 27997 16099
rect 28031 16065 28043 16099
rect 77665 16099 77723 16105
rect 77665 16096 77677 16099
rect 27985 16059 28043 16065
rect 77128 16068 77677 16096
rect 13814 16028 13820 16040
rect 12912 16000 13820 16028
rect 13814 15988 13820 16000
rect 13872 15988 13878 16040
rect 26418 15988 26424 16040
rect 26476 16028 26482 16040
rect 27065 16031 27123 16037
rect 27065 16028 27077 16031
rect 26476 16000 27077 16028
rect 26476 15988 26482 16000
rect 27065 15997 27077 16000
rect 27111 15997 27123 16031
rect 27065 15991 27123 15997
rect 13449 15963 13507 15969
rect 13449 15960 13461 15963
rect 6886 15932 13461 15960
rect 13449 15929 13461 15932
rect 13495 15929 13507 15963
rect 13449 15923 13507 15929
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 14090 15892 14096 15904
rect 14051 15864 14096 15892
rect 14090 15852 14096 15864
rect 14148 15852 14154 15904
rect 26421 15895 26479 15901
rect 26421 15861 26433 15895
rect 26467 15892 26479 15895
rect 27249 15895 27307 15901
rect 27249 15892 27261 15895
rect 26467 15864 27261 15892
rect 26467 15861 26479 15864
rect 26421 15855 26479 15861
rect 27249 15861 27261 15864
rect 27295 15892 27307 15895
rect 27706 15892 27712 15904
rect 27295 15864 27712 15892
rect 27295 15861 27307 15864
rect 27249 15855 27307 15861
rect 27706 15852 27712 15864
rect 27764 15892 27770 15904
rect 28000 15892 28028 16059
rect 77128 15901 77156 16068
rect 77665 16065 77677 16068
rect 77711 16065 77723 16099
rect 77665 16059 77723 16065
rect 27764 15864 28028 15892
rect 28077 15895 28135 15901
rect 27764 15852 27770 15864
rect 28077 15861 28089 15895
rect 28123 15892 28135 15895
rect 77113 15895 77171 15901
rect 77113 15892 77125 15895
rect 28123 15864 77125 15892
rect 28123 15861 28135 15864
rect 28077 15855 28135 15861
rect 77113 15861 77125 15864
rect 77159 15861 77171 15895
rect 77846 15892 77852 15904
rect 77807 15864 77852 15892
rect 77113 15855 77171 15861
rect 77846 15852 77852 15864
rect 77904 15852 77910 15904
rect 1104 15802 78844 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 78844 15802
rect 1104 15728 78844 15750
rect 14090 15648 14096 15700
rect 14148 15688 14154 15700
rect 27706 15688 27712 15700
rect 14148 15660 27712 15688
rect 14148 15648 14154 15660
rect 27706 15648 27712 15660
rect 27764 15648 27770 15700
rect 26697 15623 26755 15629
rect 26697 15589 26709 15623
rect 26743 15620 26755 15623
rect 27614 15620 27620 15632
rect 26743 15592 27620 15620
rect 26743 15589 26755 15592
rect 26697 15583 26755 15589
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15484 1731 15487
rect 11514 15484 11520 15496
rect 1719 15456 11520 15484
rect 1719 15453 1731 15456
rect 1673 15447 1731 15453
rect 11514 15444 11520 15456
rect 11572 15444 11578 15496
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 13081 15351 13139 15357
rect 13081 15317 13093 15351
rect 13127 15348 13139 15351
rect 13814 15348 13820 15360
rect 13127 15320 13820 15348
rect 13127 15317 13139 15320
rect 13081 15311 13139 15317
rect 13814 15308 13820 15320
rect 13872 15348 13878 15360
rect 14458 15348 14464 15360
rect 13872 15320 14464 15348
rect 13872 15308 13878 15320
rect 14458 15308 14464 15320
rect 14516 15348 14522 15360
rect 26712 15348 26740 15583
rect 27614 15580 27620 15592
rect 27672 15580 27678 15632
rect 77849 15487 77907 15493
rect 77849 15484 77861 15487
rect 77312 15456 77861 15484
rect 27798 15376 27804 15428
rect 27856 15416 27862 15428
rect 77312 15425 77340 15456
rect 77849 15453 77861 15456
rect 77895 15453 77907 15487
rect 77849 15447 77907 15453
rect 77297 15419 77355 15425
rect 77297 15416 77309 15419
rect 27856 15388 77309 15416
rect 27856 15376 27862 15388
rect 77297 15385 77309 15388
rect 77343 15385 77355 15419
rect 77297 15379 77355 15385
rect 78030 15348 78036 15360
rect 14516 15320 26740 15348
rect 77991 15320 78036 15348
rect 14516 15308 14522 15320
rect 78030 15308 78036 15320
rect 78088 15308 78094 15360
rect 1104 15258 78844 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 78844 15258
rect 1104 15184 78844 15206
rect 11514 15144 11520 15156
rect 11475 15116 11520 15144
rect 11514 15104 11520 15116
rect 11572 15104 11578 15156
rect 27709 15079 27767 15085
rect 27709 15045 27721 15079
rect 27755 15076 27767 15079
rect 27798 15076 27804 15088
rect 27755 15048 27804 15076
rect 27755 15045 27767 15048
rect 27709 15039 27767 15045
rect 27798 15036 27804 15048
rect 27856 15036 27862 15088
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 11514 15008 11520 15020
rect 1719 14980 11520 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 26421 15011 26479 15017
rect 11747 14980 12296 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 12268 14813 12296 14980
rect 26421 14977 26433 15011
rect 26467 15008 26479 15011
rect 27062 15008 27068 15020
rect 26467 14980 27068 15008
rect 26467 14977 26479 14980
rect 26421 14971 26479 14977
rect 27062 14968 27068 14980
rect 27120 15008 27126 15020
rect 27525 15011 27583 15017
rect 27525 15008 27537 15011
rect 27120 14980 27537 15008
rect 27120 14968 27126 14980
rect 27525 14977 27537 14980
rect 27571 14977 27583 15011
rect 77665 15011 77723 15017
rect 77665 15008 77677 15011
rect 27525 14971 27583 14977
rect 77128 14980 77677 15008
rect 12253 14807 12311 14813
rect 12253 14773 12265 14807
rect 12299 14804 12311 14807
rect 13354 14804 13360 14816
rect 12299 14776 13360 14804
rect 12299 14773 12311 14776
rect 12253 14767 12311 14773
rect 13354 14764 13360 14776
rect 13412 14764 13418 14816
rect 68002 14764 68008 14816
rect 68060 14804 68066 14816
rect 77128 14813 77156 14980
rect 77665 14977 77677 14980
rect 77711 14977 77723 15011
rect 77665 14971 77723 14977
rect 77113 14807 77171 14813
rect 77113 14804 77125 14807
rect 68060 14776 77125 14804
rect 68060 14764 68066 14776
rect 77113 14773 77125 14776
rect 77159 14773 77171 14807
rect 77846 14804 77852 14816
rect 77807 14776 77852 14804
rect 77113 14767 77171 14773
rect 77846 14764 77852 14776
rect 77904 14764 77910 14816
rect 1104 14714 78844 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 78844 14714
rect 1104 14640 78844 14662
rect 11514 14600 11520 14612
rect 11475 14572 11520 14600
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 11701 14399 11759 14405
rect 11701 14365 11713 14399
rect 11747 14396 11759 14399
rect 11747 14368 12296 14396
rect 11747 14365 11759 14368
rect 11701 14359 11759 14365
rect 12268 14269 12296 14368
rect 26789 14331 26847 14337
rect 26789 14297 26801 14331
rect 26835 14328 26847 14331
rect 26970 14328 26976 14340
rect 26835 14300 26976 14328
rect 26835 14297 26847 14300
rect 26789 14291 26847 14297
rect 26970 14288 26976 14300
rect 27028 14328 27034 14340
rect 27341 14331 27399 14337
rect 27341 14328 27353 14331
rect 27028 14300 27353 14328
rect 27028 14288 27034 14300
rect 27341 14297 27353 14300
rect 27387 14297 27399 14331
rect 27341 14291 27399 14297
rect 12253 14263 12311 14269
rect 12253 14229 12265 14263
rect 12299 14260 12311 14263
rect 12618 14260 12624 14272
rect 12299 14232 12624 14260
rect 12299 14229 12311 14232
rect 12253 14223 12311 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 27433 14263 27491 14269
rect 27433 14229 27445 14263
rect 27479 14260 27491 14263
rect 68002 14260 68008 14272
rect 27479 14232 68008 14260
rect 27479 14229 27491 14232
rect 27433 14223 27491 14229
rect 68002 14220 68008 14232
rect 68060 14220 68066 14272
rect 1104 14170 78844 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 78844 14170
rect 1104 14096 78844 14118
rect 10413 14059 10471 14065
rect 10413 14056 10425 14059
rect 6886 14028 10425 14056
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 6886 13920 6914 14028
rect 10413 14025 10425 14028
rect 10459 14025 10471 14059
rect 10413 14019 10471 14025
rect 12618 14016 12624 14068
rect 12676 14056 12682 14068
rect 26970 14056 26976 14068
rect 12676 14028 26976 14056
rect 12676 14016 12682 14028
rect 26970 14016 26976 14028
rect 27028 14016 27034 14068
rect 27338 14056 27344 14068
rect 27299 14028 27344 14056
rect 27338 14016 27344 14028
rect 27396 14016 27402 14068
rect 77846 14056 77852 14068
rect 77807 14028 77852 14056
rect 77846 14016 77852 14028
rect 77904 14016 77910 14068
rect 26206 13960 27108 13988
rect 1719 13892 6914 13920
rect 10597 13923 10655 13929
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 10643 13892 11652 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 11624 13861 11652 13892
rect 13354 13880 13360 13932
rect 13412 13920 13418 13932
rect 25777 13923 25835 13929
rect 25777 13920 25789 13923
rect 13412 13892 25789 13920
rect 13412 13880 13418 13892
rect 25777 13889 25789 13892
rect 25823 13920 25835 13923
rect 26206 13920 26234 13960
rect 27080 13932 27108 13960
rect 25823 13892 26234 13920
rect 26973 13923 27031 13929
rect 25823 13889 25835 13892
rect 25777 13883 25835 13889
rect 26973 13889 26985 13923
rect 27019 13889 27031 13923
rect 26973 13883 27031 13889
rect 11609 13855 11667 13861
rect 11609 13821 11621 13855
rect 11655 13852 11667 13855
rect 11882 13852 11888 13864
rect 11655 13824 11888 13852
rect 11655 13821 11667 13824
rect 11609 13815 11667 13821
rect 11882 13812 11888 13824
rect 11940 13852 11946 13864
rect 26421 13855 26479 13861
rect 26421 13852 26433 13855
rect 11940 13824 26433 13852
rect 11940 13812 11946 13824
rect 26421 13821 26433 13824
rect 26467 13852 26479 13855
rect 26988 13852 27016 13883
rect 27062 13880 27068 13932
rect 27120 13920 27126 13932
rect 27890 13920 27896 13932
rect 27120 13892 27165 13920
rect 27851 13892 27896 13920
rect 27120 13880 27126 13892
rect 27890 13880 27896 13892
rect 27948 13880 27954 13932
rect 77665 13923 77723 13929
rect 77665 13920 77677 13923
rect 77128 13892 77677 13920
rect 27908 13852 27936 13880
rect 77128 13861 77156 13892
rect 77665 13889 77677 13892
rect 77711 13889 77723 13923
rect 77665 13883 77723 13889
rect 26467 13824 27936 13852
rect 28077 13855 28135 13861
rect 26467 13821 26479 13824
rect 26421 13815 26479 13821
rect 28077 13821 28089 13855
rect 28123 13852 28135 13855
rect 77113 13855 77171 13861
rect 77113 13852 77125 13855
rect 28123 13824 77125 13852
rect 28123 13821 28135 13824
rect 28077 13815 28135 13821
rect 77113 13821 77125 13824
rect 77159 13821 77171 13855
rect 77113 13815 77171 13821
rect 1486 13784 1492 13796
rect 1447 13756 1492 13784
rect 1486 13744 1492 13756
rect 1544 13744 1550 13796
rect 26970 13716 26976 13728
rect 26931 13688 26976 13716
rect 26970 13676 26976 13688
rect 27028 13676 27034 13728
rect 1104 13626 78844 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 78844 13626
rect 1104 13552 78844 13574
rect 26697 13515 26755 13521
rect 26697 13481 26709 13515
rect 26743 13512 26755 13515
rect 26970 13512 26976 13524
rect 26743 13484 26976 13512
rect 26743 13481 26755 13484
rect 26697 13475 26755 13481
rect 26970 13472 26976 13484
rect 27028 13472 27034 13524
rect 27709 13515 27767 13521
rect 27709 13481 27721 13515
rect 27755 13512 27767 13515
rect 27890 13512 27896 13524
rect 27755 13484 27896 13512
rect 27755 13481 27767 13484
rect 27709 13475 27767 13481
rect 27890 13472 27896 13484
rect 27948 13472 27954 13524
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 9585 13311 9643 13317
rect 1719 13280 6914 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 6886 13172 6914 13280
rect 9585 13277 9597 13311
rect 9631 13277 9643 13311
rect 77849 13311 77907 13317
rect 77849 13308 77861 13311
rect 9585 13271 9643 13277
rect 77312 13280 77861 13308
rect 9600 13240 9628 13271
rect 10137 13243 10195 13249
rect 10137 13240 10149 13243
rect 9600 13212 10149 13240
rect 10137 13209 10149 13212
rect 10183 13240 10195 13243
rect 10778 13240 10784 13252
rect 10183 13212 10784 13240
rect 10183 13209 10195 13212
rect 10137 13203 10195 13209
rect 10778 13200 10784 13212
rect 10836 13240 10842 13252
rect 42153 13243 42211 13249
rect 10836 13212 35894 13240
rect 10836 13200 10842 13212
rect 9401 13175 9459 13181
rect 9401 13172 9413 13175
rect 6886 13144 9413 13172
rect 9401 13141 9413 13144
rect 9447 13141 9459 13175
rect 35866 13172 35894 13212
rect 42153 13209 42165 13243
rect 42199 13209 42211 13243
rect 42153 13203 42211 13209
rect 41506 13172 41512 13184
rect 35866 13144 41512 13172
rect 9401 13135 9459 13141
rect 41506 13132 41512 13144
rect 41564 13172 41570 13184
rect 42168 13172 42196 13203
rect 77312 13181 77340 13280
rect 77849 13277 77861 13280
rect 77895 13277 77907 13311
rect 77849 13271 77907 13277
rect 41564 13144 42196 13172
rect 42245 13175 42303 13181
rect 41564 13132 41570 13144
rect 42245 13141 42257 13175
rect 42291 13172 42303 13175
rect 77297 13175 77355 13181
rect 77297 13172 77309 13175
rect 42291 13144 77309 13172
rect 42291 13141 42303 13144
rect 42245 13135 42303 13141
rect 77297 13141 77309 13144
rect 77343 13141 77355 13175
rect 78030 13172 78036 13184
rect 77991 13144 78036 13172
rect 77297 13135 77355 13141
rect 78030 13132 78036 13144
rect 78088 13132 78094 13184
rect 1104 13082 78844 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 78844 13082
rect 1104 13008 78844 13030
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 9674 12832 9680 12844
rect 1719 12804 9680 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 77110 12792 77116 12844
rect 77168 12832 77174 12844
rect 77665 12835 77723 12841
rect 77665 12832 77677 12835
rect 77168 12804 77677 12832
rect 77168 12792 77174 12804
rect 77665 12801 77677 12804
rect 77711 12801 77723 12835
rect 77665 12795 77723 12801
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 77110 12628 77116 12640
rect 77071 12600 77116 12628
rect 77110 12588 77116 12600
rect 77168 12588 77174 12640
rect 77846 12628 77852 12640
rect 77807 12600 77852 12628
rect 77846 12588 77852 12600
rect 77904 12588 77910 12640
rect 1104 12538 78844 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 78844 12538
rect 1104 12464 78844 12486
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 9030 12220 9036 12232
rect 1719 12192 9036 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 9030 12180 9036 12192
rect 9088 12180 9094 12232
rect 9861 12223 9919 12229
rect 9861 12189 9873 12223
rect 9907 12220 9919 12223
rect 10042 12220 10048 12232
rect 9907 12192 10048 12220
rect 9907 12189 9919 12192
rect 9861 12183 9919 12189
rect 10042 12180 10048 12192
rect 10100 12220 10106 12232
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 10100 12192 12633 12220
rect 10100 12180 10106 12192
rect 12621 12189 12633 12192
rect 12667 12189 12679 12223
rect 77849 12223 77907 12229
rect 77849 12220 77861 12223
rect 12621 12183 12679 12189
rect 77312 12192 77861 12220
rect 77312 12096 77340 12192
rect 77849 12189 77861 12192
rect 77895 12189 77907 12223
rect 77849 12183 77907 12189
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12084 12863 12087
rect 77110 12084 77116 12096
rect 12851 12056 77116 12084
rect 12851 12053 12863 12056
rect 12805 12047 12863 12053
rect 77110 12044 77116 12056
rect 77168 12044 77174 12096
rect 77294 12084 77300 12096
rect 77255 12056 77300 12084
rect 77294 12044 77300 12056
rect 77352 12044 77358 12096
rect 78030 12084 78036 12096
rect 77991 12056 78036 12084
rect 78030 12044 78036 12056
rect 78088 12044 78094 12096
rect 1104 11994 78844 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 78844 11994
rect 1104 11920 78844 11942
rect 9030 11880 9036 11892
rect 8991 11852 9036 11880
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9582 11744 9588 11756
rect 9263 11716 9588 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 9582 11704 9588 11716
rect 9640 11744 9646 11756
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 9640 11716 11989 11744
rect 9640 11704 9646 11716
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12161 11543 12219 11549
rect 12161 11509 12173 11543
rect 12207 11540 12219 11543
rect 77294 11540 77300 11552
rect 12207 11512 77300 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 77294 11500 77300 11512
rect 77352 11500 77358 11552
rect 1104 11450 78844 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 78844 11450
rect 1104 11376 78844 11398
rect 1486 11268 1492 11280
rect 1447 11240 1492 11268
rect 1486 11228 1492 11240
rect 1544 11228 1550 11280
rect 78030 11268 78036 11280
rect 77991 11240 78036 11268
rect 78030 11228 78036 11240
rect 78088 11228 78094 11280
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 8294 11132 8300 11144
rect 1719 11104 8300 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 77849 11135 77907 11141
rect 77849 11132 77861 11135
rect 77312 11104 77861 11132
rect 11698 11024 11704 11076
rect 11756 11064 11762 11076
rect 77312 11073 77340 11104
rect 77849 11101 77861 11104
rect 77895 11101 77907 11135
rect 77849 11095 77907 11101
rect 77297 11067 77355 11073
rect 77297 11064 77309 11067
rect 11756 11036 77309 11064
rect 11756 11024 11762 11036
rect 77297 11033 77309 11036
rect 77343 11033 77355 11067
rect 77297 11027 77355 11033
rect 1104 10906 78844 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 78844 10906
rect 1104 10832 78844 10854
rect 8294 10792 8300 10804
rect 8255 10764 8300 10792
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 11698 10792 11704 10804
rect 11659 10764 11704 10792
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 7558 10656 7564 10668
rect 1719 10628 7564 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 7558 10616 7564 10628
rect 7616 10616 7622 10668
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 8938 10656 8944 10668
rect 8527 10628 8944 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 8938 10616 8944 10628
rect 8996 10656 9002 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 8996 10628 11529 10656
rect 8996 10616 9002 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 77665 10659 77723 10665
rect 77665 10656 77677 10659
rect 11517 10619 11575 10625
rect 77128 10628 77677 10656
rect 77128 10464 77156 10628
rect 77665 10625 77677 10628
rect 77711 10625 77723 10659
rect 77665 10619 77723 10625
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 77110 10452 77116 10464
rect 77071 10424 77116 10452
rect 77110 10412 77116 10424
rect 77168 10412 77174 10464
rect 77846 10452 77852 10464
rect 77807 10424 77852 10452
rect 77846 10412 77852 10424
rect 77904 10412 77910 10464
rect 1104 10362 78844 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 78844 10362
rect 1104 10288 78844 10310
rect 7558 10248 7564 10260
rect 7519 10220 7564 10248
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 6730 10044 6736 10056
rect 1719 10016 6736 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 8202 10044 8208 10056
rect 7791 10016 8208 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 8202 10004 8208 10016
rect 8260 10044 8266 10056
rect 10689 10047 10747 10053
rect 10689 10044 10701 10047
rect 8260 10016 10701 10044
rect 8260 10004 8266 10016
rect 10689 10013 10701 10016
rect 10735 10013 10747 10047
rect 77849 10047 77907 10053
rect 77849 10044 77861 10047
rect 10689 10007 10747 10013
rect 77312 10016 77861 10044
rect 77110 9976 77116 9988
rect 10888 9948 77116 9976
rect 1486 9908 1492 9920
rect 1447 9880 1492 9908
rect 1486 9868 1492 9880
rect 1544 9868 1550 9920
rect 10888 9917 10916 9948
rect 77110 9936 77116 9948
rect 77168 9936 77174 9988
rect 10873 9911 10931 9917
rect 10873 9877 10885 9911
rect 10919 9877 10931 9911
rect 10873 9871 10931 9877
rect 10962 9868 10968 9920
rect 11020 9908 11026 9920
rect 77312 9917 77340 10016
rect 77849 10013 77861 10016
rect 77895 10013 77907 10047
rect 77849 10007 77907 10013
rect 77297 9911 77355 9917
rect 77297 9908 77309 9911
rect 11020 9880 77309 9908
rect 11020 9868 11026 9880
rect 77297 9877 77309 9880
rect 77343 9877 77355 9911
rect 78030 9908 78036 9920
rect 77991 9880 78036 9908
rect 77297 9871 77355 9877
rect 78030 9868 78036 9880
rect 78088 9868 78094 9920
rect 1104 9818 78844 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 78844 9818
rect 1104 9744 78844 9766
rect 6730 9704 6736 9716
rect 6691 9676 6736 9704
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 10137 9707 10195 9713
rect 10137 9673 10149 9707
rect 10183 9704 10195 9707
rect 10962 9704 10968 9716
rect 10183 9676 10968 9704
rect 10183 9673 10195 9676
rect 10137 9667 10195 9673
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 5994 9568 6000 9580
rect 1719 9540 6000 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 9953 9571 10011 9577
rect 9953 9568 9965 9571
rect 6972 9540 9965 9568
rect 6972 9528 6978 9540
rect 9953 9537 9965 9540
rect 9999 9537 10011 9571
rect 77665 9571 77723 9577
rect 77665 9568 77677 9571
rect 9953 9531 10011 9537
rect 77128 9540 77677 9568
rect 1486 9364 1492 9376
rect 1447 9336 1492 9364
rect 1486 9324 1492 9336
rect 1544 9324 1550 9376
rect 69658 9324 69664 9376
rect 69716 9364 69722 9376
rect 77128 9373 77156 9540
rect 77665 9537 77677 9540
rect 77711 9537 77723 9571
rect 77665 9531 77723 9537
rect 77113 9367 77171 9373
rect 77113 9364 77125 9367
rect 69716 9336 77125 9364
rect 69716 9324 69722 9336
rect 77113 9333 77125 9336
rect 77159 9333 77171 9367
rect 77846 9364 77852 9376
rect 77807 9336 77852 9364
rect 77113 9327 77171 9333
rect 77846 9324 77852 9336
rect 77904 9324 77910 9376
rect 1104 9274 78844 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 78844 9274
rect 1104 9200 78844 9222
rect 5994 9160 6000 9172
rect 5955 9132 6000 9160
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6178 8956 6184 8968
rect 6139 8928 6184 8956
rect 6178 8916 6184 8928
rect 6236 8956 6242 8968
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 6236 8928 9321 8956
rect 6236 8916 6242 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9493 8823 9551 8829
rect 9493 8789 9505 8823
rect 9539 8820 9551 8823
rect 69658 8820 69664 8832
rect 9539 8792 69664 8820
rect 9539 8789 9551 8792
rect 9493 8783 9551 8789
rect 69658 8780 69664 8792
rect 69716 8780 69722 8832
rect 1104 8730 78844 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 78844 8730
rect 1104 8656 78844 8678
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 5258 8480 5264 8492
rect 1719 8452 5264 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 77665 8483 77723 8489
rect 77665 8480 77677 8483
rect 77128 8452 77677 8480
rect 77128 8356 77156 8452
rect 77665 8449 77677 8452
rect 77711 8449 77723 8483
rect 77665 8443 77723 8449
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 77110 8344 77116 8356
rect 77071 8316 77116 8344
rect 77110 8304 77116 8316
rect 77168 8304 77174 8356
rect 77846 8344 77852 8356
rect 77807 8316 77852 8344
rect 77846 8304 77852 8316
rect 77904 8304 77910 8356
rect 1104 8186 78844 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 78844 8186
rect 1104 8112 78844 8134
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 4522 7868 4528 7880
rect 1719 7840 4528 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7868 5503 7871
rect 5626 7868 5632 7880
rect 5491 7840 5632 7868
rect 5491 7837 5503 7840
rect 5445 7831 5503 7837
rect 5626 7828 5632 7840
rect 5684 7868 5690 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 5684 7840 8953 7868
rect 5684 7828 5690 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 77849 7871 77907 7877
rect 77849 7868 77861 7871
rect 8941 7831 8999 7837
rect 77312 7840 77861 7868
rect 77018 7760 77024 7812
rect 77076 7800 77082 7812
rect 77312 7809 77340 7840
rect 77849 7837 77861 7840
rect 77895 7837 77907 7871
rect 77849 7831 77907 7837
rect 77297 7803 77355 7809
rect 77297 7800 77309 7803
rect 77076 7772 77309 7800
rect 77076 7760 77082 7772
rect 77297 7769 77309 7772
rect 77343 7769 77355 7803
rect 77297 7763 77355 7769
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 9125 7735 9183 7741
rect 9125 7701 9137 7735
rect 9171 7732 9183 7735
rect 77110 7732 77116 7744
rect 9171 7704 77116 7732
rect 9171 7701 9183 7704
rect 9125 7695 9183 7701
rect 77110 7692 77116 7704
rect 77168 7692 77174 7744
rect 78030 7732 78036 7744
rect 77991 7704 78036 7732
rect 78030 7692 78036 7704
rect 78088 7692 78094 7744
rect 1104 7642 78844 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 78844 7642
rect 1104 7568 78844 7590
rect 4522 7528 4528 7540
rect 4483 7500 4528 7528
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 3878 7392 3884 7404
rect 1719 7364 3884 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 4706 7392 4712 7404
rect 4619 7364 4712 7392
rect 4706 7352 4712 7364
rect 4764 7392 4770 7404
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 4764 7364 8033 7392
rect 4764 7352 4770 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 77665 7395 77723 7401
rect 77665 7392 77677 7395
rect 8021 7355 8079 7361
rect 77128 7364 77677 7392
rect 8205 7259 8263 7265
rect 8205 7225 8217 7259
rect 8251 7256 8263 7259
rect 77018 7256 77024 7268
rect 8251 7228 77024 7256
rect 8251 7225 8263 7228
rect 8205 7219 8263 7225
rect 77018 7216 77024 7228
rect 77076 7216 77082 7268
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 76006 7148 76012 7200
rect 76064 7188 76070 7200
rect 77128 7197 77156 7364
rect 77665 7361 77677 7364
rect 77711 7361 77723 7395
rect 77665 7355 77723 7361
rect 77113 7191 77171 7197
rect 77113 7188 77125 7191
rect 76064 7160 77125 7188
rect 76064 7148 76070 7160
rect 77113 7157 77125 7160
rect 77159 7157 77171 7191
rect 77846 7188 77852 7200
rect 77807 7160 77852 7188
rect 77113 7151 77171 7157
rect 77846 7148 77852 7160
rect 77904 7148 77910 7200
rect 1104 7098 78844 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 78844 7098
rect 1104 7024 78844 7046
rect 3878 6984 3884 6996
rect 3839 6956 3884 6984
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 3234 6780 3240 6792
rect 1719 6752 3240 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6780 4123 6783
rect 4614 6780 4620 6792
rect 4111 6752 4620 6780
rect 4111 6749 4123 6752
rect 4065 6743 4123 6749
rect 4614 6740 4620 6752
rect 4672 6780 4678 6792
rect 7469 6783 7527 6789
rect 7469 6780 7481 6783
rect 4672 6752 7481 6780
rect 4672 6740 4678 6752
rect 7469 6749 7481 6752
rect 7515 6749 7527 6783
rect 77849 6783 77907 6789
rect 77849 6780 77861 6783
rect 7469 6743 7527 6749
rect 77312 6752 77861 6780
rect 77312 6656 77340 6752
rect 77849 6749 77861 6752
rect 77895 6749 77907 6783
rect 77849 6743 77907 6749
rect 1486 6644 1492 6656
rect 1447 6616 1492 6644
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6644 7711 6647
rect 76006 6644 76012 6656
rect 7699 6616 76012 6644
rect 7699 6613 7711 6616
rect 7653 6607 7711 6613
rect 76006 6604 76012 6616
rect 76064 6604 76070 6656
rect 77294 6644 77300 6656
rect 77255 6616 77300 6644
rect 77294 6604 77300 6616
rect 77352 6604 77358 6656
rect 78030 6644 78036 6656
rect 77991 6616 78036 6644
rect 78030 6604 78036 6616
rect 78088 6604 78094 6656
rect 1104 6554 78844 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 78844 6554
rect 1104 6480 78844 6502
rect 3234 6440 3240 6452
rect 3195 6412 3240 6440
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3786 6304 3792 6316
rect 3467 6276 3792 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3786 6264 3792 6276
rect 3844 6304 3850 6316
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 3844 6276 6929 6304
rect 3844 6264 3850 6276
rect 6917 6273 6929 6276
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 7101 6103 7159 6109
rect 7101 6069 7113 6103
rect 7147 6100 7159 6103
rect 77294 6100 77300 6112
rect 7147 6072 77300 6100
rect 7147 6069 7159 6072
rect 7101 6063 7159 6069
rect 77294 6060 77300 6072
rect 77352 6060 77358 6112
rect 1104 6010 78844 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 78844 6010
rect 1104 5936 78844 5958
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 77297 5695 77355 5701
rect 77297 5692 77309 5695
rect 6696 5664 77309 5692
rect 6696 5652 6702 5664
rect 77297 5661 77309 5664
rect 77343 5692 77355 5695
rect 77849 5695 77907 5701
rect 77849 5692 77861 5695
rect 77343 5664 77861 5692
rect 77343 5661 77355 5664
rect 77297 5655 77355 5661
rect 77849 5661 77861 5664
rect 77895 5661 77907 5695
rect 77849 5655 77907 5661
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 78030 5556 78036 5568
rect 77991 5528 78036 5556
rect 78030 5516 78036 5528
rect 78088 5516 78094 5568
rect 1104 5466 78844 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 78844 5466
rect 1104 5392 78844 5414
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 1728 5324 2605 5352
rect 1728 5312 1734 5324
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 6638 5352 6644 5364
rect 6599 5324 6644 5352
rect 2593 5315 2651 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 2038 5216 2044 5228
rect 1719 5188 2044 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 3050 5216 3056 5228
rect 2823 5188 3056 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 3050 5176 3056 5188
rect 3108 5216 3114 5228
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 3108 5188 6469 5216
rect 3108 5176 3114 5188
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 77665 5219 77723 5225
rect 77665 5216 77677 5219
rect 6457 5179 6515 5185
rect 77128 5188 77677 5216
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 69658 4972 69664 5024
rect 69716 5012 69722 5024
rect 77128 5021 77156 5188
rect 77665 5185 77677 5188
rect 77711 5185 77723 5219
rect 77665 5179 77723 5185
rect 77113 5015 77171 5021
rect 77113 5012 77125 5015
rect 69716 4984 77125 5012
rect 69716 4972 69722 4984
rect 77113 4981 77125 4984
rect 77159 4981 77171 5015
rect 77846 5012 77852 5024
rect 77807 4984 77852 5012
rect 77113 4975 77171 4981
rect 77846 4972 77852 4984
rect 77904 4972 77910 5024
rect 1104 4922 78844 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 78844 4922
rect 1104 4848 78844 4870
rect 2038 4808 2044 4820
rect 1999 4780 2044 4808
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4604 2283 4607
rect 2314 4604 2320 4616
rect 2271 4576 2320 4604
rect 2271 4573 2283 4576
rect 2225 4567 2283 4573
rect 2314 4564 2320 4576
rect 2372 4604 2378 4616
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 2372 4576 6009 4604
rect 2372 4564 2378 4576
rect 5997 4573 6009 4576
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 6181 4471 6239 4477
rect 6181 4437 6193 4471
rect 6227 4468 6239 4471
rect 69658 4468 69664 4480
rect 6227 4440 69664 4468
rect 6227 4437 6239 4440
rect 6181 4431 6239 4437
rect 69658 4428 69664 4440
rect 69716 4428 69722 4480
rect 1104 4378 78844 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 78844 4378
rect 1104 4304 78844 4326
rect 1104 3834 78844 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 78844 3834
rect 1104 3760 78844 3782
rect 53834 3720 53840 3732
rect 53795 3692 53840 3720
rect 53834 3680 53840 3692
rect 53892 3680 53898 3732
rect 64322 3720 64328 3732
rect 64283 3692 64328 3720
rect 64322 3680 64328 3692
rect 64380 3680 64386 3732
rect 27433 3587 27491 3593
rect 27433 3553 27445 3587
rect 27479 3584 27491 3587
rect 27522 3584 27528 3596
rect 27479 3556 27528 3584
rect 27479 3553 27491 3556
rect 27433 3547 27491 3553
rect 27522 3544 27528 3556
rect 27580 3544 27586 3596
rect 63862 3544 63868 3596
rect 63920 3584 63926 3596
rect 69477 3587 69535 3593
rect 69477 3584 69489 3587
rect 63920 3556 69489 3584
rect 63920 3544 63926 3556
rect 69477 3553 69489 3556
rect 69523 3584 69535 3587
rect 69658 3584 69664 3596
rect 69523 3556 69664 3584
rect 69523 3553 69535 3556
rect 69477 3547 69535 3553
rect 69658 3544 69664 3556
rect 69716 3544 69722 3596
rect 26697 3519 26755 3525
rect 26697 3485 26709 3519
rect 26743 3516 26755 3519
rect 27062 3516 27068 3528
rect 26743 3488 27068 3516
rect 26743 3485 26755 3488
rect 26697 3479 26755 3485
rect 27062 3476 27068 3488
rect 27120 3516 27126 3528
rect 27157 3519 27215 3525
rect 27157 3516 27169 3519
rect 27120 3488 27169 3516
rect 27120 3476 27126 3488
rect 27157 3485 27169 3488
rect 27203 3485 27215 3519
rect 27157 3479 27215 3485
rect 29270 3408 29276 3460
rect 29328 3448 29334 3460
rect 30469 3451 30527 3457
rect 30469 3448 30481 3451
rect 29328 3420 30481 3448
rect 29328 3408 29334 3420
rect 30469 3417 30481 3420
rect 30515 3417 30527 3451
rect 30469 3411 30527 3417
rect 66162 3408 66168 3460
rect 66220 3448 66226 3460
rect 70578 3448 70584 3460
rect 66220 3420 70584 3448
rect 66220 3408 66226 3420
rect 70578 3408 70584 3420
rect 70636 3408 70642 3460
rect 28442 3380 28448 3392
rect 28403 3352 28448 3380
rect 28442 3340 28448 3352
rect 28500 3340 28506 3392
rect 30006 3380 30012 3392
rect 29967 3352 30012 3380
rect 30006 3340 30012 3352
rect 30064 3340 30070 3392
rect 32214 3380 32220 3392
rect 32175 3352 32220 3380
rect 32214 3340 32220 3352
rect 32272 3340 32278 3392
rect 32950 3380 32956 3392
rect 32911 3352 32956 3380
rect 32950 3340 32956 3352
rect 33008 3340 33014 3392
rect 33686 3380 33692 3392
rect 33647 3352 33692 3380
rect 33686 3340 33692 3352
rect 33744 3340 33750 3392
rect 43714 3380 43720 3392
rect 43675 3352 43720 3380
rect 43714 3340 43720 3352
rect 43772 3340 43778 3392
rect 74718 3380 74724 3392
rect 74679 3352 74724 3380
rect 74718 3340 74724 3352
rect 74776 3340 74782 3392
rect 77846 3340 77852 3392
rect 77904 3380 77910 3392
rect 78033 3383 78091 3389
rect 78033 3380 78045 3383
rect 77904 3352 78045 3380
rect 77904 3340 77910 3352
rect 78033 3349 78045 3352
rect 78079 3349 78091 3383
rect 78033 3343 78091 3349
rect 1104 3290 78844 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 78844 3290
rect 1104 3216 78844 3238
rect 3786 3176 3792 3188
rect 3747 3148 3792 3176
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 8938 3176 8944 3188
rect 8899 3148 8944 3176
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 14090 3176 14096 3188
rect 14051 3148 14096 3176
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 24394 3176 24400 3188
rect 24355 3148 24400 3176
rect 24394 3136 24400 3148
rect 24452 3136 24458 3188
rect 32490 3176 32496 3188
rect 32451 3148 32496 3176
rect 32490 3136 32496 3148
rect 32548 3136 32554 3188
rect 33226 3176 33232 3188
rect 33187 3148 33232 3176
rect 33226 3136 33232 3148
rect 33284 3136 33290 3188
rect 34698 3176 34704 3188
rect 34659 3148 34704 3176
rect 34698 3136 34704 3148
rect 34756 3136 34762 3188
rect 39850 3176 39856 3188
rect 39811 3148 39856 3176
rect 39850 3136 39856 3148
rect 39908 3136 39914 3188
rect 44266 3176 44272 3188
rect 44227 3148 44272 3176
rect 44266 3136 44272 3148
rect 44324 3136 44330 3188
rect 49970 3176 49976 3188
rect 49931 3148 49976 3176
rect 49970 3136 49976 3148
rect 50028 3136 50034 3188
rect 50614 3176 50620 3188
rect 50575 3148 50620 3176
rect 50614 3136 50620 3148
rect 50672 3136 50678 3188
rect 51258 3176 51264 3188
rect 51219 3148 51264 3176
rect 51258 3136 51264 3148
rect 51316 3136 51322 3188
rect 51810 3176 51816 3188
rect 51771 3148 51816 3176
rect 51810 3136 51816 3148
rect 51868 3136 51874 3188
rect 52362 3136 52368 3188
rect 52420 3176 52426 3188
rect 52733 3179 52791 3185
rect 52733 3176 52745 3179
rect 52420 3148 52745 3176
rect 52420 3136 52426 3148
rect 52733 3145 52745 3148
rect 52779 3145 52791 3179
rect 53282 3176 53288 3188
rect 53243 3148 53288 3176
rect 52733 3139 52791 3145
rect 53282 3136 53288 3148
rect 53340 3136 53346 3188
rect 55217 3179 55275 3185
rect 55217 3145 55229 3179
rect 55263 3176 55275 3179
rect 55398 3176 55404 3188
rect 55263 3148 55404 3176
rect 55263 3145 55275 3148
rect 55217 3139 55275 3145
rect 55398 3136 55404 3148
rect 55456 3136 55462 3188
rect 56505 3179 56563 3185
rect 56505 3145 56517 3179
rect 56551 3176 56563 3179
rect 56594 3176 56600 3188
rect 56551 3148 56600 3176
rect 56551 3145 56563 3148
rect 56505 3139 56563 3145
rect 56594 3136 56600 3148
rect 56652 3136 56658 3188
rect 57146 3176 57152 3188
rect 57107 3148 57152 3176
rect 57146 3136 57152 3148
rect 57204 3136 57210 3188
rect 58434 3176 58440 3188
rect 58395 3148 58440 3176
rect 58434 3136 58440 3148
rect 58492 3136 58498 3188
rect 58986 3176 58992 3188
rect 58947 3148 58992 3176
rect 58986 3136 58992 3148
rect 59044 3136 59050 3188
rect 60274 3176 60280 3188
rect 60235 3148 60280 3176
rect 60274 3136 60280 3148
rect 60332 3136 60338 3188
rect 60642 3136 60648 3188
rect 60700 3176 60706 3188
rect 60829 3179 60887 3185
rect 60829 3176 60841 3179
rect 60700 3148 60841 3176
rect 60700 3136 60706 3148
rect 60829 3145 60841 3148
rect 60875 3145 60887 3179
rect 60829 3139 60887 3145
rect 63310 3136 63316 3188
rect 63368 3176 63374 3188
rect 64141 3179 64199 3185
rect 64141 3176 64153 3179
rect 63368 3148 64153 3176
rect 63368 3136 63374 3148
rect 64141 3145 64153 3148
rect 64187 3145 64199 3179
rect 64141 3139 64199 3145
rect 19334 3108 19340 3120
rect 19295 3080 19340 3108
rect 19334 3068 19340 3080
rect 19392 3068 19398 3120
rect 3510 3000 3516 3052
rect 3568 3040 3574 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3568 3012 3617 3040
rect 3568 3000 3574 3012
rect 3605 3009 3617 3012
rect 3651 3040 3663 3043
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 3651 3012 4261 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 8662 3040 8668 3052
rect 8343 3012 8668 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 8662 3000 8668 3012
rect 8720 3040 8726 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 8720 3012 8769 3040
rect 8720 3000 8726 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3040 13507 3043
rect 13814 3040 13820 3052
rect 13495 3012 13820 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 13814 3000 13820 3012
rect 13872 3040 13878 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13872 3012 14013 3040
rect 13872 3000 13878 3012
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 18601 3043 18659 3049
rect 18601 3009 18613 3043
rect 18647 3040 18659 3043
rect 18966 3040 18972 3052
rect 18647 3012 18972 3040
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 18966 3000 18972 3012
rect 19024 3040 19030 3052
rect 19153 3043 19211 3049
rect 19153 3040 19165 3043
rect 19024 3012 19165 3040
rect 19024 3000 19030 3012
rect 19153 3009 19165 3012
rect 19199 3009 19211 3043
rect 19153 3003 19211 3009
rect 23753 3043 23811 3049
rect 23753 3009 23765 3043
rect 23799 3040 23811 3043
rect 24118 3040 24124 3052
rect 23799 3012 24124 3040
rect 23799 3009 23811 3012
rect 23753 3003 23811 3009
rect 24118 3000 24124 3012
rect 24176 3040 24182 3052
rect 24305 3043 24363 3049
rect 24305 3040 24317 3043
rect 24176 3012 24317 3040
rect 24176 3000 24182 3012
rect 24305 3009 24317 3012
rect 24351 3009 24363 3043
rect 24305 3003 24363 3009
rect 26050 3000 26056 3052
rect 26108 3040 26114 3052
rect 26145 3043 26203 3049
rect 26145 3040 26157 3043
rect 26108 3012 26157 3040
rect 26108 3000 26114 3012
rect 26145 3009 26157 3012
rect 26191 3009 26203 3043
rect 26145 3003 26203 3009
rect 27982 3000 27988 3052
rect 28040 3040 28046 3052
rect 28077 3043 28135 3049
rect 28077 3040 28089 3043
rect 28040 3012 28089 3040
rect 28040 3000 28046 3012
rect 28077 3009 28089 3012
rect 28123 3009 28135 3043
rect 29362 3040 29368 3052
rect 29323 3012 29368 3040
rect 28077 3003 28135 3009
rect 29362 3000 29368 3012
rect 29420 3000 29426 3052
rect 30374 3040 30380 3052
rect 30335 3012 30380 3040
rect 30374 3000 30380 3012
rect 30432 3000 30438 3052
rect 32214 3000 32220 3052
rect 32272 3040 32278 3052
rect 32401 3043 32459 3049
rect 32401 3040 32413 3043
rect 32272 3012 32413 3040
rect 32272 3000 32278 3012
rect 32401 3009 32413 3012
rect 32447 3009 32459 3043
rect 32401 3003 32459 3009
rect 32950 3000 32956 3052
rect 33008 3040 33014 3052
rect 33137 3043 33195 3049
rect 33137 3040 33149 3043
rect 33008 3012 33149 3040
rect 33008 3000 33014 3012
rect 33137 3009 33149 3012
rect 33183 3009 33195 3043
rect 33137 3003 33195 3009
rect 34057 3043 34115 3049
rect 34057 3009 34069 3043
rect 34103 3040 34115 3043
rect 34422 3040 34428 3052
rect 34103 3012 34428 3040
rect 34103 3009 34115 3012
rect 34057 3003 34115 3009
rect 34422 3000 34428 3012
rect 34480 3040 34486 3052
rect 34609 3043 34667 3049
rect 34609 3040 34621 3043
rect 34480 3012 34621 3040
rect 34480 3000 34486 3012
rect 34609 3009 34621 3012
rect 34655 3009 34667 3043
rect 34609 3003 34667 3009
rect 39209 3043 39267 3049
rect 39209 3009 39221 3043
rect 39255 3040 39267 3043
rect 39574 3040 39580 3052
rect 39255 3012 39580 3040
rect 39255 3009 39267 3012
rect 39209 3003 39267 3009
rect 39574 3000 39580 3012
rect 39632 3040 39638 3052
rect 39761 3043 39819 3049
rect 39761 3040 39773 3043
rect 39632 3012 39773 3040
rect 39632 3000 39638 3012
rect 39761 3009 39773 3012
rect 39807 3009 39819 3043
rect 39761 3003 39819 3009
rect 43625 3043 43683 3049
rect 43625 3009 43637 3043
rect 43671 3040 43683 3043
rect 43990 3040 43996 3052
rect 43671 3012 43996 3040
rect 43671 3009 43683 3012
rect 43625 3003 43683 3009
rect 43990 3000 43996 3012
rect 44048 3040 44054 3052
rect 44177 3043 44235 3049
rect 44177 3040 44189 3043
rect 44048 3012 44189 3040
rect 44048 3000 44054 3012
rect 44177 3009 44189 3012
rect 44223 3009 44235 3043
rect 44177 3003 44235 3009
rect 49513 3043 49571 3049
rect 49513 3009 49525 3043
rect 49559 3040 49571 3043
rect 49988 3040 50016 3136
rect 52086 3068 52092 3120
rect 52144 3108 52150 3120
rect 53837 3111 53895 3117
rect 53837 3108 53849 3111
rect 52144 3080 53849 3108
rect 52144 3068 52150 3080
rect 53837 3077 53849 3080
rect 53883 3108 53895 3111
rect 53883 3080 54432 3108
rect 53883 3077 53895 3080
rect 53837 3071 53895 3077
rect 54404 3049 54432 3080
rect 57054 3068 57060 3120
rect 57112 3108 57118 3120
rect 57882 3108 57888 3120
rect 57112 3080 57888 3108
rect 57112 3068 57118 3080
rect 57882 3068 57888 3080
rect 57940 3108 57946 3120
rect 57977 3111 58035 3117
rect 57977 3108 57989 3111
rect 57940 3080 57989 3108
rect 57940 3068 57946 3080
rect 57977 3077 57989 3080
rect 58023 3077 58035 3111
rect 57977 3071 58035 3077
rect 49559 3012 50016 3040
rect 54389 3043 54447 3049
rect 49559 3009 49571 3012
rect 49513 3003 49571 3009
rect 54389 3009 54401 3043
rect 54435 3009 54447 3043
rect 54389 3003 54447 3009
rect 59817 3043 59875 3049
rect 59817 3009 59829 3043
rect 59863 3040 59875 3043
rect 60292 3040 60320 3136
rect 60550 3068 60556 3120
rect 60608 3108 60614 3120
rect 61381 3111 61439 3117
rect 61381 3108 61393 3111
rect 60608 3080 61393 3108
rect 60608 3068 60614 3080
rect 61381 3077 61393 3080
rect 61427 3077 61439 3111
rect 61381 3071 61439 3077
rect 62390 3068 62396 3120
rect 62448 3108 62454 3120
rect 63402 3108 63408 3120
rect 62448 3080 63408 3108
rect 62448 3068 62454 3080
rect 63402 3068 63408 3080
rect 63460 3108 63466 3120
rect 63589 3111 63647 3117
rect 63589 3108 63601 3111
rect 63460 3080 63601 3108
rect 63460 3068 63466 3080
rect 63589 3077 63601 3080
rect 63635 3077 63647 3111
rect 63589 3071 63647 3077
rect 59863 3012 60320 3040
rect 64156 3040 64184 3139
rect 65242 3136 65248 3188
rect 65300 3176 65306 3188
rect 66162 3176 66168 3188
rect 65300 3148 66168 3176
rect 65300 3136 65306 3148
rect 66162 3136 66168 3148
rect 66220 3176 66226 3188
rect 66901 3179 66959 3185
rect 66901 3176 66913 3179
rect 66220 3148 66913 3176
rect 66220 3136 66226 3148
rect 66901 3145 66913 3148
rect 66947 3145 66959 3179
rect 69290 3176 69296 3188
rect 69251 3148 69296 3176
rect 66901 3139 66959 3145
rect 69290 3136 69296 3148
rect 69348 3136 69354 3188
rect 70578 3176 70584 3188
rect 70539 3148 70584 3176
rect 70578 3136 70584 3148
rect 70636 3136 70642 3188
rect 72050 3176 72056 3188
rect 72011 3148 72056 3176
rect 72050 3136 72056 3148
rect 72108 3136 72114 3188
rect 75181 3179 75239 3185
rect 75181 3145 75193 3179
rect 75227 3176 75239 3179
rect 75914 3176 75920 3188
rect 75227 3148 75920 3176
rect 75227 3145 75239 3148
rect 75181 3139 75239 3145
rect 75914 3136 75920 3148
rect 75972 3136 75978 3188
rect 77757 3179 77815 3185
rect 77757 3145 77769 3179
rect 77803 3145 77815 3179
rect 77757 3139 77815 3145
rect 65058 3068 65064 3120
rect 65116 3108 65122 3120
rect 68186 3108 68192 3120
rect 65116 3080 68192 3108
rect 65116 3068 65122 3080
rect 68186 3068 68192 3080
rect 68244 3068 68250 3120
rect 64693 3043 64751 3049
rect 64693 3040 64705 3043
rect 64156 3012 64705 3040
rect 59863 3009 59875 3012
rect 59817 3003 59875 3009
rect 64693 3009 64705 3012
rect 64739 3009 64751 3043
rect 64693 3003 64751 3009
rect 65150 3000 65156 3052
rect 65208 3040 65214 3052
rect 68741 3043 68799 3049
rect 68741 3040 68753 3043
rect 65208 3012 68753 3040
rect 65208 3000 65214 3012
rect 68741 3009 68753 3012
rect 68787 3040 68799 3043
rect 68922 3040 68928 3052
rect 68787 3012 68928 3040
rect 68787 3009 68799 3012
rect 68741 3003 68799 3009
rect 68922 3000 68928 3012
rect 68980 3000 68986 3052
rect 69308 3040 69336 3136
rect 77772 3108 77800 3139
rect 69952 3080 77800 3108
rect 69845 3043 69903 3049
rect 69845 3040 69857 3043
rect 69308 3012 69857 3040
rect 69845 3009 69857 3012
rect 69891 3009 69903 3043
rect 69845 3003 69903 3009
rect 25590 2932 25596 2984
rect 25648 2972 25654 2984
rect 26421 2975 26479 2981
rect 26421 2972 26433 2975
rect 25648 2944 26433 2972
rect 25648 2932 25654 2944
rect 26421 2941 26433 2944
rect 26467 2972 26479 2975
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26467 2944 26985 2972
rect 26467 2941 26479 2944
rect 26421 2935 26479 2941
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 27798 2932 27804 2984
rect 27856 2972 27862 2984
rect 28353 2975 28411 2981
rect 28353 2972 28365 2975
rect 27856 2944 28365 2972
rect 27856 2932 27862 2944
rect 28353 2941 28365 2944
rect 28399 2972 28411 2975
rect 28442 2972 28448 2984
rect 28399 2944 28448 2972
rect 28399 2941 28411 2944
rect 28353 2935 28411 2941
rect 28442 2932 28448 2944
rect 28500 2932 28506 2984
rect 29270 2932 29276 2984
rect 29328 2972 29334 2984
rect 29641 2975 29699 2981
rect 29641 2972 29653 2975
rect 29328 2944 29653 2972
rect 29328 2932 29334 2944
rect 29641 2941 29653 2944
rect 29687 2941 29699 2975
rect 29641 2935 29699 2941
rect 30006 2932 30012 2984
rect 30064 2972 30070 2984
rect 30101 2975 30159 2981
rect 30101 2972 30113 2975
rect 30064 2944 30113 2972
rect 30064 2932 30070 2944
rect 30101 2941 30113 2944
rect 30147 2941 30159 2975
rect 30101 2935 30159 2941
rect 59906 2932 59912 2984
rect 59964 2972 59970 2984
rect 61930 2972 61936 2984
rect 59964 2944 61936 2972
rect 59964 2932 59970 2944
rect 61930 2932 61936 2944
rect 61988 2932 61994 2984
rect 62482 2932 62488 2984
rect 62540 2972 62546 2984
rect 65426 2972 65432 2984
rect 62540 2944 65432 2972
rect 62540 2932 62546 2944
rect 65426 2932 65432 2944
rect 65484 2932 65490 2984
rect 65518 2932 65524 2984
rect 65576 2972 65582 2984
rect 69952 2972 69980 3080
rect 74537 3043 74595 3049
rect 74537 3009 74549 3043
rect 74583 3040 74595 3043
rect 74902 3040 74908 3052
rect 74583 3012 74908 3040
rect 74583 3009 74595 3012
rect 74537 3003 74595 3009
rect 74902 3000 74908 3012
rect 74960 3040 74966 3052
rect 74997 3043 75055 3049
rect 74997 3040 75009 3043
rect 74960 3012 75009 3040
rect 74960 3000 74966 3012
rect 74997 3009 75009 3012
rect 75043 3009 75055 3043
rect 74997 3003 75055 3009
rect 77846 3000 77852 3052
rect 77904 3040 77910 3052
rect 77941 3043 77999 3049
rect 77941 3040 77953 3043
rect 77904 3012 77953 3040
rect 77904 3000 77910 3012
rect 77941 3009 77953 3012
rect 77987 3009 77999 3043
rect 77941 3003 77999 3009
rect 65576 2944 69980 2972
rect 65576 2932 65582 2944
rect 62298 2864 62304 2916
rect 62356 2904 62362 2916
rect 66257 2907 66315 2913
rect 66257 2904 66269 2907
rect 62356 2876 66269 2904
rect 62356 2864 62362 2876
rect 66257 2873 66269 2876
rect 66303 2904 66315 2907
rect 66346 2904 66352 2916
rect 66303 2876 66352 2904
rect 66303 2873 66315 2876
rect 66257 2867 66315 2873
rect 66346 2864 66352 2876
rect 66404 2864 66410 2916
rect 71317 2907 71375 2913
rect 71317 2904 71329 2907
rect 69676 2876 71329 2904
rect 2774 2836 2780 2848
rect 2735 2808 2780 2836
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 4982 2796 4988 2848
rect 5040 2836 5046 2848
rect 5169 2839 5227 2845
rect 5169 2836 5181 2839
rect 5040 2808 5181 2836
rect 5040 2796 5046 2808
rect 5169 2805 5181 2808
rect 5215 2805 5227 2839
rect 5718 2836 5724 2848
rect 5679 2808 5724 2836
rect 5169 2799 5227 2805
rect 5718 2796 5724 2808
rect 5776 2796 5782 2848
rect 6454 2836 6460 2848
rect 6415 2808 6460 2836
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 7190 2836 7196 2848
rect 7151 2808 7196 2836
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 7745 2839 7803 2845
rect 7745 2805 7757 2839
rect 7791 2836 7803 2839
rect 7926 2836 7932 2848
rect 7791 2808 7932 2836
rect 7791 2805 7803 2808
rect 7745 2799 7803 2805
rect 7926 2796 7932 2808
rect 7984 2796 7990 2848
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9677 2839 9735 2845
rect 9677 2836 9689 2839
rect 9456 2808 9689 2836
rect 9456 2796 9462 2808
rect 9677 2805 9689 2808
rect 9723 2805 9735 2839
rect 9677 2799 9735 2805
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10321 2839 10379 2845
rect 10321 2836 10333 2839
rect 10192 2808 10333 2836
rect 10192 2796 10198 2808
rect 10321 2805 10333 2808
rect 10367 2805 10379 2839
rect 10870 2836 10876 2848
rect 10831 2808 10876 2836
rect 10321 2799 10379 2805
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 11606 2836 11612 2848
rect 11567 2808 11612 2836
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 12342 2836 12348 2848
rect 12303 2808 12348 2836
rect 12342 2796 12348 2808
rect 12400 2796 12406 2848
rect 12897 2839 12955 2845
rect 12897 2805 12909 2839
rect 12943 2836 12955 2839
rect 13078 2836 13084 2848
rect 12943 2808 13084 2836
rect 12943 2805 12955 2808
rect 12897 2799 12955 2805
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 14737 2839 14795 2845
rect 14737 2836 14749 2839
rect 14608 2808 14749 2836
rect 14608 2796 14614 2808
rect 14737 2805 14749 2808
rect 14783 2805 14795 2839
rect 14737 2799 14795 2805
rect 15286 2796 15292 2848
rect 15344 2836 15350 2848
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 15344 2808 15485 2836
rect 15344 2796 15350 2808
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 16022 2836 16028 2848
rect 15983 2808 16028 2836
rect 15473 2799 15531 2805
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 16758 2836 16764 2848
rect 16719 2808 16764 2836
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 17494 2836 17500 2848
rect 17455 2808 17500 2836
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 18049 2839 18107 2845
rect 18049 2805 18061 2839
rect 18095 2836 18107 2839
rect 18230 2836 18236 2848
rect 18095 2808 18236 2836
rect 18095 2805 18107 2808
rect 18049 2799 18107 2805
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 19978 2836 19984 2848
rect 19939 2808 19984 2836
rect 19978 2796 19984 2808
rect 20036 2796 20042 2848
rect 20438 2796 20444 2848
rect 20496 2836 20502 2848
rect 20717 2839 20775 2845
rect 20717 2836 20729 2839
rect 20496 2808 20729 2836
rect 20496 2796 20502 2808
rect 20717 2805 20729 2808
rect 20763 2805 20775 2839
rect 21174 2836 21180 2848
rect 21135 2808 21180 2836
rect 20717 2799 20775 2805
rect 21174 2796 21180 2808
rect 21232 2796 21238 2848
rect 21910 2836 21916 2848
rect 21871 2808 21916 2836
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 22646 2836 22652 2848
rect 22607 2808 22652 2836
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 23201 2839 23259 2845
rect 23201 2805 23213 2839
rect 23247 2836 23259 2839
rect 23382 2836 23388 2848
rect 23247 2808 23388 2836
rect 23247 2805 23259 2808
rect 23201 2799 23259 2805
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 24854 2796 24860 2848
rect 24912 2836 24918 2848
rect 25041 2839 25099 2845
rect 25041 2836 25053 2839
rect 24912 2808 25053 2836
rect 24912 2796 24918 2808
rect 25041 2805 25053 2808
rect 25087 2805 25099 2839
rect 31478 2836 31484 2848
rect 31439 2808 31484 2836
rect 25041 2799 25099 2805
rect 31478 2796 31484 2808
rect 31536 2796 31542 2848
rect 35342 2836 35348 2848
rect 35303 2808 35348 2836
rect 35342 2796 35348 2808
rect 35400 2796 35406 2848
rect 35894 2796 35900 2848
rect 35952 2836 35958 2848
rect 36081 2839 36139 2845
rect 36081 2836 36093 2839
rect 35952 2808 36093 2836
rect 35952 2796 35958 2808
rect 36081 2805 36093 2808
rect 36127 2805 36139 2839
rect 36630 2836 36636 2848
rect 36591 2808 36636 2836
rect 36081 2799 36139 2805
rect 36630 2796 36636 2808
rect 36688 2796 36694 2848
rect 37366 2836 37372 2848
rect 37327 2808 37372 2836
rect 37366 2796 37372 2808
rect 37424 2796 37430 2848
rect 38102 2836 38108 2848
rect 38063 2808 38108 2836
rect 38102 2796 38108 2808
rect 38160 2796 38166 2848
rect 38657 2839 38715 2845
rect 38657 2805 38669 2839
rect 38703 2836 38715 2839
rect 38838 2836 38844 2848
rect 38703 2808 38844 2836
rect 38703 2805 38715 2808
rect 38657 2799 38715 2805
rect 38838 2796 38844 2808
rect 38896 2796 38902 2848
rect 41046 2836 41052 2848
rect 41007 2808 41052 2836
rect 41046 2796 41052 2808
rect 41104 2796 41110 2848
rect 42426 2836 42432 2848
rect 42387 2808 42432 2836
rect 42426 2796 42432 2808
rect 42484 2796 42490 2848
rect 42794 2796 42800 2848
rect 42852 2836 42858 2848
rect 42981 2839 43039 2845
rect 42981 2836 42993 2839
rect 42852 2808 42993 2836
rect 42852 2796 42858 2808
rect 42981 2805 42993 2808
rect 43027 2805 43039 2839
rect 42981 2799 43039 2805
rect 44726 2796 44732 2848
rect 44784 2836 44790 2848
rect 44821 2839 44879 2845
rect 44821 2836 44833 2839
rect 44784 2808 44833 2836
rect 44784 2796 44790 2808
rect 44821 2805 44833 2808
rect 44867 2805 44879 2839
rect 45646 2836 45652 2848
rect 45607 2808 45652 2836
rect 44821 2799 44879 2805
rect 45646 2796 45652 2808
rect 45704 2796 45710 2848
rect 46198 2796 46204 2848
rect 46256 2836 46262 2848
rect 46293 2839 46351 2845
rect 46293 2836 46305 2839
rect 46256 2808 46305 2836
rect 46256 2796 46262 2808
rect 46293 2805 46305 2808
rect 46339 2805 46351 2839
rect 47578 2836 47584 2848
rect 47539 2808 47584 2836
rect 46293 2799 46351 2805
rect 47578 2796 47584 2808
rect 47636 2796 47642 2848
rect 47670 2796 47676 2848
rect 47728 2836 47734 2848
rect 48133 2839 48191 2845
rect 48133 2836 48145 2839
rect 47728 2808 48145 2836
rect 47728 2796 47734 2808
rect 48133 2805 48145 2808
rect 48179 2836 48191 2839
rect 48406 2836 48412 2848
rect 48179 2808 48412 2836
rect 48179 2805 48191 2808
rect 48133 2799 48191 2805
rect 48406 2796 48412 2808
rect 48464 2796 48470 2848
rect 48774 2836 48780 2848
rect 48735 2808 48780 2836
rect 48774 2796 48780 2808
rect 48832 2796 48838 2848
rect 49142 2796 49148 2848
rect 49200 2836 49206 2848
rect 49329 2839 49387 2845
rect 49329 2836 49341 2839
rect 49200 2808 49341 2836
rect 49200 2796 49206 2808
rect 49329 2805 49341 2808
rect 49375 2805 49387 2839
rect 49329 2799 49387 2805
rect 54294 2796 54300 2848
rect 54352 2836 54358 2848
rect 54573 2839 54631 2845
rect 54573 2836 54585 2839
rect 54352 2808 54585 2836
rect 54352 2796 54358 2808
rect 54573 2805 54585 2808
rect 54619 2805 54631 2839
rect 54573 2799 54631 2805
rect 59446 2796 59452 2848
rect 59504 2836 59510 2848
rect 59633 2839 59691 2845
rect 59633 2836 59645 2839
rect 59504 2808 59645 2836
rect 59504 2796 59510 2808
rect 59633 2805 59645 2808
rect 59679 2805 59691 2839
rect 59633 2799 59691 2805
rect 59814 2796 59820 2848
rect 59872 2836 59878 2848
rect 63034 2836 63040 2848
rect 59872 2808 63040 2836
rect 59872 2796 59878 2808
rect 63034 2796 63040 2808
rect 63092 2796 63098 2848
rect 64598 2796 64604 2848
rect 64656 2836 64662 2848
rect 64877 2839 64935 2845
rect 64877 2836 64889 2839
rect 64656 2808 64889 2836
rect 64656 2796 64662 2808
rect 64877 2805 64889 2808
rect 64923 2805 64935 2839
rect 64877 2799 64935 2805
rect 66070 2796 66076 2848
rect 66128 2836 66134 2848
rect 69676 2836 69704 2876
rect 71317 2873 71329 2876
rect 71363 2904 71375 2907
rect 71498 2904 71504 2916
rect 71363 2876 71504 2904
rect 71363 2873 71375 2876
rect 71317 2867 71375 2873
rect 71498 2864 71504 2876
rect 71556 2864 71562 2916
rect 77110 2904 77116 2916
rect 77071 2876 77116 2904
rect 77110 2864 77116 2876
rect 77168 2904 77174 2916
rect 77386 2904 77392 2916
rect 77168 2876 77392 2904
rect 77168 2864 77174 2876
rect 77386 2864 77392 2876
rect 77444 2864 77450 2916
rect 66128 2808 69704 2836
rect 66128 2796 66134 2808
rect 69750 2796 69756 2848
rect 69808 2836 69814 2848
rect 70029 2839 70087 2845
rect 70029 2836 70041 2839
rect 69808 2808 70041 2836
rect 69808 2796 69814 2808
rect 70029 2805 70041 2808
rect 70075 2805 70087 2839
rect 73338 2836 73344 2848
rect 73299 2808 73344 2836
rect 70029 2799 70087 2805
rect 73338 2796 73344 2808
rect 73396 2796 73402 2848
rect 73890 2836 73896 2848
rect 73851 2808 73896 2836
rect 73890 2796 73896 2808
rect 73948 2796 73954 2848
rect 75730 2836 75736 2848
rect 75691 2808 75736 2836
rect 75730 2796 75736 2808
rect 75788 2796 75794 2848
rect 76374 2796 76380 2848
rect 76432 2836 76438 2848
rect 76469 2839 76527 2845
rect 76469 2836 76481 2839
rect 76432 2808 76481 2836
rect 76432 2796 76438 2808
rect 76469 2805 76481 2808
rect 76515 2805 76527 2839
rect 76469 2799 76527 2805
rect 1104 2746 78844 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 78844 2746
rect 1104 2672 78844 2694
rect 2314 2632 2320 2644
rect 2275 2604 2320 2632
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 4525 2635 4583 2641
rect 4525 2601 4537 2635
rect 4571 2632 4583 2635
rect 4614 2632 4620 2644
rect 4571 2604 4620 2632
rect 4571 2601 4583 2604
rect 4525 2595 4583 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 4764 2604 5181 2632
rect 4764 2592 4770 2604
rect 5169 2601 5181 2604
rect 5215 2601 5227 2635
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5169 2595 5227 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6178 2592 6184 2644
rect 6236 2632 6242 2644
rect 6733 2635 6791 2641
rect 6733 2632 6745 2635
rect 6236 2604 6745 2632
rect 6236 2592 6242 2604
rect 6733 2601 6745 2604
rect 6779 2601 6791 2635
rect 6733 2595 6791 2601
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 6972 2604 7481 2632
rect 6972 2592 6978 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 8202 2632 8208 2644
rect 8163 2604 8208 2632
rect 7469 2595 7527 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10778 2632 10784 2644
rect 10739 2604 10784 2632
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 11882 2632 11888 2644
rect 11843 2604 11888 2632
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12618 2632 12624 2644
rect 12579 2604 12624 2632
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 13354 2632 13360 2644
rect 13315 2604 13360 2632
rect 13354 2592 13360 2604
rect 13412 2592 13418 2644
rect 14458 2632 14464 2644
rect 14419 2604 14464 2632
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 15930 2632 15936 2644
rect 15891 2604 15936 2632
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 17034 2632 17040 2644
rect 16995 2604 17040 2632
rect 17034 2592 17040 2604
rect 17092 2592 17098 2644
rect 17770 2632 17776 2644
rect 17731 2604 17776 2632
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 18506 2632 18512 2644
rect 18467 2604 18512 2632
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 20346 2632 20352 2644
rect 20307 2604 20352 2632
rect 20346 2592 20352 2604
rect 20404 2592 20410 2644
rect 22922 2632 22928 2644
rect 22883 2604 22928 2632
rect 22922 2592 22928 2604
rect 22980 2592 22986 2644
rect 23658 2632 23664 2644
rect 23619 2604 23664 2632
rect 23658 2592 23664 2604
rect 23716 2592 23722 2644
rect 24946 2632 24952 2644
rect 24907 2604 24952 2632
rect 24946 2592 24952 2604
rect 25004 2592 25010 2644
rect 33962 2632 33968 2644
rect 33923 2604 33968 2632
rect 33962 2592 33968 2604
rect 34020 2592 34026 2644
rect 35805 2635 35863 2641
rect 35805 2601 35817 2635
rect 35851 2632 35863 2635
rect 36262 2632 36268 2644
rect 35851 2604 36268 2632
rect 35851 2601 35863 2604
rect 35805 2595 35863 2601
rect 36262 2592 36268 2604
rect 36320 2592 36326 2644
rect 36538 2632 36544 2644
rect 36499 2604 36544 2632
rect 36538 2592 36544 2604
rect 36596 2592 36602 2644
rect 37642 2632 37648 2644
rect 37603 2604 37648 2632
rect 37642 2592 37648 2604
rect 37700 2592 37706 2644
rect 38378 2632 38384 2644
rect 38339 2604 38384 2632
rect 38378 2592 38384 2604
rect 38436 2592 38442 2644
rect 39114 2632 39120 2644
rect 39075 2604 39120 2632
rect 39114 2592 39120 2604
rect 39172 2592 39178 2644
rect 40586 2632 40592 2644
rect 40547 2604 40592 2632
rect 40586 2592 40592 2604
rect 40644 2592 40650 2644
rect 42610 2632 42616 2644
rect 42571 2604 42616 2632
rect 42610 2592 42616 2604
rect 42668 2592 42674 2644
rect 43346 2632 43352 2644
rect 43307 2604 43352 2632
rect 43346 2592 43352 2604
rect 43404 2592 43410 2644
rect 45186 2632 45192 2644
rect 45147 2604 45192 2632
rect 45186 2592 45192 2604
rect 45244 2592 45250 2644
rect 45922 2632 45928 2644
rect 45883 2604 45928 2632
rect 45922 2592 45928 2604
rect 45980 2592 45986 2644
rect 46658 2632 46664 2644
rect 46619 2604 46664 2632
rect 46658 2592 46664 2604
rect 46716 2592 46722 2644
rect 47762 2632 47768 2644
rect 47723 2604 47768 2632
rect 47762 2592 47768 2604
rect 47820 2592 47826 2644
rect 49234 2632 49240 2644
rect 49195 2604 49240 2632
rect 49234 2592 49240 2604
rect 49292 2592 49298 2644
rect 73522 2632 73528 2644
rect 73483 2604 73528 2632
rect 73522 2592 73528 2604
rect 73580 2592 73586 2644
rect 74258 2632 74264 2644
rect 74219 2604 74264 2632
rect 74258 2592 74264 2604
rect 74316 2592 74322 2644
rect 74994 2632 75000 2644
rect 74955 2604 75000 2632
rect 74994 2592 75000 2604
rect 75052 2592 75058 2644
rect 76101 2635 76159 2641
rect 76101 2601 76113 2635
rect 76147 2632 76159 2635
rect 76282 2632 76288 2644
rect 76147 2604 76288 2632
rect 76147 2601 76159 2604
rect 76101 2595 76159 2601
rect 76282 2592 76288 2604
rect 76340 2592 76346 2644
rect 15102 2564 15108 2576
rect 15063 2536 15108 2564
rect 15102 2524 15108 2536
rect 15160 2524 15166 2576
rect 19426 2524 19432 2576
rect 19484 2564 19490 2576
rect 19521 2567 19579 2573
rect 19521 2564 19533 2567
rect 19484 2536 19533 2564
rect 19484 2524 19490 2536
rect 19521 2533 19533 2536
rect 19567 2533 19579 2567
rect 19521 2527 19579 2533
rect 22281 2567 22339 2573
rect 22281 2533 22293 2567
rect 22327 2564 22339 2567
rect 26326 2564 26332 2576
rect 22327 2536 26332 2564
rect 22327 2533 22339 2536
rect 22281 2527 22339 2533
rect 26326 2524 26332 2536
rect 26384 2524 26390 2576
rect 34790 2524 34796 2576
rect 34848 2564 34854 2576
rect 34977 2567 35035 2573
rect 34977 2564 34989 2567
rect 34848 2536 34989 2564
rect 34848 2524 34854 2536
rect 34977 2533 34989 2536
rect 35023 2533 35035 2567
rect 41414 2564 41420 2576
rect 41375 2536 41420 2564
rect 34977 2527 35035 2533
rect 41414 2524 41420 2536
rect 41472 2524 41478 2576
rect 44174 2564 44180 2576
rect 44135 2536 44180 2564
rect 44174 2524 44180 2536
rect 44232 2524 44238 2576
rect 47486 2524 47492 2576
rect 47544 2564 47550 2576
rect 48593 2567 48651 2573
rect 48593 2564 48605 2567
rect 47544 2536 48605 2564
rect 47544 2524 47550 2536
rect 48593 2533 48605 2536
rect 48639 2533 48651 2567
rect 48593 2527 48651 2533
rect 52822 2524 52828 2576
rect 52880 2564 52886 2576
rect 53561 2567 53619 2573
rect 53561 2564 53573 2567
rect 52880 2536 53573 2564
rect 52880 2524 52886 2536
rect 53561 2533 53573 2536
rect 53607 2533 53619 2567
rect 53561 2527 53619 2533
rect 57974 2524 57980 2576
rect 58032 2564 58038 2576
rect 58805 2567 58863 2573
rect 58805 2564 58817 2567
rect 58032 2536 58817 2564
rect 58032 2524 58038 2536
rect 58805 2533 58817 2536
rect 58851 2533 58863 2567
rect 58805 2527 58863 2533
rect 63862 2524 63868 2576
rect 63920 2564 63926 2576
rect 64693 2567 64751 2573
rect 64693 2564 64705 2567
rect 63920 2536 64705 2564
rect 63920 2524 63926 2536
rect 64693 2533 64705 2536
rect 64739 2533 64751 2567
rect 64693 2527 64751 2533
rect 69014 2524 69020 2576
rect 69072 2564 69078 2576
rect 69845 2567 69903 2573
rect 69845 2564 69857 2567
rect 69072 2536 69857 2564
rect 69072 2524 69078 2536
rect 69845 2533 69857 2536
rect 69891 2533 69903 2567
rect 69845 2527 69903 2533
rect 26142 2496 26148 2508
rect 26103 2468 26148 2496
rect 26142 2456 26148 2468
rect 26200 2456 26206 2508
rect 28718 2496 28724 2508
rect 28679 2468 28724 2496
rect 28718 2456 28724 2468
rect 28776 2456 28782 2508
rect 31018 2496 31024 2508
rect 30979 2468 31024 2496
rect 31018 2456 31024 2468
rect 31076 2456 31082 2508
rect 31938 2456 31944 2508
rect 31996 2496 32002 2508
rect 32401 2499 32459 2505
rect 32401 2496 32413 2499
rect 31996 2468 32413 2496
rect 31996 2456 32002 2468
rect 32401 2465 32413 2468
rect 32447 2465 32459 2499
rect 32401 2459 32459 2465
rect 53282 2456 53288 2508
rect 53340 2496 53346 2508
rect 53340 2468 54248 2496
rect 53340 2456 53346 2468
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 2038 2428 2044 2440
rect 1719 2400 2044 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2038 2388 2044 2400
rect 2096 2428 2102 2440
rect 2133 2431 2191 2437
rect 2133 2428 2145 2431
rect 2096 2400 2145 2428
rect 2096 2388 2102 2400
rect 2133 2397 2145 2400
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 2869 2431 2927 2437
rect 2869 2428 2881 2431
rect 2832 2400 2881 2428
rect 2832 2388 2838 2400
rect 2869 2397 2881 2400
rect 2915 2397 2927 2431
rect 2869 2391 2927 2397
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 4246 2428 4252 2440
rect 3927 2400 4252 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 4246 2388 4252 2400
rect 4304 2428 4310 2440
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4304 2400 4353 2428
rect 4304 2388 4310 2400
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 4982 2428 4988 2440
rect 4943 2400 4988 2428
rect 4341 2391 4399 2397
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 5776 2400 5825 2428
rect 5776 2388 5782 2400
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6512 2400 6561 2428
rect 6512 2388 6518 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 7248 2400 7297 2428
rect 7248 2388 7254 2400
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 8021 2431 8079 2437
rect 8021 2428 8033 2431
rect 7984 2400 8033 2428
rect 7984 2388 7990 2400
rect 8021 2397 8033 2400
rect 8067 2397 8079 2431
rect 9398 2428 9404 2440
rect 9359 2400 9404 2428
rect 8021 2391 8079 2397
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 10134 2388 10140 2440
rect 10192 2428 10198 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 10192 2400 10241 2428
rect 10192 2388 10198 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10870 2388 10876 2440
rect 10928 2428 10934 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10928 2400 10977 2428
rect 10928 2388 10934 2400
rect 10965 2397 10977 2400
rect 11011 2397 11023 2431
rect 22094 2428 22100 2440
rect 22055 2400 22100 2428
rect 10965 2391 11023 2397
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23532 2400 23581 2428
rect 23532 2388 23538 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 23569 2391 23627 2397
rect 26326 2388 26332 2440
rect 26384 2428 26390 2440
rect 26421 2431 26479 2437
rect 26421 2428 26433 2431
rect 26384 2400 26433 2428
rect 26384 2388 26390 2400
rect 26421 2397 26433 2400
rect 26467 2428 26479 2431
rect 26973 2431 27031 2437
rect 26973 2428 26985 2431
rect 26467 2400 26985 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 26973 2397 26985 2400
rect 27019 2397 27031 2431
rect 26973 2391 27031 2397
rect 28534 2388 28540 2440
rect 28592 2428 28598 2440
rect 28997 2431 29055 2437
rect 28997 2428 29009 2431
rect 28592 2400 29009 2428
rect 28592 2388 28598 2400
rect 28997 2397 29009 2400
rect 29043 2428 29055 2431
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29043 2400 29561 2428
rect 29043 2397 29055 2400
rect 28997 2391 29055 2397
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 30285 2431 30343 2437
rect 30285 2397 30297 2431
rect 30331 2428 30343 2431
rect 30742 2428 30748 2440
rect 30331 2400 30748 2428
rect 30331 2397 30343 2400
rect 30285 2391 30343 2397
rect 30742 2388 30748 2400
rect 30800 2388 30806 2440
rect 31478 2388 31484 2440
rect 31536 2428 31542 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31536 2400 32137 2428
rect 31536 2388 31542 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 45646 2388 45652 2440
rect 45704 2428 45710 2440
rect 45833 2431 45891 2437
rect 45833 2428 45845 2431
rect 45704 2400 45845 2428
rect 45704 2388 45710 2400
rect 45833 2397 45845 2400
rect 45879 2397 45891 2431
rect 48406 2428 48412 2440
rect 48367 2400 48412 2428
rect 45833 2391 45891 2397
rect 48406 2388 48412 2400
rect 48464 2388 48470 2440
rect 50433 2431 50491 2437
rect 50433 2397 50445 2431
rect 50479 2428 50491 2431
rect 50614 2428 50620 2440
rect 50479 2400 50620 2428
rect 50479 2397 50491 2400
rect 50433 2391 50491 2397
rect 50614 2388 50620 2400
rect 50672 2388 50678 2440
rect 51169 2431 51227 2437
rect 51169 2397 51181 2431
rect 51215 2428 51227 2431
rect 51258 2428 51264 2440
rect 51215 2400 51264 2428
rect 51215 2397 51227 2400
rect 51169 2391 51227 2397
rect 51258 2388 51264 2400
rect 51316 2388 51322 2440
rect 51810 2388 51816 2440
rect 51868 2428 51874 2440
rect 51905 2431 51963 2437
rect 51905 2428 51917 2431
rect 51868 2400 51917 2428
rect 51868 2388 51874 2400
rect 51905 2397 51917 2400
rect 51951 2397 51963 2431
rect 51905 2391 51963 2397
rect 52362 2388 52368 2440
rect 52420 2428 52426 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52420 2400 52745 2428
rect 52420 2388 52426 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 53745 2431 53803 2437
rect 53745 2397 53757 2431
rect 53791 2428 53803 2431
rect 53834 2428 53840 2440
rect 53791 2400 53840 2428
rect 53791 2397 53803 2400
rect 53745 2391 53803 2397
rect 53834 2388 53840 2400
rect 53892 2388 53898 2440
rect 54220 2437 54248 2468
rect 60550 2456 60556 2508
rect 60608 2496 60614 2508
rect 60608 2468 61516 2496
rect 60608 2456 60614 2468
rect 54205 2431 54263 2437
rect 54205 2397 54217 2431
rect 54251 2397 54263 2431
rect 54205 2391 54263 2397
rect 55309 2431 55367 2437
rect 55309 2397 55321 2431
rect 55355 2428 55367 2431
rect 55398 2428 55404 2440
rect 55355 2400 55404 2428
rect 55355 2397 55367 2400
rect 55309 2391 55367 2397
rect 55398 2388 55404 2400
rect 55456 2388 55462 2440
rect 56321 2431 56379 2437
rect 56321 2397 56333 2431
rect 56367 2428 56379 2431
rect 56594 2428 56600 2440
rect 56367 2400 56600 2428
rect 56367 2397 56379 2400
rect 56321 2391 56379 2397
rect 56594 2388 56600 2400
rect 56652 2388 56658 2440
rect 57057 2431 57115 2437
rect 57057 2397 57069 2431
rect 57103 2428 57115 2431
rect 57146 2428 57152 2440
rect 57103 2400 57152 2428
rect 57103 2397 57115 2400
rect 57057 2391 57115 2397
rect 57146 2388 57152 2400
rect 57204 2388 57210 2440
rect 57882 2428 57888 2440
rect 57843 2400 57888 2428
rect 57882 2388 57888 2400
rect 57940 2388 57946 2440
rect 58434 2388 58440 2440
rect 58492 2428 58498 2440
rect 58621 2431 58679 2437
rect 58621 2428 58633 2431
rect 58492 2400 58633 2428
rect 58492 2388 58498 2400
rect 58621 2397 58633 2400
rect 58667 2397 58679 2431
rect 58621 2391 58679 2397
rect 58986 2388 58992 2440
rect 59044 2428 59050 2440
rect 59357 2431 59415 2437
rect 59357 2428 59369 2431
rect 59044 2400 59369 2428
rect 59044 2388 59050 2400
rect 59357 2397 59369 2400
rect 59403 2397 59415 2431
rect 59357 2391 59415 2397
rect 60642 2388 60648 2440
rect 60700 2428 60706 2440
rect 61488 2437 61516 2468
rect 66162 2456 66168 2508
rect 66220 2496 66226 2508
rect 66220 2468 67128 2496
rect 66220 2456 66226 2468
rect 60737 2431 60795 2437
rect 60737 2428 60749 2431
rect 60700 2400 60749 2428
rect 60700 2388 60706 2400
rect 60737 2397 60749 2400
rect 60783 2397 60795 2431
rect 60737 2391 60795 2397
rect 61473 2431 61531 2437
rect 61473 2397 61485 2431
rect 61519 2397 61531 2431
rect 61930 2428 61936 2440
rect 61891 2400 61936 2428
rect 61473 2391 61531 2397
rect 61930 2388 61936 2400
rect 61988 2388 61994 2440
rect 63034 2428 63040 2440
rect 62995 2400 63040 2428
rect 63034 2388 63040 2400
rect 63092 2388 63098 2440
rect 63402 2388 63408 2440
rect 63460 2428 63466 2440
rect 63773 2431 63831 2437
rect 63773 2428 63785 2431
rect 63460 2400 63785 2428
rect 63460 2388 63466 2400
rect 63773 2397 63785 2400
rect 63819 2397 63831 2431
rect 63773 2391 63831 2397
rect 64322 2388 64328 2440
rect 64380 2428 64386 2440
rect 64509 2431 64567 2437
rect 64509 2428 64521 2431
rect 64380 2400 64521 2428
rect 64380 2388 64386 2400
rect 64509 2397 64521 2400
rect 64555 2397 64567 2431
rect 64509 2391 64567 2397
rect 65426 2388 65432 2440
rect 65484 2428 65490 2440
rect 65613 2431 65671 2437
rect 65613 2428 65625 2431
rect 65484 2400 65625 2428
rect 65484 2388 65490 2400
rect 65613 2397 65625 2400
rect 65659 2397 65671 2431
rect 66346 2428 66352 2440
rect 66307 2400 66352 2428
rect 65613 2391 65671 2397
rect 66346 2388 66352 2400
rect 66404 2388 66410 2440
rect 67100 2437 67128 2468
rect 67085 2431 67143 2437
rect 67085 2397 67097 2431
rect 67131 2397 67143 2431
rect 68186 2428 68192 2440
rect 68147 2400 68192 2428
rect 67085 2391 67143 2397
rect 68186 2388 68192 2400
rect 68244 2388 68250 2440
rect 68922 2428 68928 2440
rect 68883 2400 68928 2428
rect 68922 2388 68928 2400
rect 68980 2388 68986 2440
rect 69658 2428 69664 2440
rect 69619 2400 69664 2428
rect 69658 2388 69664 2400
rect 69716 2388 69722 2440
rect 70578 2388 70584 2440
rect 70636 2428 70642 2440
rect 70765 2431 70823 2437
rect 70765 2428 70777 2431
rect 70636 2400 70777 2428
rect 70636 2388 70642 2400
rect 70765 2397 70777 2400
rect 70811 2397 70823 2431
rect 71498 2428 71504 2440
rect 71459 2400 71504 2428
rect 70765 2391 70823 2397
rect 71498 2388 71504 2400
rect 71556 2388 71562 2440
rect 72050 2388 72056 2440
rect 72108 2428 72114 2440
rect 72237 2431 72295 2437
rect 72237 2428 72249 2431
rect 72108 2400 72249 2428
rect 72108 2388 72114 2400
rect 72237 2397 72249 2400
rect 72283 2397 72295 2431
rect 72237 2391 72295 2397
rect 72694 2388 72700 2440
rect 72752 2428 72758 2440
rect 73338 2428 73344 2440
rect 72752 2400 73344 2428
rect 72752 2388 72758 2400
rect 73338 2388 73344 2400
rect 73396 2388 73402 2440
rect 73430 2388 73436 2440
rect 73488 2428 73494 2440
rect 73890 2428 73896 2440
rect 73488 2400 73896 2428
rect 73488 2388 73494 2400
rect 73890 2388 73896 2400
rect 73948 2428 73954 2440
rect 74077 2431 74135 2437
rect 74077 2428 74089 2431
rect 73948 2400 74089 2428
rect 73948 2388 73954 2400
rect 74077 2397 74089 2400
rect 74123 2397 74135 2431
rect 74077 2391 74135 2397
rect 74718 2388 74724 2440
rect 74776 2428 74782 2440
rect 74813 2431 74871 2437
rect 74813 2428 74825 2431
rect 74776 2400 74825 2428
rect 74776 2388 74782 2400
rect 74813 2397 74825 2400
rect 74859 2397 74871 2431
rect 75914 2428 75920 2440
rect 75875 2400 75920 2428
rect 74813 2391 74871 2397
rect 75914 2388 75920 2400
rect 75972 2388 75978 2440
rect 76374 2388 76380 2440
rect 76432 2428 76438 2440
rect 76653 2431 76711 2437
rect 76653 2428 76665 2431
rect 76432 2400 76665 2428
rect 76432 2388 76438 2400
rect 76653 2397 76665 2400
rect 76699 2397 76711 2431
rect 77386 2428 77392 2440
rect 77347 2400 77392 2428
rect 76653 2391 76711 2397
rect 77386 2388 77392 2400
rect 77444 2388 77450 2440
rect 11606 2320 11612 2372
rect 11664 2360 11670 2372
rect 11793 2363 11851 2369
rect 11793 2360 11805 2363
rect 11664 2332 11805 2360
rect 11664 2320 11670 2332
rect 11793 2329 11805 2332
rect 11839 2329 11851 2363
rect 11793 2323 11851 2329
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 12529 2363 12587 2369
rect 12529 2360 12541 2363
rect 12492 2332 12541 2360
rect 12492 2320 12498 2332
rect 12529 2329 12541 2332
rect 12575 2329 12587 2363
rect 12529 2323 12587 2329
rect 13078 2320 13084 2372
rect 13136 2360 13142 2372
rect 13265 2363 13323 2369
rect 13265 2360 13277 2363
rect 13136 2332 13277 2360
rect 13136 2320 13142 2332
rect 13265 2329 13277 2332
rect 13311 2329 13323 2363
rect 14550 2360 14556 2372
rect 14511 2332 14556 2360
rect 13265 2323 13323 2329
rect 14550 2320 14556 2332
rect 14608 2320 14614 2372
rect 15286 2360 15292 2372
rect 15247 2332 15292 2360
rect 15286 2320 15292 2332
rect 15344 2320 15350 2372
rect 16022 2360 16028 2372
rect 15983 2332 16028 2360
rect 16022 2320 16028 2332
rect 16080 2320 16086 2372
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 16945 2363 17003 2369
rect 16945 2360 16957 2363
rect 16816 2332 16957 2360
rect 16816 2320 16822 2332
rect 16945 2329 16957 2332
rect 16991 2329 17003 2363
rect 16945 2323 17003 2329
rect 17494 2320 17500 2372
rect 17552 2360 17558 2372
rect 17681 2363 17739 2369
rect 17681 2360 17693 2363
rect 17552 2332 17693 2360
rect 17552 2320 17558 2332
rect 17681 2329 17693 2332
rect 17727 2329 17739 2363
rect 17681 2323 17739 2329
rect 18230 2320 18236 2372
rect 18288 2360 18294 2372
rect 18417 2363 18475 2369
rect 18417 2360 18429 2363
rect 18288 2332 18429 2360
rect 18288 2320 18294 2332
rect 18417 2329 18429 2332
rect 18463 2329 18475 2363
rect 18417 2323 18475 2329
rect 19705 2363 19763 2369
rect 19705 2329 19717 2363
rect 19751 2360 19763 2363
rect 19978 2360 19984 2372
rect 19751 2332 19984 2360
rect 19751 2329 19763 2332
rect 19705 2323 19763 2329
rect 19978 2320 19984 2332
rect 20036 2320 20042 2372
rect 20438 2360 20444 2372
rect 20399 2332 20444 2360
rect 20438 2320 20444 2332
rect 20496 2320 20502 2372
rect 21174 2360 21180 2372
rect 21135 2332 21180 2360
rect 21174 2320 21180 2332
rect 21232 2320 21238 2372
rect 22112 2332 22600 2360
rect 21085 2295 21143 2301
rect 21085 2261 21097 2295
rect 21131 2292 21143 2295
rect 22112 2292 22140 2332
rect 21131 2264 22140 2292
rect 22572 2292 22600 2332
rect 22646 2320 22652 2372
rect 22704 2360 22710 2372
rect 22833 2363 22891 2369
rect 22833 2360 22845 2363
rect 22704 2332 22845 2360
rect 22704 2320 22710 2332
rect 22833 2329 22845 2332
rect 22879 2329 22891 2363
rect 22833 2323 22891 2329
rect 24854 2320 24860 2372
rect 24912 2360 24918 2372
rect 25041 2363 25099 2369
rect 25041 2360 25053 2363
rect 24912 2332 25053 2360
rect 24912 2320 24918 2332
rect 25041 2329 25053 2332
rect 25087 2329 25099 2363
rect 25041 2323 25099 2329
rect 33686 2320 33692 2372
rect 33744 2360 33750 2372
rect 33873 2363 33931 2369
rect 33873 2360 33885 2363
rect 33744 2332 33885 2360
rect 33744 2320 33750 2332
rect 33873 2329 33885 2332
rect 33919 2329 33931 2363
rect 35158 2360 35164 2372
rect 35119 2332 35164 2360
rect 33873 2323 33931 2329
rect 35158 2320 35164 2332
rect 35216 2320 35222 2372
rect 35894 2320 35900 2372
rect 35952 2360 35958 2372
rect 36630 2360 36636 2372
rect 35952 2332 35997 2360
rect 36591 2332 36636 2360
rect 35952 2320 35958 2332
rect 36630 2320 36636 2332
rect 36688 2320 36694 2372
rect 37366 2320 37372 2372
rect 37424 2360 37430 2372
rect 37553 2363 37611 2369
rect 37553 2360 37565 2363
rect 37424 2332 37565 2360
rect 37424 2320 37430 2332
rect 37553 2329 37565 2332
rect 37599 2329 37611 2363
rect 37553 2323 37611 2329
rect 38102 2320 38108 2372
rect 38160 2360 38166 2372
rect 38289 2363 38347 2369
rect 38289 2360 38301 2363
rect 38160 2332 38301 2360
rect 38160 2320 38166 2332
rect 38289 2329 38301 2332
rect 38335 2329 38347 2363
rect 38289 2323 38347 2329
rect 38838 2320 38844 2372
rect 38896 2360 38902 2372
rect 39025 2363 39083 2369
rect 39025 2360 39037 2363
rect 38896 2332 39037 2360
rect 38896 2320 38902 2332
rect 39025 2329 39037 2332
rect 39071 2329 39083 2363
rect 39025 2323 39083 2329
rect 39945 2363 40003 2369
rect 39945 2329 39957 2363
rect 39991 2360 40003 2363
rect 40310 2360 40316 2372
rect 39991 2332 40316 2360
rect 39991 2329 40003 2332
rect 39945 2323 40003 2329
rect 40310 2320 40316 2332
rect 40368 2360 40374 2372
rect 40497 2363 40555 2369
rect 40497 2360 40509 2363
rect 40368 2332 40509 2360
rect 40368 2320 40374 2332
rect 40497 2329 40509 2332
rect 40543 2329 40555 2363
rect 40497 2323 40555 2329
rect 41046 2320 41052 2372
rect 41104 2360 41110 2372
rect 41233 2363 41291 2369
rect 41233 2360 41245 2363
rect 41104 2332 41245 2360
rect 41104 2320 41110 2332
rect 41233 2329 41245 2332
rect 41279 2329 41291 2363
rect 41233 2323 41291 2329
rect 41782 2320 41788 2372
rect 41840 2360 41846 2372
rect 42426 2360 42432 2372
rect 41840 2332 42432 2360
rect 41840 2320 41846 2332
rect 42426 2320 42432 2332
rect 42484 2360 42490 2372
rect 42521 2363 42579 2369
rect 42521 2360 42533 2363
rect 42484 2332 42533 2360
rect 42484 2320 42490 2332
rect 42521 2329 42533 2332
rect 42567 2329 42579 2363
rect 42521 2323 42579 2329
rect 42794 2320 42800 2372
rect 42852 2360 42858 2372
rect 43257 2363 43315 2369
rect 43257 2360 43269 2363
rect 42852 2332 43269 2360
rect 42852 2320 42858 2332
rect 43257 2329 43269 2332
rect 43303 2329 43315 2363
rect 43257 2323 43315 2329
rect 43346 2320 43352 2372
rect 43404 2360 43410 2372
rect 43714 2360 43720 2372
rect 43404 2332 43720 2360
rect 43404 2320 43410 2332
rect 43714 2320 43720 2332
rect 43772 2360 43778 2372
rect 43993 2363 44051 2369
rect 43993 2360 44005 2363
rect 43772 2332 44005 2360
rect 43772 2320 43778 2332
rect 43993 2329 44005 2332
rect 44039 2329 44051 2363
rect 43993 2323 44051 2329
rect 44726 2320 44732 2372
rect 44784 2360 44790 2372
rect 45097 2363 45155 2369
rect 45097 2360 45109 2363
rect 44784 2332 45109 2360
rect 44784 2320 44790 2332
rect 45097 2329 45109 2332
rect 45143 2329 45155 2363
rect 45097 2323 45155 2329
rect 46198 2320 46204 2372
rect 46256 2360 46262 2372
rect 46569 2363 46627 2369
rect 46569 2360 46581 2363
rect 46256 2332 46581 2360
rect 46256 2320 46262 2332
rect 46569 2329 46581 2332
rect 46615 2329 46627 2363
rect 46569 2323 46627 2329
rect 46934 2320 46940 2372
rect 46992 2360 46998 2372
rect 47578 2360 47584 2372
rect 46992 2332 47584 2360
rect 46992 2320 46998 2332
rect 47578 2320 47584 2332
rect 47636 2360 47642 2372
rect 47673 2363 47731 2369
rect 47673 2360 47685 2363
rect 47636 2332 47685 2360
rect 47636 2320 47642 2332
rect 47673 2329 47685 2332
rect 47719 2329 47731 2363
rect 48774 2360 48780 2372
rect 47673 2323 47731 2329
rect 48424 2332 48780 2360
rect 48424 2304 48452 2332
rect 48774 2320 48780 2332
rect 48832 2360 48838 2372
rect 49145 2363 49203 2369
rect 49145 2360 49157 2363
rect 48832 2332 49157 2360
rect 48832 2320 48838 2332
rect 49145 2329 49157 2332
rect 49191 2329 49203 2363
rect 49145 2323 49203 2329
rect 67358 2320 67364 2372
rect 67416 2360 67422 2372
rect 67416 2332 74534 2360
rect 67416 2320 67422 2332
rect 26510 2292 26516 2304
rect 22572 2264 26516 2292
rect 21131 2261 21143 2264
rect 21085 2255 21143 2261
rect 26510 2252 26516 2264
rect 26568 2252 26574 2304
rect 48406 2252 48412 2304
rect 48464 2252 48470 2304
rect 49878 2252 49884 2304
rect 49936 2292 49942 2304
rect 50249 2295 50307 2301
rect 50249 2292 50261 2295
rect 49936 2264 50261 2292
rect 49936 2252 49942 2264
rect 50249 2261 50261 2264
rect 50295 2261 50307 2295
rect 50249 2255 50307 2261
rect 50614 2252 50620 2304
rect 50672 2292 50678 2304
rect 50985 2295 51043 2301
rect 50985 2292 50997 2295
rect 50672 2264 50997 2292
rect 50672 2252 50678 2264
rect 50985 2261 50997 2264
rect 51031 2261 51043 2295
rect 50985 2255 51043 2261
rect 51350 2252 51356 2304
rect 51408 2292 51414 2304
rect 51721 2295 51779 2301
rect 51721 2292 51733 2295
rect 51408 2264 51733 2292
rect 51408 2252 51414 2264
rect 51721 2261 51733 2264
rect 51767 2261 51779 2295
rect 51721 2255 51779 2261
rect 52086 2252 52092 2304
rect 52144 2292 52150 2304
rect 52917 2295 52975 2301
rect 52917 2292 52929 2295
rect 52144 2264 52929 2292
rect 52144 2252 52150 2264
rect 52917 2261 52929 2264
rect 52963 2261 52975 2295
rect 52917 2255 52975 2261
rect 53558 2252 53564 2304
rect 53616 2292 53622 2304
rect 54389 2295 54447 2301
rect 54389 2292 54401 2295
rect 53616 2264 54401 2292
rect 53616 2252 53622 2264
rect 54389 2261 54401 2264
rect 54435 2261 54447 2295
rect 54389 2255 54447 2261
rect 55030 2252 55036 2304
rect 55088 2292 55094 2304
rect 55493 2295 55551 2301
rect 55493 2292 55505 2295
rect 55088 2264 55505 2292
rect 55088 2252 55094 2264
rect 55493 2261 55505 2264
rect 55539 2261 55551 2295
rect 55493 2255 55551 2261
rect 55766 2252 55772 2304
rect 55824 2292 55830 2304
rect 56137 2295 56195 2301
rect 56137 2292 56149 2295
rect 55824 2264 56149 2292
rect 55824 2252 55830 2264
rect 56137 2261 56149 2264
rect 56183 2261 56195 2295
rect 56137 2255 56195 2261
rect 56502 2252 56508 2304
rect 56560 2292 56566 2304
rect 56873 2295 56931 2301
rect 56873 2292 56885 2295
rect 56560 2264 56885 2292
rect 56560 2252 56566 2264
rect 56873 2261 56885 2264
rect 56919 2261 56931 2295
rect 56873 2255 56931 2261
rect 57238 2252 57244 2304
rect 57296 2292 57302 2304
rect 58069 2295 58127 2301
rect 58069 2292 58081 2295
rect 57296 2264 58081 2292
rect 57296 2252 57302 2264
rect 58069 2261 58081 2264
rect 58115 2261 58127 2295
rect 58069 2255 58127 2261
rect 58710 2252 58716 2304
rect 58768 2292 58774 2304
rect 59541 2295 59599 2301
rect 59541 2292 59553 2295
rect 58768 2264 59553 2292
rect 58768 2252 58774 2264
rect 59541 2261 59553 2264
rect 59587 2261 59599 2295
rect 59541 2255 59599 2261
rect 60182 2252 60188 2304
rect 60240 2292 60246 2304
rect 60553 2295 60611 2301
rect 60553 2292 60565 2295
rect 60240 2264 60565 2292
rect 60240 2252 60246 2264
rect 60553 2261 60565 2264
rect 60599 2261 60611 2295
rect 60553 2255 60611 2261
rect 60918 2252 60924 2304
rect 60976 2292 60982 2304
rect 61289 2295 61347 2301
rect 61289 2292 61301 2295
rect 60976 2264 61301 2292
rect 60976 2252 60982 2264
rect 61289 2261 61301 2264
rect 61335 2261 61347 2295
rect 61289 2255 61347 2261
rect 61654 2252 61660 2304
rect 61712 2292 61718 2304
rect 62117 2295 62175 2301
rect 62117 2292 62129 2295
rect 61712 2264 62129 2292
rect 61712 2252 61718 2264
rect 62117 2261 62129 2264
rect 62163 2261 62175 2295
rect 62117 2255 62175 2261
rect 62390 2252 62396 2304
rect 62448 2292 62454 2304
rect 63221 2295 63279 2301
rect 63221 2292 63233 2295
rect 62448 2264 63233 2292
rect 62448 2252 62454 2264
rect 63221 2261 63233 2264
rect 63267 2261 63279 2295
rect 63221 2255 63279 2261
rect 63402 2252 63408 2304
rect 63460 2292 63466 2304
rect 63957 2295 64015 2301
rect 63957 2292 63969 2295
rect 63460 2264 63969 2292
rect 63460 2252 63466 2264
rect 63957 2261 63969 2264
rect 64003 2261 64015 2295
rect 63957 2255 64015 2261
rect 65334 2252 65340 2304
rect 65392 2292 65398 2304
rect 65797 2295 65855 2301
rect 65797 2292 65809 2295
rect 65392 2264 65809 2292
rect 65392 2252 65398 2264
rect 65797 2261 65809 2264
rect 65843 2261 65855 2295
rect 65797 2255 65855 2261
rect 66070 2252 66076 2304
rect 66128 2292 66134 2304
rect 66533 2295 66591 2301
rect 66533 2292 66545 2295
rect 66128 2264 66545 2292
rect 66128 2252 66134 2264
rect 66533 2261 66545 2264
rect 66579 2261 66591 2295
rect 66533 2255 66591 2261
rect 66806 2252 66812 2304
rect 66864 2292 66870 2304
rect 67269 2295 67327 2301
rect 67269 2292 67281 2295
rect 66864 2264 67281 2292
rect 66864 2252 66870 2264
rect 67269 2261 67281 2264
rect 67315 2261 67327 2295
rect 67269 2255 67327 2261
rect 67542 2252 67548 2304
rect 67600 2292 67606 2304
rect 68373 2295 68431 2301
rect 68373 2292 68385 2295
rect 67600 2264 68385 2292
rect 67600 2252 67606 2264
rect 68373 2261 68385 2264
rect 68419 2261 68431 2295
rect 68373 2255 68431 2261
rect 68554 2252 68560 2304
rect 68612 2292 68618 2304
rect 69109 2295 69167 2301
rect 69109 2292 69121 2295
rect 68612 2264 69121 2292
rect 68612 2252 68618 2264
rect 69109 2261 69121 2264
rect 69155 2261 69167 2295
rect 69109 2255 69167 2261
rect 70486 2252 70492 2304
rect 70544 2292 70550 2304
rect 70949 2295 71007 2301
rect 70949 2292 70961 2295
rect 70544 2264 70961 2292
rect 70544 2252 70550 2264
rect 70949 2261 70961 2264
rect 70995 2261 71007 2295
rect 70949 2255 71007 2261
rect 71222 2252 71228 2304
rect 71280 2292 71286 2304
rect 71685 2295 71743 2301
rect 71685 2292 71697 2295
rect 71280 2264 71697 2292
rect 71280 2252 71286 2264
rect 71685 2261 71697 2264
rect 71731 2261 71743 2295
rect 71685 2255 71743 2261
rect 71958 2252 71964 2304
rect 72016 2292 72022 2304
rect 72421 2295 72479 2301
rect 72421 2292 72433 2295
rect 72016 2264 72433 2292
rect 72016 2252 72022 2264
rect 72421 2261 72433 2264
rect 72467 2261 72479 2295
rect 74506 2292 74534 2332
rect 76837 2295 76895 2301
rect 76837 2292 76849 2295
rect 74506 2264 76849 2292
rect 72421 2255 72479 2261
rect 76837 2261 76849 2264
rect 76883 2261 76895 2295
rect 76837 2255 76895 2261
rect 77110 2252 77116 2304
rect 77168 2292 77174 2304
rect 77573 2295 77631 2301
rect 77573 2292 77585 2295
rect 77168 2264 77585 2292
rect 77168 2252 77174 2264
rect 77573 2261 77585 2264
rect 77619 2261 77631 2295
rect 77573 2255 77631 2261
rect 1104 2202 78844 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 78844 2202
rect 1104 2128 78844 2150
<< via1 >>
rect 4214 77766 4266 77818
rect 4278 77766 4330 77818
rect 4342 77766 4394 77818
rect 4406 77766 4458 77818
rect 4470 77766 4522 77818
rect 34934 77766 34986 77818
rect 34998 77766 35050 77818
rect 35062 77766 35114 77818
rect 35126 77766 35178 77818
rect 35190 77766 35242 77818
rect 65654 77766 65706 77818
rect 65718 77766 65770 77818
rect 65782 77766 65834 77818
rect 65846 77766 65898 77818
rect 65910 77766 65962 77818
rect 19574 77222 19626 77274
rect 19638 77222 19690 77274
rect 19702 77222 19754 77274
rect 19766 77222 19818 77274
rect 19830 77222 19882 77274
rect 50294 77222 50346 77274
rect 50358 77222 50410 77274
rect 50422 77222 50474 77274
rect 50486 77222 50538 77274
rect 50550 77222 50602 77274
rect 4214 76678 4266 76730
rect 4278 76678 4330 76730
rect 4342 76678 4394 76730
rect 4406 76678 4458 76730
rect 4470 76678 4522 76730
rect 34934 76678 34986 76730
rect 34998 76678 35050 76730
rect 35062 76678 35114 76730
rect 35126 76678 35178 76730
rect 35190 76678 35242 76730
rect 65654 76678 65706 76730
rect 65718 76678 65770 76730
rect 65782 76678 65834 76730
rect 65846 76678 65898 76730
rect 65910 76678 65962 76730
rect 19574 76134 19626 76186
rect 19638 76134 19690 76186
rect 19702 76134 19754 76186
rect 19766 76134 19818 76186
rect 19830 76134 19882 76186
rect 50294 76134 50346 76186
rect 50358 76134 50410 76186
rect 50422 76134 50474 76186
rect 50486 76134 50538 76186
rect 50550 76134 50602 76186
rect 4214 75590 4266 75642
rect 4278 75590 4330 75642
rect 4342 75590 4394 75642
rect 4406 75590 4458 75642
rect 4470 75590 4522 75642
rect 34934 75590 34986 75642
rect 34998 75590 35050 75642
rect 35062 75590 35114 75642
rect 35126 75590 35178 75642
rect 35190 75590 35242 75642
rect 65654 75590 65706 75642
rect 65718 75590 65770 75642
rect 65782 75590 65834 75642
rect 65846 75590 65898 75642
rect 65910 75590 65962 75642
rect 1676 75327 1728 75336
rect 1676 75293 1685 75327
rect 1685 75293 1719 75327
rect 1719 75293 1728 75327
rect 1676 75284 1728 75293
rect 1492 75191 1544 75200
rect 1492 75157 1501 75191
rect 1501 75157 1535 75191
rect 1535 75157 1544 75191
rect 1492 75148 1544 75157
rect 76564 75148 76616 75200
rect 78036 75191 78088 75200
rect 78036 75157 78045 75191
rect 78045 75157 78079 75191
rect 78079 75157 78088 75191
rect 78036 75148 78088 75157
rect 19574 75046 19626 75098
rect 19638 75046 19690 75098
rect 19702 75046 19754 75098
rect 19766 75046 19818 75098
rect 19830 75046 19882 75098
rect 50294 75046 50346 75098
rect 50358 75046 50410 75098
rect 50422 75046 50474 75098
rect 50486 75046 50538 75098
rect 50550 75046 50602 75098
rect 1400 74851 1452 74860
rect 1400 74817 1409 74851
rect 1409 74817 1443 74851
rect 1443 74817 1452 74851
rect 1400 74808 1452 74817
rect 78128 74808 78180 74860
rect 77576 74672 77628 74724
rect 2412 74604 2464 74656
rect 4214 74502 4266 74554
rect 4278 74502 4330 74554
rect 4342 74502 4394 74554
rect 4406 74502 4458 74554
rect 4470 74502 4522 74554
rect 34934 74502 34986 74554
rect 34998 74502 35050 74554
rect 35062 74502 35114 74554
rect 35126 74502 35178 74554
rect 35190 74502 35242 74554
rect 65654 74502 65706 74554
rect 65718 74502 65770 74554
rect 65782 74502 65834 74554
rect 65846 74502 65898 74554
rect 65910 74502 65962 74554
rect 1400 74375 1452 74384
rect 1400 74341 1409 74375
rect 1409 74341 1443 74375
rect 1443 74341 1452 74375
rect 1400 74332 1452 74341
rect 78128 74375 78180 74384
rect 78128 74341 78137 74375
rect 78137 74341 78171 74375
rect 78171 74341 78180 74375
rect 78128 74332 78180 74341
rect 19574 73958 19626 74010
rect 19638 73958 19690 74010
rect 19702 73958 19754 74010
rect 19766 73958 19818 74010
rect 19830 73958 19882 74010
rect 50294 73958 50346 74010
rect 50358 73958 50410 74010
rect 50422 73958 50474 74010
rect 50486 73958 50538 74010
rect 50550 73958 50602 74010
rect 1492 73627 1544 73636
rect 1492 73593 1501 73627
rect 1501 73593 1535 73627
rect 1535 73593 1544 73627
rect 1492 73584 1544 73593
rect 2688 73516 2740 73568
rect 77024 73516 77076 73568
rect 77852 73627 77904 73636
rect 77852 73593 77861 73627
rect 77861 73593 77895 73627
rect 77895 73593 77904 73627
rect 77852 73584 77904 73593
rect 4214 73414 4266 73466
rect 4278 73414 4330 73466
rect 4342 73414 4394 73466
rect 4406 73414 4458 73466
rect 4470 73414 4522 73466
rect 34934 73414 34986 73466
rect 34998 73414 35050 73466
rect 35062 73414 35114 73466
rect 35126 73414 35178 73466
rect 35190 73414 35242 73466
rect 65654 73414 65706 73466
rect 65718 73414 65770 73466
rect 65782 73414 65834 73466
rect 65846 73414 65898 73466
rect 65910 73414 65962 73466
rect 1492 73015 1544 73024
rect 1492 72981 1501 73015
rect 1501 72981 1535 73015
rect 1535 72981 1544 73015
rect 1492 72972 1544 72981
rect 76196 73108 76248 73160
rect 2320 72972 2372 73024
rect 78036 73015 78088 73024
rect 78036 72981 78045 73015
rect 78045 72981 78079 73015
rect 78079 72981 78088 73015
rect 78036 72972 78088 72981
rect 19574 72870 19626 72922
rect 19638 72870 19690 72922
rect 19702 72870 19754 72922
rect 19766 72870 19818 72922
rect 19830 72870 19882 72922
rect 50294 72870 50346 72922
rect 50358 72870 50410 72922
rect 50422 72870 50474 72922
rect 50486 72870 50538 72922
rect 50550 72870 50602 72922
rect 1492 72471 1544 72480
rect 1492 72437 1501 72471
rect 1501 72437 1535 72471
rect 1535 72437 1544 72471
rect 1492 72428 1544 72437
rect 76104 72632 76156 72684
rect 2412 72428 2464 72480
rect 77852 72471 77904 72480
rect 77852 72437 77861 72471
rect 77861 72437 77895 72471
rect 77895 72437 77904 72471
rect 77852 72428 77904 72437
rect 4214 72326 4266 72378
rect 4278 72326 4330 72378
rect 4342 72326 4394 72378
rect 4406 72326 4458 72378
rect 4470 72326 4522 72378
rect 34934 72326 34986 72378
rect 34998 72326 35050 72378
rect 35062 72326 35114 72378
rect 35126 72326 35178 72378
rect 35190 72326 35242 72378
rect 65654 72326 65706 72378
rect 65718 72326 65770 72378
rect 65782 72326 65834 72378
rect 65846 72326 65898 72378
rect 65910 72326 65962 72378
rect 75920 72020 75972 72072
rect 1492 71927 1544 71936
rect 1492 71893 1501 71927
rect 1501 71893 1535 71927
rect 1535 71893 1544 71927
rect 1492 71884 1544 71893
rect 2228 71927 2280 71936
rect 2228 71893 2237 71927
rect 2237 71893 2271 71927
rect 2271 71893 2280 71927
rect 2228 71884 2280 71893
rect 78036 71927 78088 71936
rect 78036 71893 78045 71927
rect 78045 71893 78079 71927
rect 78079 71893 78088 71927
rect 78036 71884 78088 71893
rect 19574 71782 19626 71834
rect 19638 71782 19690 71834
rect 19702 71782 19754 71834
rect 19766 71782 19818 71834
rect 19830 71782 19882 71834
rect 50294 71782 50346 71834
rect 50358 71782 50410 71834
rect 50422 71782 50474 71834
rect 50486 71782 50538 71834
rect 50550 71782 50602 71834
rect 76196 71723 76248 71732
rect 76196 71689 76205 71723
rect 76205 71689 76239 71723
rect 76239 71689 76248 71723
rect 76196 71680 76248 71689
rect 76288 71544 76340 71596
rect 2320 71340 2372 71392
rect 76288 71340 76340 71392
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 34934 71238 34986 71290
rect 34998 71238 35050 71290
rect 35062 71238 35114 71290
rect 35126 71238 35178 71290
rect 35190 71238 35242 71290
rect 65654 71238 65706 71290
rect 65718 71238 65770 71290
rect 65782 71238 65834 71290
rect 65846 71238 65898 71290
rect 65910 71238 65962 71290
rect 76104 71179 76156 71188
rect 76104 71145 76113 71179
rect 76113 71145 76147 71179
rect 76147 71145 76156 71179
rect 76104 71136 76156 71145
rect 1492 70839 1544 70848
rect 1492 70805 1501 70839
rect 1501 70805 1535 70839
rect 1535 70805 1544 70839
rect 1492 70796 1544 70805
rect 76012 70932 76064 70984
rect 2412 70864 2464 70916
rect 2320 70796 2372 70848
rect 75828 70864 75880 70916
rect 78036 70839 78088 70848
rect 78036 70805 78045 70839
rect 78045 70805 78079 70839
rect 78079 70805 78088 70839
rect 78036 70796 78088 70805
rect 19574 70694 19626 70746
rect 19638 70694 19690 70746
rect 19702 70694 19754 70746
rect 19766 70694 19818 70746
rect 19830 70694 19882 70746
rect 50294 70694 50346 70746
rect 50358 70694 50410 70746
rect 50422 70694 50474 70746
rect 50486 70694 50538 70746
rect 50550 70694 50602 70746
rect 2228 70524 2280 70576
rect 75920 70592 75972 70644
rect 75000 70456 75052 70508
rect 2228 70431 2280 70440
rect 2228 70397 2237 70431
rect 2237 70397 2271 70431
rect 2271 70397 2280 70431
rect 2228 70388 2280 70397
rect 73344 70388 73396 70440
rect 1492 70295 1544 70304
rect 1492 70261 1501 70295
rect 1501 70261 1535 70295
rect 1535 70261 1544 70295
rect 1492 70252 1544 70261
rect 77852 70295 77904 70304
rect 77852 70261 77861 70295
rect 77861 70261 77895 70295
rect 77895 70261 77904 70295
rect 77852 70252 77904 70261
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 34934 70150 34986 70202
rect 34998 70150 35050 70202
rect 35062 70150 35114 70202
rect 35126 70150 35178 70202
rect 35190 70150 35242 70202
rect 65654 70150 65706 70202
rect 65718 70150 65770 70202
rect 65782 70150 65834 70202
rect 65846 70150 65898 70202
rect 65910 70150 65962 70202
rect 75828 70048 75880 70100
rect 1400 69887 1452 69896
rect 1400 69853 1409 69887
rect 1409 69853 1443 69887
rect 1443 69853 1452 69887
rect 1400 69844 1452 69853
rect 2320 69776 2372 69828
rect 1768 69708 1820 69760
rect 78128 69887 78180 69896
rect 78128 69853 78137 69887
rect 78137 69853 78171 69887
rect 78171 69853 78180 69887
rect 78128 69844 78180 69853
rect 74264 69708 74316 69760
rect 77944 69751 77996 69760
rect 77944 69717 77953 69751
rect 77953 69717 77987 69751
rect 77987 69717 77996 69751
rect 77944 69708 77996 69717
rect 19574 69606 19626 69658
rect 19638 69606 19690 69658
rect 19702 69606 19754 69658
rect 19766 69606 19818 69658
rect 19830 69606 19882 69658
rect 50294 69606 50346 69658
rect 50358 69606 50410 69658
rect 50422 69606 50474 69658
rect 50486 69606 50538 69658
rect 50550 69606 50602 69658
rect 65984 69504 66036 69556
rect 77944 69504 77996 69556
rect 1400 69411 1452 69420
rect 1400 69377 1409 69411
rect 1409 69377 1443 69411
rect 1443 69377 1452 69411
rect 1400 69368 1452 69377
rect 77944 69411 77996 69420
rect 77944 69377 77953 69411
rect 77953 69377 77987 69411
rect 77987 69377 77996 69411
rect 77944 69368 77996 69377
rect 1676 69164 1728 69216
rect 76656 69164 76708 69216
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 34934 69062 34986 69114
rect 34998 69062 35050 69114
rect 35062 69062 35114 69114
rect 35126 69062 35178 69114
rect 35190 69062 35242 69114
rect 65654 69062 65706 69114
rect 65718 69062 65770 69114
rect 65782 69062 65834 69114
rect 65846 69062 65898 69114
rect 65910 69062 65962 69114
rect 73344 69003 73396 69012
rect 73344 68969 73353 69003
rect 73353 68969 73387 69003
rect 73387 68969 73396 69003
rect 73344 68960 73396 68969
rect 1400 68663 1452 68672
rect 1400 68629 1409 68663
rect 1409 68629 1443 68663
rect 1443 68629 1452 68663
rect 1400 68620 1452 68629
rect 2228 68620 2280 68672
rect 73528 68620 73580 68672
rect 77944 68620 77996 68672
rect 19574 68518 19626 68570
rect 19638 68518 19690 68570
rect 19702 68518 19754 68570
rect 19766 68518 19818 68570
rect 19830 68518 19882 68570
rect 50294 68518 50346 68570
rect 50358 68518 50410 68570
rect 50422 68518 50474 68570
rect 50486 68518 50538 68570
rect 50550 68518 50602 68570
rect 1400 68323 1452 68332
rect 1400 68289 1409 68323
rect 1409 68289 1443 68323
rect 1443 68289 1452 68323
rect 1400 68280 1452 68289
rect 77944 68323 77996 68332
rect 77944 68289 77953 68323
rect 77953 68289 77987 68323
rect 77987 68289 77996 68323
rect 77944 68280 77996 68289
rect 66168 68076 66220 68128
rect 75184 68076 75236 68128
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 34934 67974 34986 68026
rect 34998 67974 35050 68026
rect 35062 67974 35114 68026
rect 35126 67974 35178 68026
rect 35190 67974 35242 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 1860 67804 1912 67856
rect 66996 67804 67048 67856
rect 1400 67711 1452 67720
rect 1400 67677 1409 67711
rect 1409 67677 1443 67711
rect 1443 67677 1452 67711
rect 1400 67668 1452 67677
rect 78128 67711 78180 67720
rect 78128 67677 78137 67711
rect 78137 67677 78171 67711
rect 78171 67677 78180 67711
rect 78128 67668 78180 67677
rect 19574 67430 19626 67482
rect 19638 67430 19690 67482
rect 19702 67430 19754 67482
rect 19766 67430 19818 67482
rect 19830 67430 19882 67482
rect 50294 67430 50346 67482
rect 50358 67430 50410 67482
rect 50422 67430 50474 67482
rect 50486 67430 50538 67482
rect 50550 67430 50602 67482
rect 1400 67235 1452 67244
rect 1400 67201 1409 67235
rect 1409 67201 1443 67235
rect 1443 67201 1452 67235
rect 1400 67192 1452 67201
rect 77944 67235 77996 67244
rect 77944 67201 77953 67235
rect 77953 67201 77987 67235
rect 77987 67201 77996 67235
rect 77944 67192 77996 67201
rect 72332 67056 72384 67108
rect 1584 67031 1636 67040
rect 1584 66997 1593 67031
rect 1593 66997 1627 67031
rect 1627 66997 1636 67031
rect 1584 66988 1636 66997
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 1584 66784 1636 66836
rect 63132 66784 63184 66836
rect 1400 66623 1452 66632
rect 1400 66589 1409 66623
rect 1409 66589 1443 66623
rect 1443 66589 1452 66623
rect 1400 66580 1452 66589
rect 78128 66623 78180 66632
rect 78128 66589 78137 66623
rect 78137 66589 78171 66623
rect 78171 66589 78180 66623
rect 78128 66580 78180 66589
rect 1584 66487 1636 66496
rect 1584 66453 1593 66487
rect 1593 66453 1627 66487
rect 1627 66453 1636 66487
rect 1584 66444 1636 66453
rect 77944 66487 77996 66496
rect 77944 66453 77953 66487
rect 77953 66453 77987 66487
rect 77987 66453 77996 66487
rect 77944 66444 77996 66453
rect 19574 66342 19626 66394
rect 19638 66342 19690 66394
rect 19702 66342 19754 66394
rect 19766 66342 19818 66394
rect 19830 66342 19882 66394
rect 50294 66342 50346 66394
rect 50358 66342 50410 66394
rect 50422 66342 50474 66394
rect 50486 66342 50538 66394
rect 50550 66342 50602 66394
rect 66076 66240 66128 66292
rect 77944 66240 77996 66292
rect 1400 65943 1452 65952
rect 1400 65909 1409 65943
rect 1409 65909 1443 65943
rect 1443 65909 1452 65943
rect 1400 65900 1452 65909
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 1400 65535 1452 65544
rect 1400 65501 1409 65535
rect 1409 65501 1443 65535
rect 1443 65501 1452 65535
rect 1400 65492 1452 65501
rect 78128 65535 78180 65544
rect 78128 65501 78137 65535
rect 78137 65501 78171 65535
rect 78171 65501 78180 65535
rect 78128 65492 78180 65501
rect 64512 65356 64564 65408
rect 76012 65356 76064 65408
rect 19574 65254 19626 65306
rect 19638 65254 19690 65306
rect 19702 65254 19754 65306
rect 19766 65254 19818 65306
rect 19830 65254 19882 65306
rect 50294 65254 50346 65306
rect 50358 65254 50410 65306
rect 50422 65254 50474 65306
rect 50486 65254 50538 65306
rect 50550 65254 50602 65306
rect 2320 65152 2372 65204
rect 1400 65059 1452 65068
rect 1400 65025 1409 65059
rect 1409 65025 1443 65059
rect 1443 65025 1452 65059
rect 1400 65016 1452 65025
rect 77944 65059 77996 65068
rect 77944 65025 77953 65059
rect 77953 65025 77987 65059
rect 77987 65025 77996 65059
rect 77944 65016 77996 65025
rect 72424 64948 72476 65000
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 34934 64710 34986 64762
rect 34998 64710 35050 64762
rect 35062 64710 35114 64762
rect 35126 64710 35178 64762
rect 35190 64710 35242 64762
rect 65654 64710 65706 64762
rect 65718 64710 65770 64762
rect 65782 64710 65834 64762
rect 65846 64710 65898 64762
rect 65910 64710 65962 64762
rect 1400 64447 1452 64456
rect 1400 64413 1409 64447
rect 1409 64413 1443 64447
rect 1443 64413 1452 64447
rect 1400 64404 1452 64413
rect 78128 64447 78180 64456
rect 78128 64413 78137 64447
rect 78137 64413 78171 64447
rect 78171 64413 78180 64447
rect 78128 64404 78180 64413
rect 1492 64268 1544 64320
rect 77484 64268 77536 64320
rect 19574 64166 19626 64218
rect 19638 64166 19690 64218
rect 19702 64166 19754 64218
rect 19766 64166 19818 64218
rect 19830 64166 19882 64218
rect 50294 64166 50346 64218
rect 50358 64166 50410 64218
rect 50422 64166 50474 64218
rect 50486 64166 50538 64218
rect 50550 64166 50602 64218
rect 1400 63971 1452 63980
rect 1400 63937 1409 63971
rect 1409 63937 1443 63971
rect 1443 63937 1452 63971
rect 1400 63928 1452 63937
rect 77944 63971 77996 63980
rect 77944 63937 77953 63971
rect 77953 63937 77987 63971
rect 77987 63937 77996 63971
rect 77944 63928 77996 63937
rect 2228 63724 2280 63776
rect 62672 63724 62724 63776
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 34934 63622 34986 63674
rect 34998 63622 35050 63674
rect 35062 63622 35114 63674
rect 35126 63622 35178 63674
rect 35190 63622 35242 63674
rect 65654 63622 65706 63674
rect 65718 63622 65770 63674
rect 65782 63622 65834 63674
rect 65846 63622 65898 63674
rect 65910 63622 65962 63674
rect 1400 63223 1452 63232
rect 1400 63189 1409 63223
rect 1409 63189 1443 63223
rect 1443 63189 1452 63223
rect 1400 63180 1452 63189
rect 77944 63180 77996 63232
rect 19574 63078 19626 63130
rect 19638 63078 19690 63130
rect 19702 63078 19754 63130
rect 19766 63078 19818 63130
rect 19830 63078 19882 63130
rect 50294 63078 50346 63130
rect 50358 63078 50410 63130
rect 50422 63078 50474 63130
rect 50486 63078 50538 63130
rect 50550 63078 50602 63130
rect 1400 62883 1452 62892
rect 1400 62849 1409 62883
rect 1409 62849 1443 62883
rect 1443 62849 1452 62883
rect 1400 62840 1452 62849
rect 77944 62883 77996 62892
rect 77944 62849 77953 62883
rect 77953 62849 77987 62883
rect 77987 62849 77996 62883
rect 77944 62840 77996 62849
rect 2136 62636 2188 62688
rect 77300 62636 77352 62688
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 34934 62534 34986 62586
rect 34998 62534 35050 62586
rect 35062 62534 35114 62586
rect 35126 62534 35178 62586
rect 35190 62534 35242 62586
rect 65654 62534 65706 62586
rect 65718 62534 65770 62586
rect 65782 62534 65834 62586
rect 65846 62534 65898 62586
rect 65910 62534 65962 62586
rect 65432 62432 65484 62484
rect 65984 62432 66036 62484
rect 1400 62271 1452 62280
rect 1400 62237 1409 62271
rect 1409 62237 1443 62271
rect 1443 62237 1452 62271
rect 1400 62228 1452 62237
rect 78128 62271 78180 62280
rect 78128 62237 78137 62271
rect 78137 62237 78171 62271
rect 78171 62237 78180 62271
rect 78128 62228 78180 62237
rect 1768 62160 1820 62212
rect 1952 62092 2004 62144
rect 64420 62092 64472 62144
rect 77392 62092 77444 62144
rect 19574 61990 19626 62042
rect 19638 61990 19690 62042
rect 19702 61990 19754 62042
rect 19766 61990 19818 62042
rect 19830 61990 19882 62042
rect 50294 61990 50346 62042
rect 50358 61990 50410 62042
rect 50422 61990 50474 62042
rect 50486 61990 50538 62042
rect 50550 61990 50602 62042
rect 64512 61931 64564 61940
rect 64512 61897 64521 61931
rect 64521 61897 64555 61931
rect 64555 61897 64564 61931
rect 64512 61888 64564 61897
rect 65524 61888 65576 61940
rect 66168 61931 66220 61940
rect 66168 61897 66177 61931
rect 66177 61897 66211 61931
rect 66211 61897 66220 61931
rect 66168 61888 66220 61897
rect 65340 61820 65392 61872
rect 66076 61820 66128 61872
rect 1400 61795 1452 61804
rect 1400 61761 1409 61795
rect 1409 61761 1443 61795
rect 1443 61761 1452 61795
rect 1400 61752 1452 61761
rect 64052 61795 64104 61804
rect 64052 61761 64061 61795
rect 64061 61761 64095 61795
rect 64095 61761 64104 61795
rect 64052 61752 64104 61761
rect 77944 61795 77996 61804
rect 77944 61761 77953 61795
rect 77953 61761 77987 61795
rect 77987 61761 77996 61795
rect 77944 61752 77996 61761
rect 61660 61616 61712 61668
rect 64328 61616 64380 61668
rect 2412 61548 2464 61600
rect 2688 61548 2740 61600
rect 66076 61548 66128 61600
rect 77760 61591 77812 61600
rect 77760 61557 77769 61591
rect 77769 61557 77803 61591
rect 77803 61557 77812 61591
rect 77760 61548 77812 61557
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 65654 61446 65706 61498
rect 65718 61446 65770 61498
rect 65782 61446 65834 61498
rect 65846 61446 65898 61498
rect 65910 61446 65962 61498
rect 1584 61344 1636 61396
rect 61660 61344 61712 61396
rect 63132 61387 63184 61396
rect 63132 61353 63141 61387
rect 63141 61353 63175 61387
rect 63175 61353 63184 61387
rect 63132 61344 63184 61353
rect 63224 61344 63276 61396
rect 64972 61319 65024 61328
rect 64972 61285 64981 61319
rect 64981 61285 65015 61319
rect 65015 61285 65024 61319
rect 64972 61276 65024 61285
rect 66168 61319 66220 61328
rect 66168 61285 66177 61319
rect 66177 61285 66211 61319
rect 66211 61285 66220 61319
rect 66168 61276 66220 61285
rect 77760 61208 77812 61260
rect 1400 61183 1452 61192
rect 1400 61149 1409 61183
rect 1409 61149 1443 61183
rect 1443 61149 1452 61183
rect 1400 61140 1452 61149
rect 63960 61183 64012 61192
rect 63960 61149 63969 61183
rect 63969 61149 64003 61183
rect 64003 61149 64012 61183
rect 63960 61140 64012 61149
rect 64420 61183 64472 61192
rect 64420 61149 64429 61183
rect 64429 61149 64463 61183
rect 64463 61149 64472 61183
rect 64420 61140 64472 61149
rect 65248 61140 65300 61192
rect 65524 61140 65576 61192
rect 65984 61183 66036 61192
rect 65984 61149 65998 61183
rect 65998 61149 66032 61183
rect 66032 61149 66036 61183
rect 66720 61183 66772 61192
rect 65984 61140 66036 61149
rect 66720 61149 66729 61183
rect 66729 61149 66763 61183
rect 66763 61149 66772 61183
rect 66720 61140 66772 61149
rect 63684 61072 63736 61124
rect 2044 61004 2096 61056
rect 63776 61047 63828 61056
rect 63776 61013 63785 61047
rect 63785 61013 63819 61047
rect 63819 61013 63828 61047
rect 63776 61004 63828 61013
rect 65432 61072 65484 61124
rect 75184 61140 75236 61192
rect 78128 61183 78180 61192
rect 78128 61149 78137 61183
rect 78137 61149 78171 61183
rect 78171 61149 78180 61183
rect 78128 61140 78180 61149
rect 77024 61072 77076 61124
rect 77944 61047 77996 61056
rect 77944 61013 77953 61047
rect 77953 61013 77987 61047
rect 77987 61013 77996 61047
rect 77944 61004 77996 61013
rect 19574 60902 19626 60954
rect 19638 60902 19690 60954
rect 19702 60902 19754 60954
rect 19766 60902 19818 60954
rect 19830 60902 19882 60954
rect 50294 60902 50346 60954
rect 50358 60902 50410 60954
rect 50422 60902 50474 60954
rect 50486 60902 50538 60954
rect 50550 60902 50602 60954
rect 64052 60800 64104 60852
rect 60004 60732 60056 60784
rect 77944 60732 77996 60784
rect 63684 60664 63736 60716
rect 64328 60664 64380 60716
rect 64604 60707 64656 60716
rect 64604 60673 64613 60707
rect 64613 60673 64647 60707
rect 64647 60673 64656 60707
rect 64604 60664 64656 60673
rect 64788 60707 64840 60716
rect 64788 60673 64802 60707
rect 64802 60673 64836 60707
rect 64836 60673 64840 60707
rect 64788 60664 64840 60673
rect 65248 60664 65300 60716
rect 65432 60664 65484 60716
rect 65984 60664 66036 60716
rect 65340 60596 65392 60648
rect 65524 60639 65576 60648
rect 65524 60605 65533 60639
rect 65533 60605 65567 60639
rect 65567 60605 65576 60639
rect 65524 60596 65576 60605
rect 76564 60596 76616 60648
rect 67364 60528 67416 60580
rect 1400 60503 1452 60512
rect 1400 60469 1409 60503
rect 1409 60469 1443 60503
rect 1443 60469 1452 60503
rect 1400 60460 1452 60469
rect 63040 60503 63092 60512
rect 63040 60469 63049 60503
rect 63049 60469 63083 60503
rect 63083 60469 63092 60503
rect 63040 60460 63092 60469
rect 65156 60460 65208 60512
rect 65524 60460 65576 60512
rect 66076 60460 66128 60512
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 65654 60358 65706 60410
rect 65718 60358 65770 60410
rect 65782 60358 65834 60410
rect 65846 60358 65898 60410
rect 65910 60358 65962 60410
rect 62672 60299 62724 60308
rect 62672 60265 62681 60299
rect 62681 60265 62715 60299
rect 62715 60265 62724 60299
rect 62672 60256 62724 60265
rect 63960 60299 64012 60308
rect 63960 60265 63969 60299
rect 63969 60265 64003 60299
rect 64003 60265 64012 60299
rect 63960 60256 64012 60265
rect 59544 60188 59596 60240
rect 65248 60256 65300 60308
rect 66720 60299 66772 60308
rect 66720 60265 66729 60299
rect 66729 60265 66763 60299
rect 66763 60265 66772 60299
rect 66720 60256 66772 60265
rect 65064 60188 65116 60240
rect 1400 60095 1452 60104
rect 1400 60061 1409 60095
rect 1409 60061 1443 60095
rect 1443 60061 1452 60095
rect 1400 60052 1452 60061
rect 63592 60095 63644 60104
rect 63592 60061 63601 60095
rect 63601 60061 63635 60095
rect 63635 60061 63644 60095
rect 63592 60052 63644 60061
rect 63684 60052 63736 60104
rect 64512 60052 64564 60104
rect 64788 60095 64840 60104
rect 64788 60061 64802 60095
rect 64802 60061 64836 60095
rect 64836 60061 64840 60095
rect 65616 60095 65668 60104
rect 64788 60052 64840 60061
rect 65616 60061 65625 60095
rect 65625 60061 65659 60095
rect 65659 60061 65668 60095
rect 65616 60052 65668 60061
rect 66076 60188 66128 60240
rect 68100 60231 68152 60240
rect 68100 60197 68109 60231
rect 68109 60197 68143 60231
rect 68143 60197 68152 60231
rect 68100 60188 68152 60197
rect 76656 60256 76708 60308
rect 65984 60095 66036 60104
rect 65984 60061 65998 60095
rect 65998 60061 66032 60095
rect 66032 60061 66036 60095
rect 65984 60052 66036 60061
rect 67364 60052 67416 60104
rect 78128 60095 78180 60104
rect 78128 60061 78137 60095
rect 78137 60061 78171 60095
rect 78171 60061 78180 60095
rect 78128 60052 78180 60061
rect 64604 60027 64656 60036
rect 64604 59993 64613 60027
rect 64613 59993 64647 60027
rect 64647 59993 64656 60027
rect 64604 59984 64656 59993
rect 2596 59916 2648 59968
rect 65708 59984 65760 60036
rect 66996 59984 67048 60036
rect 76012 59984 76064 60036
rect 77944 59959 77996 59968
rect 77944 59925 77953 59959
rect 77953 59925 77987 59959
rect 77987 59925 77996 59959
rect 77944 59916 77996 59925
rect 19574 59814 19626 59866
rect 19638 59814 19690 59866
rect 19702 59814 19754 59866
rect 19766 59814 19818 59866
rect 19830 59814 19882 59866
rect 50294 59814 50346 59866
rect 50358 59814 50410 59866
rect 50422 59814 50474 59866
rect 50486 59814 50538 59866
rect 50550 59814 50602 59866
rect 62120 59712 62172 59764
rect 63224 59712 63276 59764
rect 64880 59712 64932 59764
rect 64696 59687 64748 59696
rect 1400 59619 1452 59628
rect 1400 59585 1409 59619
rect 1409 59585 1443 59619
rect 1443 59585 1452 59619
rect 1400 59576 1452 59585
rect 63132 59576 63184 59628
rect 63776 59619 63828 59628
rect 63776 59585 63779 59619
rect 63779 59585 63828 59619
rect 2320 59508 2372 59560
rect 63776 59576 63828 59585
rect 64420 59619 64472 59628
rect 64420 59585 64429 59619
rect 64429 59585 64463 59619
rect 64463 59585 64472 59619
rect 64420 59576 64472 59585
rect 64696 59653 64705 59687
rect 64705 59653 64739 59687
rect 64739 59653 64748 59687
rect 64696 59644 64748 59653
rect 65248 59712 65300 59764
rect 77944 59712 77996 59764
rect 64604 59619 64656 59628
rect 64604 59585 64613 59619
rect 64613 59585 64647 59619
rect 64647 59585 64656 59619
rect 64604 59576 64656 59585
rect 2228 59440 2280 59492
rect 2688 59372 2740 59424
rect 64420 59440 64472 59492
rect 61844 59372 61896 59424
rect 63868 59415 63920 59424
rect 63868 59381 63877 59415
rect 63877 59381 63911 59415
rect 63911 59381 63920 59415
rect 63868 59372 63920 59381
rect 65248 59508 65300 59560
rect 65340 59440 65392 59492
rect 65800 59619 65852 59628
rect 65800 59585 65809 59619
rect 65809 59585 65843 59619
rect 65843 59585 65852 59619
rect 67180 59644 67232 59696
rect 72424 59644 72476 59696
rect 65800 59576 65852 59585
rect 77944 59619 77996 59628
rect 77944 59585 77953 59619
rect 77953 59585 77987 59619
rect 77987 59585 77996 59619
rect 77944 59576 77996 59585
rect 65708 59440 65760 59492
rect 72332 59508 72384 59560
rect 65984 59372 66036 59424
rect 67180 59415 67232 59424
rect 67180 59381 67189 59415
rect 67189 59381 67223 59415
rect 67223 59381 67232 59415
rect 67180 59372 67232 59381
rect 77760 59415 77812 59424
rect 77760 59381 77769 59415
rect 77769 59381 77803 59415
rect 77803 59381 77812 59415
rect 77760 59372 77812 59381
rect 4214 59270 4266 59322
rect 4278 59270 4330 59322
rect 4342 59270 4394 59322
rect 4406 59270 4458 59322
rect 4470 59270 4522 59322
rect 34934 59270 34986 59322
rect 34998 59270 35050 59322
rect 35062 59270 35114 59322
rect 35126 59270 35178 59322
rect 35190 59270 35242 59322
rect 65654 59270 65706 59322
rect 65718 59270 65770 59322
rect 65782 59270 65834 59322
rect 65846 59270 65898 59322
rect 65910 59270 65962 59322
rect 63684 59168 63736 59220
rect 64604 59168 64656 59220
rect 65432 59168 65484 59220
rect 62488 59100 62540 59152
rect 64696 59100 64748 59152
rect 67180 59100 67232 59152
rect 60280 59032 60332 59084
rect 1400 59007 1452 59016
rect 1400 58973 1409 59007
rect 1409 58973 1443 59007
rect 1443 58973 1452 59007
rect 1400 58964 1452 58973
rect 2412 58964 2464 59016
rect 61660 58964 61712 59016
rect 61844 59007 61896 59016
rect 61844 58973 61853 59007
rect 61853 58973 61887 59007
rect 61887 58973 61896 59007
rect 61844 58964 61896 58973
rect 62212 59007 62264 59016
rect 62212 58973 62226 59007
rect 62226 58973 62260 59007
rect 62260 58973 62264 59007
rect 63132 59007 63184 59016
rect 62212 58964 62264 58973
rect 63132 58973 63141 59007
rect 63141 58973 63175 59007
rect 63175 58973 63184 59007
rect 63132 58964 63184 58973
rect 65616 59007 65668 59016
rect 61936 58896 61988 58948
rect 62672 58896 62724 58948
rect 65616 58973 65625 59007
rect 65625 58973 65659 59007
rect 65659 58973 65668 59007
rect 65616 58964 65668 58973
rect 78128 59007 78180 59016
rect 78128 58973 78137 59007
rect 78137 58973 78171 59007
rect 78171 58973 78180 59007
rect 78128 58964 78180 58973
rect 77760 58896 77812 58948
rect 1584 58871 1636 58880
rect 1584 58837 1593 58871
rect 1593 58837 1627 58871
rect 1627 58837 1636 58871
rect 1584 58828 1636 58837
rect 59820 58871 59872 58880
rect 59820 58837 59829 58871
rect 59829 58837 59863 58871
rect 59863 58837 59872 58871
rect 59820 58828 59872 58837
rect 61292 58871 61344 58880
rect 61292 58837 61301 58871
rect 61301 58837 61335 58871
rect 61335 58837 61344 58871
rect 61292 58828 61344 58837
rect 67364 58871 67416 58880
rect 67364 58837 67373 58871
rect 67373 58837 67407 58871
rect 67407 58837 67416 58871
rect 67364 58828 67416 58837
rect 77944 58871 77996 58880
rect 77944 58837 77953 58871
rect 77953 58837 77987 58871
rect 77987 58837 77996 58871
rect 77944 58828 77996 58837
rect 19574 58726 19626 58778
rect 19638 58726 19690 58778
rect 19702 58726 19754 58778
rect 19766 58726 19818 58778
rect 19830 58726 19882 58778
rect 50294 58726 50346 58778
rect 50358 58726 50410 58778
rect 50422 58726 50474 58778
rect 50486 58726 50538 58778
rect 50550 58726 50602 58778
rect 2688 58624 2740 58676
rect 59544 58667 59596 58676
rect 1584 58556 1636 58608
rect 1400 58531 1452 58540
rect 1400 58497 1409 58531
rect 1409 58497 1443 58531
rect 1443 58497 1452 58531
rect 1400 58488 1452 58497
rect 59544 58633 59553 58667
rect 59553 58633 59587 58667
rect 59587 58633 59596 58667
rect 59544 58624 59596 58633
rect 61292 58624 61344 58676
rect 60280 58599 60332 58608
rect 60280 58565 60289 58599
rect 60289 58565 60323 58599
rect 60323 58565 60332 58599
rect 60280 58556 60332 58565
rect 62120 58599 62172 58608
rect 62120 58565 62129 58599
rect 62129 58565 62163 58599
rect 62163 58565 62172 58599
rect 62120 58556 62172 58565
rect 64420 58624 64472 58676
rect 66996 58624 67048 58676
rect 77944 58624 77996 58676
rect 59820 58488 59872 58540
rect 60188 58531 60240 58540
rect 60188 58497 60197 58531
rect 60197 58497 60231 58531
rect 60231 58497 60240 58531
rect 60188 58488 60240 58497
rect 60372 58531 60424 58540
rect 60372 58497 60386 58531
rect 60386 58497 60420 58531
rect 60420 58497 60424 58531
rect 60372 58488 60424 58497
rect 61660 58488 61712 58540
rect 61936 58488 61988 58540
rect 62212 58531 62264 58540
rect 62212 58497 62226 58531
rect 62226 58497 62260 58531
rect 62260 58497 62264 58531
rect 62212 58488 62264 58497
rect 63776 58488 63828 58540
rect 77944 58531 77996 58540
rect 77944 58497 77953 58531
rect 77953 58497 77987 58531
rect 77987 58497 77996 58531
rect 77944 58488 77996 58497
rect 2136 58352 2188 58404
rect 61016 58352 61068 58404
rect 64880 58420 64932 58472
rect 65616 58420 65668 58472
rect 2688 58284 2740 58336
rect 60556 58327 60608 58336
rect 60556 58293 60565 58327
rect 60565 58293 60599 58327
rect 60599 58293 60608 58327
rect 60556 58284 60608 58293
rect 61108 58327 61160 58336
rect 61108 58293 61117 58327
rect 61117 58293 61151 58327
rect 61151 58293 61160 58327
rect 61108 58284 61160 58293
rect 62396 58327 62448 58336
rect 62396 58293 62405 58327
rect 62405 58293 62439 58327
rect 62439 58293 62448 58327
rect 62396 58284 62448 58293
rect 63592 58327 63644 58336
rect 63592 58293 63601 58327
rect 63601 58293 63635 58327
rect 63635 58293 63644 58327
rect 63592 58284 63644 58293
rect 77760 58327 77812 58336
rect 77760 58293 77769 58327
rect 77769 58293 77803 58327
rect 77803 58293 77812 58327
rect 77760 58284 77812 58293
rect 4214 58182 4266 58234
rect 4278 58182 4330 58234
rect 4342 58182 4394 58234
rect 4406 58182 4458 58234
rect 4470 58182 4522 58234
rect 34934 58182 34986 58234
rect 34998 58182 35050 58234
rect 35062 58182 35114 58234
rect 35126 58182 35178 58234
rect 35190 58182 35242 58234
rect 65654 58182 65706 58234
rect 65718 58182 65770 58234
rect 65782 58182 65834 58234
rect 65846 58182 65898 58234
rect 65910 58182 65962 58234
rect 62212 58080 62264 58132
rect 63224 58080 63276 58132
rect 59544 57919 59596 57928
rect 2596 57808 2648 57860
rect 59544 57885 59553 57919
rect 59553 57885 59587 57919
rect 59587 57885 59596 57919
rect 59544 57876 59596 57885
rect 59728 57919 59780 57928
rect 59728 57885 59731 57919
rect 59731 57885 59780 57919
rect 59728 57876 59780 57885
rect 60372 57876 60424 57928
rect 61292 58012 61344 58064
rect 61016 57944 61068 57996
rect 63592 58012 63644 58064
rect 61108 57919 61160 57928
rect 61108 57885 61117 57919
rect 61117 57885 61151 57919
rect 61151 57885 61160 57919
rect 61108 57876 61160 57885
rect 61752 57919 61804 57928
rect 61752 57885 61761 57919
rect 61761 57885 61795 57919
rect 61795 57885 61804 57919
rect 61752 57876 61804 57885
rect 62120 57919 62172 57928
rect 62120 57885 62134 57919
rect 62134 57885 62168 57919
rect 62168 57885 62172 57919
rect 62120 57876 62172 57885
rect 62304 57919 62356 57928
rect 62304 57885 62330 57919
rect 62330 57885 62356 57919
rect 62304 57876 62356 57885
rect 60188 57808 60240 57860
rect 60464 57808 60516 57860
rect 1400 57783 1452 57792
rect 1400 57749 1409 57783
rect 1409 57749 1443 57783
rect 1443 57749 1452 57783
rect 1400 57740 1452 57749
rect 59544 57740 59596 57792
rect 59820 57783 59872 57792
rect 59820 57749 59837 57783
rect 59837 57749 59871 57783
rect 59871 57749 59872 57783
rect 59820 57740 59872 57749
rect 60648 57740 60700 57792
rect 61384 57808 61436 57860
rect 61936 57851 61988 57860
rect 61936 57817 61945 57851
rect 61945 57817 61979 57851
rect 61979 57817 61988 57851
rect 61936 57808 61988 57817
rect 63224 57919 63276 57928
rect 63224 57885 63238 57919
rect 63238 57885 63272 57919
rect 63272 57885 63276 57919
rect 63224 57876 63276 57885
rect 63592 57876 63644 57928
rect 65340 57876 65392 57928
rect 77300 57808 77352 57860
rect 63224 57740 63276 57792
rect 63316 57740 63368 57792
rect 63592 57740 63644 57792
rect 77484 57740 77536 57792
rect 77944 57740 77996 57792
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 1492 57536 1544 57588
rect 1400 57443 1452 57452
rect 1400 57409 1409 57443
rect 1409 57409 1443 57443
rect 1443 57409 1452 57443
rect 1400 57400 1452 57409
rect 59636 57511 59688 57520
rect 59636 57477 59645 57511
rect 59645 57477 59679 57511
rect 59679 57477 59688 57511
rect 59636 57468 59688 57477
rect 77760 57468 77812 57520
rect 59544 57443 59596 57452
rect 59544 57409 59553 57443
rect 59553 57409 59587 57443
rect 59587 57409 59596 57443
rect 59544 57400 59596 57409
rect 59728 57443 59780 57452
rect 59728 57409 59742 57443
rect 59742 57409 59776 57443
rect 59776 57409 59780 57443
rect 59728 57400 59780 57409
rect 61752 57400 61804 57452
rect 63040 57443 63092 57452
rect 63040 57409 63049 57443
rect 63049 57409 63083 57443
rect 63083 57409 63092 57443
rect 63040 57400 63092 57409
rect 63224 57443 63276 57452
rect 63224 57409 63233 57443
rect 63233 57409 63267 57443
rect 63267 57409 63276 57443
rect 63224 57400 63276 57409
rect 61384 57375 61436 57384
rect 61384 57341 61393 57375
rect 61393 57341 61427 57375
rect 61427 57341 61436 57375
rect 61384 57332 61436 57341
rect 63408 57443 63460 57452
rect 63408 57409 63422 57443
rect 63422 57409 63456 57443
rect 63456 57409 63460 57443
rect 77944 57443 77996 57452
rect 63408 57400 63460 57409
rect 77944 57409 77953 57443
rect 77953 57409 77987 57443
rect 77987 57409 77996 57443
rect 77944 57400 77996 57409
rect 1584 57239 1636 57248
rect 1584 57205 1593 57239
rect 1593 57205 1627 57239
rect 1627 57205 1636 57239
rect 1584 57196 1636 57205
rect 2688 57196 2740 57248
rect 60832 57264 60884 57316
rect 64328 57264 64380 57316
rect 77392 57264 77444 57316
rect 59636 57196 59688 57248
rect 60280 57196 60332 57248
rect 77760 57239 77812 57248
rect 77760 57205 77769 57239
rect 77769 57205 77803 57239
rect 77803 57205 77812 57239
rect 77760 57196 77812 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 63040 57035 63092 57044
rect 1952 56856 2004 56908
rect 63040 57001 63049 57035
rect 63049 57001 63083 57035
rect 63083 57001 63092 57035
rect 63040 56992 63092 57001
rect 59820 56967 59872 56976
rect 59820 56933 59829 56967
rect 59829 56933 59863 56967
rect 59863 56933 59872 56967
rect 59820 56924 59872 56933
rect 60464 56924 60516 56976
rect 59084 56856 59136 56908
rect 1400 56831 1452 56840
rect 1400 56797 1409 56831
rect 1409 56797 1443 56831
rect 1443 56797 1452 56831
rect 1400 56788 1452 56797
rect 59452 56831 59504 56840
rect 2044 56720 2096 56772
rect 59452 56797 59461 56831
rect 59461 56797 59495 56831
rect 59495 56797 59504 56831
rect 59452 56788 59504 56797
rect 59728 56831 59780 56840
rect 59728 56797 59731 56831
rect 59731 56797 59780 56831
rect 59728 56788 59780 56797
rect 77760 56992 77812 57044
rect 59544 56763 59596 56772
rect 59544 56729 59553 56763
rect 59553 56729 59587 56763
rect 59587 56729 59596 56763
rect 59544 56720 59596 56729
rect 60004 56720 60056 56772
rect 2688 56652 2740 56704
rect 60740 56720 60792 56772
rect 62120 56788 62172 56840
rect 78128 56831 78180 56840
rect 78128 56797 78137 56831
rect 78137 56797 78171 56831
rect 78171 56797 78180 56831
rect 78128 56788 78180 56797
rect 60832 56652 60884 56704
rect 76196 56652 76248 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 1584 56448 1636 56500
rect 57704 56448 57756 56500
rect 59544 56448 59596 56500
rect 57888 56380 57940 56432
rect 1400 56355 1452 56364
rect 1400 56321 1409 56355
rect 1409 56321 1443 56355
rect 1443 56321 1452 56355
rect 1400 56312 1452 56321
rect 59728 56312 59780 56364
rect 76196 56312 76248 56364
rect 77944 56355 77996 56364
rect 77944 56321 77953 56355
rect 77953 56321 77987 56355
rect 77987 56321 77996 56355
rect 77944 56312 77996 56321
rect 60740 56287 60792 56296
rect 60740 56253 60749 56287
rect 60749 56253 60783 56287
rect 60783 56253 60792 56287
rect 61200 56287 61252 56296
rect 60740 56244 60792 56253
rect 61200 56253 61209 56287
rect 61209 56253 61243 56287
rect 61243 56253 61252 56287
rect 61200 56244 61252 56253
rect 63132 56244 63184 56296
rect 55956 56176 56008 56228
rect 56784 56176 56836 56228
rect 57152 56108 57204 56160
rect 60832 56108 60884 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 55956 55947 56008 55956
rect 55956 55913 55965 55947
rect 55965 55913 55999 55947
rect 55999 55913 56008 55947
rect 55956 55904 56008 55913
rect 57152 55904 57204 55956
rect 2688 55700 2740 55752
rect 1492 55675 1544 55684
rect 1492 55641 1501 55675
rect 1501 55641 1535 55675
rect 1535 55641 1544 55675
rect 1492 55632 1544 55641
rect 57060 55879 57112 55888
rect 57060 55845 57069 55879
rect 57069 55845 57103 55879
rect 57103 55845 57112 55879
rect 57060 55836 57112 55845
rect 58440 55836 58492 55888
rect 60740 55836 60792 55888
rect 56784 55743 56836 55752
rect 56784 55709 56793 55743
rect 56793 55709 56827 55743
rect 56827 55709 56836 55743
rect 56784 55700 56836 55709
rect 56876 55743 56928 55752
rect 56876 55709 56890 55743
rect 56890 55709 56924 55743
rect 56924 55709 56928 55743
rect 56876 55700 56928 55709
rect 57888 55743 57940 55752
rect 57888 55709 57897 55743
rect 57897 55709 57931 55743
rect 57931 55709 57940 55743
rect 57888 55700 57940 55709
rect 57796 55675 57848 55684
rect 55680 55564 55732 55616
rect 56600 55564 56652 55616
rect 57796 55641 57805 55675
rect 57805 55641 57839 55675
rect 57839 55641 57848 55675
rect 57796 55632 57848 55641
rect 56876 55564 56928 55616
rect 57888 55564 57940 55616
rect 60464 55700 60516 55752
rect 64880 55700 64932 55752
rect 78128 55743 78180 55752
rect 78128 55709 78137 55743
rect 78137 55709 78171 55743
rect 78171 55709 78180 55743
rect 78128 55700 78180 55709
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 55680 55403 55732 55412
rect 55680 55369 55689 55403
rect 55689 55369 55723 55403
rect 55723 55369 55732 55403
rect 55680 55360 55732 55369
rect 57888 55360 57940 55412
rect 57152 55292 57204 55344
rect 57796 55292 57848 55344
rect 56692 55267 56744 55276
rect 56692 55233 56695 55267
rect 56695 55233 56744 55267
rect 56692 55224 56744 55233
rect 57704 55224 57756 55276
rect 56600 55088 56652 55140
rect 58992 55224 59044 55276
rect 60464 55224 60516 55276
rect 61200 55267 61252 55276
rect 61200 55233 61209 55267
rect 61209 55233 61243 55267
rect 61243 55233 61252 55267
rect 61200 55224 61252 55233
rect 59084 55156 59136 55208
rect 1492 55063 1544 55072
rect 1492 55029 1501 55063
rect 1501 55029 1535 55063
rect 1535 55029 1544 55063
rect 1492 55020 1544 55029
rect 57152 55020 57204 55072
rect 78128 55020 78180 55072
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 59084 54816 59136 54868
rect 53104 54680 53156 54732
rect 60832 54748 60884 54800
rect 56692 54680 56744 54732
rect 1492 54655 1544 54664
rect 1492 54621 1501 54655
rect 1501 54621 1535 54655
rect 1535 54621 1544 54655
rect 1492 54612 1544 54621
rect 56600 54655 56652 54664
rect 56600 54621 56609 54655
rect 56609 54621 56643 54655
rect 56643 54621 56652 54655
rect 56600 54612 56652 54621
rect 53380 54544 53432 54596
rect 60740 54612 60792 54664
rect 77944 54612 77996 54664
rect 78128 54655 78180 54664
rect 78128 54621 78137 54655
rect 78137 54621 78171 54655
rect 78171 54621 78180 54655
rect 78128 54612 78180 54621
rect 55496 54476 55548 54528
rect 76196 54476 76248 54528
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 55496 54315 55548 54324
rect 55496 54281 55505 54315
rect 55505 54281 55539 54315
rect 55539 54281 55548 54315
rect 55496 54272 55548 54281
rect 1492 54179 1544 54188
rect 1492 54145 1501 54179
rect 1501 54145 1535 54179
rect 1535 54145 1544 54179
rect 1492 54136 1544 54145
rect 56600 54204 56652 54256
rect 56692 54136 56744 54188
rect 1676 54043 1728 54052
rect 1676 54009 1685 54043
rect 1685 54009 1719 54043
rect 1719 54009 1728 54043
rect 1676 54000 1728 54009
rect 56600 53975 56652 53984
rect 56600 53941 56609 53975
rect 56609 53941 56643 53975
rect 56643 53941 56652 53975
rect 56600 53932 56652 53941
rect 77484 54068 77536 54120
rect 77944 54111 77996 54120
rect 77944 54077 77953 54111
rect 77953 54077 77987 54111
rect 77987 54077 77996 54111
rect 77944 54068 77996 54077
rect 76196 53932 76248 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 77300 53567 77352 53576
rect 77300 53533 77309 53567
rect 77309 53533 77343 53567
rect 77343 53533 77352 53567
rect 77300 53524 77352 53533
rect 77392 53524 77444 53576
rect 1492 53499 1544 53508
rect 1492 53465 1501 53499
rect 1501 53465 1535 53499
rect 1535 53465 1544 53499
rect 1492 53456 1544 53465
rect 53288 53456 53340 53508
rect 77668 53456 77720 53508
rect 2688 53388 2740 53440
rect 54116 53388 54168 53440
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 1676 53116 1728 53168
rect 53288 53159 53340 53168
rect 1492 53091 1544 53100
rect 1492 53057 1501 53091
rect 1501 53057 1535 53091
rect 1535 53057 1544 53091
rect 1492 53048 1544 53057
rect 52828 53048 52880 53100
rect 53288 53125 53297 53159
rect 53297 53125 53331 53159
rect 53331 53125 53340 53159
rect 53288 53116 53340 53125
rect 53196 53091 53248 53100
rect 53196 53057 53205 53091
rect 53205 53057 53239 53091
rect 53239 53057 53248 53091
rect 53196 53048 53248 53057
rect 53840 53048 53892 53100
rect 54116 53091 54168 53100
rect 54116 53057 54125 53091
rect 54125 53057 54159 53091
rect 54159 53057 54168 53091
rect 54116 53048 54168 53057
rect 77668 53091 77720 53100
rect 53196 52912 53248 52964
rect 77668 53057 77677 53091
rect 77677 53057 77711 53091
rect 77711 53057 77720 53091
rect 77668 53048 77720 53057
rect 53288 52844 53340 52896
rect 55220 52844 55272 52896
rect 77576 52980 77628 53032
rect 77484 52844 77536 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 52828 52683 52880 52692
rect 52828 52649 52837 52683
rect 52837 52649 52871 52683
rect 52871 52649 52880 52683
rect 52828 52640 52880 52649
rect 77576 52615 77628 52624
rect 77576 52581 77585 52615
rect 77585 52581 77619 52615
rect 77619 52581 77628 52615
rect 77576 52572 77628 52581
rect 51816 52504 51868 52556
rect 77392 52504 77444 52556
rect 53380 52479 53432 52488
rect 53380 52445 53389 52479
rect 53389 52445 53423 52479
rect 53423 52445 53432 52479
rect 53380 52436 53432 52445
rect 52184 52368 52236 52420
rect 53840 52436 53892 52488
rect 1492 52343 1544 52352
rect 1492 52309 1501 52343
rect 1501 52309 1535 52343
rect 1535 52309 1544 52343
rect 1492 52300 1544 52309
rect 55036 52300 55088 52352
rect 77944 52300 77996 52352
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 51816 52071 51868 52080
rect 51816 52037 51825 52071
rect 51825 52037 51859 52071
rect 51859 52037 51868 52071
rect 51816 52028 51868 52037
rect 1492 52003 1544 52012
rect 1492 51969 1501 52003
rect 1501 51969 1535 52003
rect 1535 51969 1544 52003
rect 1492 51960 1544 51969
rect 51724 52003 51776 52012
rect 2688 51824 2740 51876
rect 51724 51969 51733 52003
rect 51733 51969 51767 52003
rect 51767 51969 51776 52003
rect 51724 51960 51776 51969
rect 52184 51960 52236 52012
rect 53196 51960 53248 52012
rect 53840 51960 53892 52012
rect 55036 52003 55088 52012
rect 53104 51935 53156 51944
rect 53104 51901 53113 51935
rect 53113 51901 53147 51935
rect 53147 51901 53156 51935
rect 55036 51969 55045 52003
rect 55045 51969 55079 52003
rect 55079 51969 55088 52003
rect 55036 51960 55088 51969
rect 53104 51892 53156 51901
rect 1584 51799 1636 51808
rect 1584 51765 1593 51799
rect 1593 51765 1627 51799
rect 1627 51765 1636 51799
rect 1584 51756 1636 51765
rect 52092 51799 52144 51808
rect 52092 51765 52101 51799
rect 52101 51765 52135 51799
rect 52135 51765 52144 51799
rect 52092 51756 52144 51765
rect 53840 51756 53892 51808
rect 77944 51935 77996 51944
rect 77944 51901 77953 51935
rect 77953 51901 77987 51935
rect 77987 51901 77996 51935
rect 77944 51892 77996 51901
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 1584 51552 1636 51604
rect 55036 51552 55088 51604
rect 52368 51527 52420 51536
rect 52368 51493 52377 51527
rect 52377 51493 52411 51527
rect 52411 51493 52420 51527
rect 52368 51484 52420 51493
rect 51724 51416 51776 51468
rect 53104 51416 53156 51468
rect 1492 51323 1544 51332
rect 1492 51289 1501 51323
rect 1501 51289 1535 51323
rect 1535 51289 1544 51323
rect 1492 51280 1544 51289
rect 52184 51391 52236 51400
rect 52184 51357 52198 51391
rect 52198 51357 52232 51391
rect 52232 51357 52236 51391
rect 52184 51348 52236 51357
rect 53012 51348 53064 51400
rect 77300 51391 77352 51400
rect 77300 51357 77309 51391
rect 77309 51357 77343 51391
rect 77343 51357 77352 51391
rect 77300 51348 77352 51357
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 1492 50915 1544 50924
rect 1492 50881 1501 50915
rect 1501 50881 1535 50915
rect 1535 50881 1544 50915
rect 1492 50872 1544 50881
rect 53380 50872 53432 50924
rect 53472 50847 53524 50856
rect 53472 50813 53481 50847
rect 53481 50813 53515 50847
rect 53515 50813 53524 50847
rect 53472 50804 53524 50813
rect 77116 50847 77168 50856
rect 77116 50813 77125 50847
rect 77125 50813 77159 50847
rect 77159 50813 77168 50847
rect 77116 50804 77168 50813
rect 77208 50804 77260 50856
rect 50252 50668 50304 50720
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 50252 50507 50304 50516
rect 50252 50473 50261 50507
rect 50261 50473 50295 50507
rect 50295 50473 50304 50507
rect 50252 50464 50304 50473
rect 2504 50328 2556 50380
rect 1492 50235 1544 50244
rect 1492 50201 1501 50235
rect 1501 50201 1535 50235
rect 1535 50201 1544 50235
rect 1492 50192 1544 50201
rect 51816 50396 51868 50448
rect 53380 50439 53432 50448
rect 53380 50405 53389 50439
rect 53389 50405 53423 50439
rect 53423 50405 53432 50439
rect 53380 50396 53432 50405
rect 51172 50260 51224 50312
rect 52736 50260 52788 50312
rect 53472 50260 53524 50312
rect 49792 50124 49844 50176
rect 50988 50235 51040 50244
rect 50988 50201 50997 50235
rect 50997 50201 51031 50235
rect 51031 50201 51040 50235
rect 53012 50235 53064 50244
rect 50988 50192 51040 50201
rect 53012 50201 53021 50235
rect 53021 50201 53055 50235
rect 53055 50201 53064 50235
rect 53012 50192 53064 50201
rect 77392 50260 77444 50312
rect 77576 50303 77628 50312
rect 77576 50269 77585 50303
rect 77585 50269 77619 50303
rect 77619 50269 77628 50303
rect 77576 50260 77628 50269
rect 52736 50124 52788 50176
rect 77208 50192 77260 50244
rect 77760 50124 77812 50176
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 49792 49963 49844 49972
rect 49792 49929 49801 49963
rect 49801 49929 49835 49963
rect 49835 49929 49844 49963
rect 49792 49920 49844 49929
rect 50344 49920 50396 49972
rect 50988 49920 51040 49972
rect 52736 49963 52788 49972
rect 52736 49929 52745 49963
rect 52745 49929 52779 49963
rect 52779 49929 52788 49963
rect 52736 49920 52788 49929
rect 77392 49895 77444 49904
rect 50712 49784 50764 49836
rect 51172 49784 51224 49836
rect 51264 49716 51316 49768
rect 77392 49861 77401 49895
rect 77401 49861 77435 49895
rect 77435 49861 77444 49895
rect 77392 49852 77444 49861
rect 77576 49716 77628 49768
rect 1492 49623 1544 49632
rect 1492 49589 1501 49623
rect 1501 49589 1535 49623
rect 1535 49589 1544 49623
rect 1492 49580 1544 49589
rect 78128 49580 78180 49632
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 50620 49308 50672 49360
rect 1492 49215 1544 49224
rect 1492 49181 1501 49215
rect 1501 49181 1535 49215
rect 1535 49181 1544 49215
rect 1492 49172 1544 49181
rect 50344 49215 50396 49224
rect 50344 49181 50353 49215
rect 50353 49181 50387 49215
rect 50387 49181 50396 49215
rect 50344 49172 50396 49181
rect 50712 49172 50764 49224
rect 78128 49215 78180 49224
rect 78128 49181 78137 49215
rect 78137 49181 78171 49215
rect 78171 49181 78180 49215
rect 78128 49172 78180 49181
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 50160 48832 50212 48884
rect 1492 48739 1544 48748
rect 1492 48705 1501 48739
rect 1501 48705 1535 48739
rect 1535 48705 1544 48739
rect 1492 48696 1544 48705
rect 50712 48696 50764 48748
rect 49976 48492 50028 48544
rect 77116 48671 77168 48680
rect 77116 48637 77125 48671
rect 77125 48637 77159 48671
rect 77159 48637 77168 48671
rect 77116 48628 77168 48637
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 47768 48016 47820 48068
rect 1492 47991 1544 48000
rect 1492 47957 1501 47991
rect 1501 47957 1535 47991
rect 1535 47957 1544 47991
rect 1492 47948 1544 47957
rect 48320 47948 48372 48000
rect 77024 47948 77076 48000
rect 78036 47991 78088 48000
rect 78036 47957 78045 47991
rect 78045 47957 78079 47991
rect 78079 47957 78088 47991
rect 78036 47948 78088 47957
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 47768 47787 47820 47796
rect 47768 47753 47777 47787
rect 47777 47753 47811 47787
rect 47811 47753 47820 47787
rect 47768 47744 47820 47753
rect 47124 47608 47176 47660
rect 48320 47608 48372 47660
rect 49240 47608 49292 47660
rect 77024 47472 77076 47524
rect 1492 47447 1544 47456
rect 1492 47413 1501 47447
rect 1501 47413 1535 47447
rect 1535 47413 1544 47447
rect 1492 47404 1544 47413
rect 49240 47404 49292 47456
rect 69664 47404 69716 47456
rect 77852 47447 77904 47456
rect 77852 47413 77861 47447
rect 77861 47413 77895 47447
rect 77895 47413 77904 47447
rect 77852 47404 77904 47413
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 47124 47243 47176 47252
rect 47124 47209 47133 47243
rect 47133 47209 47167 47243
rect 47167 47209 47176 47243
rect 47124 47200 47176 47209
rect 47676 46996 47728 47048
rect 69664 46928 69716 46980
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 47676 46699 47728 46708
rect 47676 46665 47685 46699
rect 47685 46665 47719 46699
rect 47719 46665 47728 46699
rect 47676 46656 47728 46665
rect 46388 46520 46440 46572
rect 1492 46427 1544 46436
rect 1492 46393 1501 46427
rect 1501 46393 1535 46427
rect 1535 46393 1544 46427
rect 1492 46384 1544 46393
rect 46940 46316 46992 46368
rect 69664 46316 69716 46368
rect 77852 46427 77904 46436
rect 77852 46393 77861 46427
rect 77861 46393 77895 46427
rect 77895 46393 77904 46427
rect 77852 46384 77904 46393
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 46388 46155 46440 46164
rect 46388 46121 46397 46155
rect 46397 46121 46431 46155
rect 46431 46121 46440 46155
rect 46388 46112 46440 46121
rect 46848 45976 46900 46028
rect 46940 45908 46992 45960
rect 47768 45908 47820 45960
rect 1492 45815 1544 45824
rect 1492 45781 1501 45815
rect 1501 45781 1535 45815
rect 1535 45781 1544 45815
rect 1492 45772 1544 45781
rect 2228 45815 2280 45824
rect 2228 45781 2237 45815
rect 2237 45781 2271 45815
rect 2271 45781 2280 45815
rect 2228 45772 2280 45781
rect 69664 45772 69716 45824
rect 78036 45815 78088 45824
rect 78036 45781 78045 45815
rect 78045 45781 78079 45815
rect 78079 45781 78088 45815
rect 78036 45772 78088 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 46848 45543 46900 45552
rect 46848 45509 46857 45543
rect 46857 45509 46891 45543
rect 46891 45509 46900 45543
rect 46848 45500 46900 45509
rect 44916 45432 44968 45484
rect 46664 45475 46716 45484
rect 46664 45441 46673 45475
rect 46673 45441 46707 45475
rect 46707 45441 46716 45475
rect 46664 45432 46716 45441
rect 2228 45296 2280 45348
rect 1492 45271 1544 45280
rect 1492 45237 1501 45271
rect 1501 45237 1535 45271
rect 1535 45237 1544 45271
rect 1492 45228 1544 45237
rect 69664 45228 69716 45280
rect 77852 45271 77904 45280
rect 77852 45237 77861 45271
rect 77861 45237 77895 45271
rect 77895 45237 77904 45271
rect 77852 45228 77904 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 44916 45024 44968 45076
rect 44272 44820 44324 44872
rect 45928 44795 45980 44804
rect 45928 44761 45937 44795
rect 45937 44761 45971 44795
rect 45971 44761 45980 44795
rect 45928 44752 45980 44761
rect 1492 44727 1544 44736
rect 1492 44693 1501 44727
rect 1501 44693 1535 44727
rect 1535 44693 1544 44727
rect 1492 44684 1544 44693
rect 69664 44684 69716 44736
rect 77300 44727 77352 44736
rect 77300 44693 77309 44727
rect 77309 44693 77343 44727
rect 77343 44693 77352 44727
rect 77300 44684 77352 44693
rect 78036 44727 78088 44736
rect 78036 44693 78045 44727
rect 78045 44693 78079 44727
rect 78079 44693 78088 44727
rect 78036 44684 78088 44693
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 44272 44523 44324 44532
rect 44272 44489 44281 44523
rect 44281 44489 44315 44523
rect 44315 44489 44324 44523
rect 44272 44480 44324 44489
rect 45192 44387 45244 44396
rect 45192 44353 45201 44387
rect 45201 44353 45235 44387
rect 45235 44353 45244 44387
rect 45192 44344 45244 44353
rect 45928 44140 45980 44192
rect 77300 44140 77352 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 43536 43732 43588 43784
rect 1492 43639 1544 43648
rect 1492 43605 1501 43639
rect 1501 43605 1535 43639
rect 1535 43605 1544 43639
rect 1492 43596 1544 43605
rect 44272 43596 44324 43648
rect 77300 43639 77352 43648
rect 77300 43605 77309 43639
rect 77309 43605 77343 43639
rect 77343 43605 77352 43639
rect 77300 43596 77352 43605
rect 78036 43639 78088 43648
rect 78036 43605 78045 43639
rect 78045 43605 78079 43639
rect 78079 43605 78088 43639
rect 78036 43596 78088 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 43536 43435 43588 43444
rect 43536 43401 43545 43435
rect 43545 43401 43579 43435
rect 43579 43401 43588 43435
rect 43536 43392 43588 43401
rect 1492 43095 1544 43104
rect 1492 43061 1501 43095
rect 1501 43061 1535 43095
rect 1535 43061 1544 43095
rect 1492 43052 1544 43061
rect 44272 43256 44324 43308
rect 77300 43120 77352 43172
rect 2320 43052 2372 43104
rect 76932 43052 76984 43104
rect 77852 43095 77904 43104
rect 77852 43061 77861 43095
rect 77861 43061 77895 43095
rect 77895 43061 77904 43095
rect 77852 43052 77904 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 2320 42644 2372 42696
rect 42524 42576 42576 42628
rect 1492 42551 1544 42560
rect 1492 42517 1501 42551
rect 1501 42517 1535 42551
rect 1535 42517 1544 42551
rect 1492 42508 1544 42517
rect 44180 42508 44232 42560
rect 76932 42508 76984 42560
rect 77024 42508 77076 42560
rect 78036 42551 78088 42560
rect 78036 42517 78045 42551
rect 78045 42517 78079 42551
rect 78079 42517 78088 42551
rect 78036 42508 78088 42517
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 42524 42347 42576 42356
rect 42524 42313 42533 42347
rect 42533 42313 42567 42347
rect 42567 42313 42576 42347
rect 42524 42304 42576 42313
rect 43352 42168 43404 42220
rect 41328 42032 41380 42084
rect 77024 42032 77076 42084
rect 1492 42007 1544 42016
rect 1492 41973 1501 42007
rect 1501 41973 1535 42007
rect 1535 41973 1544 42007
rect 1492 41964 1544 41973
rect 69664 41964 69716 42016
rect 77852 42007 77904 42016
rect 77852 41973 77861 42007
rect 77861 41973 77895 42007
rect 77895 41973 77904 42007
rect 77852 41964 77904 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 41328 41735 41380 41744
rect 41328 41701 41337 41735
rect 41337 41701 41371 41735
rect 41371 41701 41380 41735
rect 41328 41692 41380 41701
rect 42616 41556 42668 41608
rect 43352 41420 43404 41472
rect 69664 41420 69716 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 1492 40987 1544 40996
rect 1492 40953 1501 40987
rect 1501 40953 1535 40987
rect 1535 40953 1544 40987
rect 1492 40944 1544 40953
rect 40684 40944 40736 40996
rect 77852 40987 77904 40996
rect 77852 40953 77861 40987
rect 77861 40953 77895 40987
rect 77895 40953 77904 40987
rect 77852 40944 77904 40953
rect 41420 40876 41472 40928
rect 42616 40919 42668 40928
rect 42616 40885 42625 40919
rect 42625 40885 42659 40919
rect 42659 40885 42668 40919
rect 42616 40876 42668 40885
rect 77116 40919 77168 40928
rect 77116 40885 77125 40919
rect 77125 40885 77159 40919
rect 77159 40885 77168 40919
rect 77116 40876 77168 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 40684 40715 40736 40724
rect 40684 40681 40693 40715
rect 40693 40681 40727 40715
rect 40727 40681 40736 40715
rect 40684 40672 40736 40681
rect 1492 40375 1544 40384
rect 1492 40341 1501 40375
rect 1501 40341 1535 40375
rect 1535 40341 1544 40375
rect 1492 40332 1544 40341
rect 41420 40400 41472 40452
rect 77116 40400 77168 40452
rect 2320 40332 2372 40384
rect 41052 40332 41104 40384
rect 78036 40375 78088 40384
rect 78036 40341 78045 40375
rect 78045 40341 78079 40375
rect 78079 40341 78088 40375
rect 78036 40332 78088 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 40592 39992 40644 40044
rect 41052 40035 41104 40044
rect 41052 40001 41061 40035
rect 41061 40001 41095 40035
rect 41095 40001 41104 40035
rect 41052 39992 41104 40001
rect 2320 39924 2372 39976
rect 39120 39856 39172 39908
rect 1492 39831 1544 39840
rect 1492 39797 1501 39831
rect 1501 39797 1535 39831
rect 1535 39797 1544 39831
rect 1492 39788 1544 39797
rect 41420 39788 41472 39840
rect 69664 39788 69716 39840
rect 77852 39831 77904 39840
rect 77852 39797 77861 39831
rect 77861 39797 77895 39831
rect 77895 39797 77904 39831
rect 77852 39788 77904 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 39120 39627 39172 39636
rect 39120 39593 39129 39627
rect 39129 39593 39163 39627
rect 39163 39593 39172 39627
rect 39120 39584 39172 39593
rect 38384 39312 38436 39364
rect 39856 39312 39908 39364
rect 1492 39287 1544 39296
rect 1492 39253 1501 39287
rect 1501 39253 1535 39287
rect 1535 39253 1544 39287
rect 1492 39244 1544 39253
rect 40592 39244 40644 39296
rect 69664 39244 69716 39296
rect 77300 39287 77352 39296
rect 77300 39253 77309 39287
rect 77309 39253 77343 39287
rect 77343 39253 77352 39287
rect 77300 39244 77352 39253
rect 78036 39287 78088 39296
rect 78036 39253 78045 39287
rect 78045 39253 78079 39287
rect 78079 39253 78088 39287
rect 78036 39244 78088 39253
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 38384 39040 38436 39092
rect 39120 38904 39172 38956
rect 39856 38700 39908 38752
rect 77300 38700 77352 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 37740 38224 37792 38276
rect 1492 38199 1544 38208
rect 1492 38165 1501 38199
rect 1501 38165 1535 38199
rect 1535 38165 1544 38199
rect 1492 38156 1544 38165
rect 38384 38199 38436 38208
rect 38384 38165 38393 38199
rect 38393 38165 38427 38199
rect 38427 38165 38436 38199
rect 38384 38156 38436 38165
rect 39120 38199 39172 38208
rect 39120 38165 39129 38199
rect 39129 38165 39163 38199
rect 39163 38165 39172 38199
rect 39120 38156 39172 38165
rect 77024 38156 77076 38208
rect 78036 38199 78088 38208
rect 78036 38165 78045 38199
rect 78045 38165 78079 38199
rect 78079 38165 78088 38199
rect 78036 38156 78088 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 37740 37995 37792 38004
rect 37740 37961 37749 37995
rect 37749 37961 37783 37995
rect 37783 37961 37792 37995
rect 37740 37952 37792 37961
rect 38384 37816 38436 37868
rect 37004 37680 37056 37732
rect 77024 37680 77076 37732
rect 1492 37655 1544 37664
rect 1492 37621 1501 37655
rect 1501 37621 1535 37655
rect 1535 37621 1544 37655
rect 1492 37612 1544 37621
rect 69664 37612 69716 37664
rect 77852 37655 77904 37664
rect 77852 37621 77861 37655
rect 77861 37621 77895 37655
rect 77895 37621 77904 37655
rect 77852 37612 77904 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 37004 37451 37056 37460
rect 37004 37417 37013 37451
rect 37013 37417 37047 37451
rect 37047 37417 37056 37451
rect 37004 37408 37056 37417
rect 38384 37340 38436 37392
rect 69664 37272 69716 37324
rect 36268 37136 36320 37188
rect 37648 37136 37700 37188
rect 38016 37136 38068 37188
rect 1492 37111 1544 37120
rect 1492 37077 1501 37111
rect 1501 37077 1535 37111
rect 1535 37077 1544 37111
rect 1492 37068 1544 37077
rect 77300 37111 77352 37120
rect 77300 37077 77309 37111
rect 77309 37077 77343 37111
rect 77343 37077 77352 37111
rect 77300 37068 77352 37077
rect 78036 37111 78088 37120
rect 78036 37077 78045 37111
rect 78045 37077 78079 37111
rect 78079 37077 78088 37111
rect 78036 37068 78088 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 36268 36907 36320 36916
rect 36268 36873 36277 36907
rect 36277 36873 36311 36907
rect 36311 36873 36320 36907
rect 36268 36864 36320 36873
rect 38016 36907 38068 36916
rect 38016 36873 38025 36907
rect 38025 36873 38059 36907
rect 38059 36873 38068 36907
rect 38016 36864 38068 36873
rect 35624 36728 35676 36780
rect 36636 36728 36688 36780
rect 37188 36728 37240 36780
rect 77300 36796 77352 36848
rect 1492 36567 1544 36576
rect 1492 36533 1501 36567
rect 1501 36533 1535 36567
rect 1535 36533 1544 36567
rect 1492 36524 1544 36533
rect 69664 36524 69716 36576
rect 77852 36567 77904 36576
rect 77852 36533 77861 36567
rect 77861 36533 77895 36567
rect 77895 36533 77904 36567
rect 77852 36524 77904 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 35624 36363 35676 36372
rect 35624 36329 35633 36363
rect 35633 36329 35667 36363
rect 35667 36329 35676 36363
rect 35624 36320 35676 36329
rect 37188 36363 37240 36372
rect 37188 36329 37197 36363
rect 37197 36329 37231 36363
rect 37231 36329 37240 36363
rect 37188 36320 37240 36329
rect 36268 36048 36320 36100
rect 69664 35980 69716 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 1492 35547 1544 35556
rect 1492 35513 1501 35547
rect 1501 35513 1535 35547
rect 1535 35513 1544 35547
rect 1492 35504 1544 35513
rect 34704 35504 34756 35556
rect 35716 35436 35768 35488
rect 36268 35479 36320 35488
rect 36268 35445 36277 35479
rect 36277 35445 36311 35479
rect 36311 35445 36320 35479
rect 36268 35436 36320 35445
rect 68008 35436 68060 35488
rect 77852 35547 77904 35556
rect 77852 35513 77861 35547
rect 77861 35513 77895 35547
rect 77895 35513 77904 35547
rect 77852 35504 77904 35513
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 34704 35232 34756 35284
rect 34152 35028 34204 35080
rect 34796 34960 34848 35012
rect 35716 34960 35768 35012
rect 1492 34935 1544 34944
rect 1492 34901 1501 34935
rect 1501 34901 1535 34935
rect 1535 34901 1544 34935
rect 1492 34892 1544 34901
rect 68008 34892 68060 34944
rect 77300 34935 77352 34944
rect 77300 34901 77309 34935
rect 77309 34901 77343 34935
rect 77343 34901 77352 34935
rect 77300 34892 77352 34901
rect 78036 34935 78088 34944
rect 78036 34901 78045 34935
rect 78045 34901 78079 34935
rect 78079 34901 78088 34935
rect 78036 34892 78088 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 34152 34731 34204 34740
rect 34152 34697 34161 34731
rect 34161 34697 34195 34731
rect 34195 34697 34204 34731
rect 34152 34688 34204 34697
rect 35716 34731 35768 34740
rect 35716 34697 35725 34731
rect 35725 34697 35759 34731
rect 35759 34697 35768 34731
rect 35716 34688 35768 34697
rect 77300 34620 77352 34672
rect 34704 34552 34756 34604
rect 2320 34484 2372 34536
rect 77116 34527 77168 34536
rect 77116 34493 77125 34527
rect 77125 34493 77159 34527
rect 77159 34493 77168 34527
rect 77116 34484 77168 34493
rect 1492 34391 1544 34400
rect 1492 34357 1501 34391
rect 1501 34357 1535 34391
rect 1535 34357 1544 34391
rect 1492 34348 1544 34357
rect 77852 34391 77904 34400
rect 77852 34357 77861 34391
rect 77861 34357 77895 34391
rect 77895 34357 77904 34391
rect 77852 34348 77904 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 2320 33940 2372 33992
rect 32680 33872 32732 33924
rect 1492 33847 1544 33856
rect 1492 33813 1501 33847
rect 1501 33813 1535 33847
rect 1535 33813 1544 33847
rect 1492 33804 1544 33813
rect 33968 33804 34020 33856
rect 34704 33804 34756 33856
rect 77116 33804 77168 33856
rect 77300 33847 77352 33856
rect 77300 33813 77309 33847
rect 77309 33813 77343 33847
rect 77343 33813 77352 33847
rect 77300 33804 77352 33813
rect 78036 33847 78088 33856
rect 78036 33813 78045 33847
rect 78045 33813 78079 33847
rect 78079 33813 78088 33847
rect 78036 33804 78088 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 32680 33643 32732 33652
rect 32680 33609 32689 33643
rect 32689 33609 32723 33643
rect 32723 33609 32732 33643
rect 32680 33600 32732 33609
rect 33232 33464 33284 33516
rect 77300 33260 77352 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 32220 32784 32272 32836
rect 1492 32759 1544 32768
rect 1492 32725 1501 32759
rect 1501 32725 1535 32759
rect 1535 32725 1544 32759
rect 1492 32716 1544 32725
rect 32956 32716 33008 32768
rect 33232 32716 33284 32768
rect 77024 32716 77076 32768
rect 78036 32759 78088 32768
rect 78036 32725 78045 32759
rect 78045 32725 78079 32759
rect 78079 32725 78088 32759
rect 78036 32716 78088 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 32220 32555 32272 32564
rect 32220 32521 32229 32555
rect 32229 32521 32263 32555
rect 32263 32521 32272 32555
rect 32220 32512 32272 32521
rect 31208 32376 31260 32428
rect 32956 32419 33008 32428
rect 32956 32385 32965 32419
rect 32965 32385 32999 32419
rect 32999 32385 33008 32419
rect 32956 32376 33008 32385
rect 77024 32240 77076 32292
rect 1492 32215 1544 32224
rect 1492 32181 1501 32215
rect 1501 32181 1535 32215
rect 1535 32181 1544 32215
rect 1492 32172 1544 32181
rect 69664 32172 69716 32224
rect 77852 32215 77904 32224
rect 77852 32181 77861 32215
rect 77861 32181 77895 32215
rect 77895 32181 77904 32215
rect 77852 32172 77904 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 31208 32011 31260 32020
rect 31208 31977 31217 32011
rect 31217 31977 31251 32011
rect 31251 31977 31260 32011
rect 31208 31968 31260 31977
rect 32404 31900 32456 31952
rect 78036 31943 78088 31952
rect 69664 31832 69716 31884
rect 2320 31764 2372 31816
rect 32588 31764 32640 31816
rect 32956 31807 33008 31816
rect 32956 31773 32965 31807
rect 32965 31773 32999 31807
rect 32999 31773 33008 31807
rect 32956 31764 33008 31773
rect 78036 31909 78045 31943
rect 78045 31909 78079 31943
rect 78079 31909 78088 31943
rect 78036 31900 78088 31909
rect 31944 31696 31996 31748
rect 1492 31671 1544 31680
rect 1492 31637 1501 31671
rect 1501 31637 1535 31671
rect 1535 31637 1544 31671
rect 1492 31628 1544 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 32404 31399 32456 31408
rect 32404 31365 32413 31399
rect 32413 31365 32447 31399
rect 32447 31365 32456 31399
rect 32404 31356 32456 31365
rect 31668 31288 31720 31340
rect 2320 31220 2372 31272
rect 29736 31152 29788 31204
rect 1492 31127 1544 31136
rect 1492 31093 1501 31127
rect 1501 31093 1535 31127
rect 1535 31093 1544 31127
rect 1492 31084 1544 31093
rect 31944 31084 31996 31136
rect 68008 31084 68060 31136
rect 77852 31127 77904 31136
rect 77852 31093 77861 31127
rect 77861 31093 77895 31127
rect 77895 31093 77904 31127
rect 77852 31084 77904 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 29736 30923 29788 30932
rect 29736 30889 29745 30923
rect 29745 30889 29779 30923
rect 29779 30889 29788 30923
rect 29736 30880 29788 30889
rect 30380 30608 30432 30660
rect 31024 30540 31076 30592
rect 31668 30540 31720 30592
rect 68008 30540 68060 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 1492 30107 1544 30116
rect 1492 30073 1501 30107
rect 1501 30073 1535 30107
rect 1535 30073 1544 30107
rect 1492 30064 1544 30073
rect 28816 30064 28868 30116
rect 29368 29996 29420 30048
rect 30380 29996 30432 30048
rect 69664 29996 69716 30048
rect 77852 30107 77904 30116
rect 77852 30073 77861 30107
rect 77861 30073 77895 30107
rect 77895 30073 77904 30107
rect 77852 30064 77904 30073
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 28816 29835 28868 29844
rect 28816 29801 28825 29835
rect 28825 29801 28859 29835
rect 28859 29801 28868 29835
rect 28816 29792 28868 29801
rect 28264 29588 28316 29640
rect 1492 29495 1544 29504
rect 1492 29461 1501 29495
rect 1501 29461 1535 29495
rect 1535 29461 1544 29495
rect 1492 29452 1544 29461
rect 29368 29452 29420 29504
rect 69664 29452 69716 29504
rect 77300 29495 77352 29504
rect 77300 29461 77309 29495
rect 77309 29461 77343 29495
rect 77343 29461 77352 29495
rect 77300 29452 77352 29461
rect 78036 29495 78088 29504
rect 78036 29461 78045 29495
rect 78045 29461 78079 29495
rect 78079 29461 78088 29495
rect 78036 29452 78088 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 28264 29291 28316 29300
rect 28264 29257 28273 29291
rect 28273 29257 28307 29291
rect 28307 29257 28316 29291
rect 28264 29248 28316 29257
rect 26148 29044 26200 29096
rect 77300 29112 77352 29164
rect 1492 29019 1544 29028
rect 1492 28985 1501 29019
rect 1501 28985 1535 29019
rect 1535 28985 1544 29019
rect 1492 28976 1544 28985
rect 28724 28976 28776 29028
rect 77116 29019 77168 29028
rect 77116 28985 77125 29019
rect 77125 28985 77159 29019
rect 77159 28985 77168 29019
rect 77116 28976 77168 28985
rect 77852 29019 77904 29028
rect 77852 28985 77861 29019
rect 77861 28985 77895 29019
rect 77895 28985 77904 29019
rect 77852 28976 77904 28985
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 26148 28636 26200 28688
rect 27068 28500 27120 28552
rect 1492 28407 1544 28416
rect 1492 28373 1501 28407
rect 1501 28373 1535 28407
rect 1535 28373 1544 28407
rect 1492 28364 1544 28373
rect 27988 28364 28040 28416
rect 77116 28364 77168 28416
rect 77300 28407 77352 28416
rect 77300 28373 77309 28407
rect 77309 28373 77343 28407
rect 77343 28373 77352 28407
rect 77300 28364 77352 28373
rect 78036 28407 78088 28416
rect 78036 28373 78045 28407
rect 78045 28373 78079 28407
rect 78079 28373 78088 28407
rect 78036 28364 78088 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 27068 28203 27120 28212
rect 27068 28169 27077 28203
rect 27077 28169 27111 28203
rect 27111 28169 27120 28203
rect 27068 28160 27120 28169
rect 27436 28024 27488 28076
rect 77300 27820 77352 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 26056 27412 26108 27464
rect 1492 27319 1544 27328
rect 1492 27285 1501 27319
rect 1501 27285 1535 27319
rect 1535 27285 1544 27319
rect 1492 27276 1544 27285
rect 26148 27276 26200 27328
rect 27436 27319 27488 27328
rect 27436 27285 27445 27319
rect 27445 27285 27479 27319
rect 27479 27285 27488 27319
rect 27436 27276 27488 27285
rect 77024 27276 77076 27328
rect 78036 27319 78088 27328
rect 78036 27285 78045 27319
rect 78045 27285 78079 27319
rect 78079 27285 78088 27319
rect 78036 27276 78088 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 26056 27115 26108 27124
rect 26056 27081 26065 27115
rect 26065 27081 26099 27115
rect 26099 27081 26108 27115
rect 26056 27072 26108 27081
rect 25228 26936 25280 26988
rect 26148 26979 26200 26988
rect 26148 26945 26157 26979
rect 26157 26945 26191 26979
rect 26191 26945 26200 26979
rect 26148 26936 26200 26945
rect 77024 26800 77076 26852
rect 1492 26775 1544 26784
rect 1492 26741 1501 26775
rect 1501 26741 1535 26775
rect 1535 26741 1544 26775
rect 1492 26732 1544 26741
rect 69664 26732 69716 26784
rect 77852 26775 77904 26784
rect 77852 26741 77861 26775
rect 77861 26741 77895 26775
rect 77895 26741 77904 26775
rect 77852 26732 77904 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 25228 26571 25280 26580
rect 25228 26537 25237 26571
rect 25237 26537 25271 26571
rect 25271 26537 25280 26571
rect 25228 26528 25280 26537
rect 78036 26503 78088 26512
rect 78036 26469 78045 26503
rect 78045 26469 78079 26503
rect 78079 26469 78088 26503
rect 78036 26460 78088 26469
rect 26148 26392 26200 26444
rect 22836 26324 22888 26376
rect 77392 26367 77444 26376
rect 1492 26231 1544 26240
rect 1492 26197 1501 26231
rect 1501 26197 1535 26231
rect 1535 26197 1544 26231
rect 1492 26188 1544 26197
rect 77392 26333 77401 26367
rect 77401 26333 77435 26367
rect 77435 26333 77444 26367
rect 77392 26324 77444 26333
rect 69664 26256 69716 26308
rect 26056 26231 26108 26240
rect 26056 26197 26065 26231
rect 26065 26197 26099 26231
rect 26099 26197 26108 26231
rect 26056 26188 26108 26197
rect 32680 26188 32732 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 22836 25959 22888 25968
rect 22836 25925 22845 25959
rect 22845 25925 22879 25959
rect 22879 25925 22888 25959
rect 22836 25916 22888 25925
rect 31668 25916 31720 25968
rect 32680 25959 32732 25968
rect 32680 25925 32689 25959
rect 32689 25925 32723 25959
rect 32723 25925 32732 25959
rect 32680 25916 32732 25925
rect 24952 25848 25004 25900
rect 22284 25712 22336 25764
rect 69664 25712 69716 25764
rect 1492 25687 1544 25696
rect 1492 25653 1501 25687
rect 1501 25653 1535 25687
rect 1535 25653 1544 25687
rect 1492 25644 1544 25653
rect 26056 25644 26108 25696
rect 77392 25644 77444 25696
rect 77852 25687 77904 25696
rect 77852 25653 77861 25687
rect 77861 25653 77895 25687
rect 77895 25653 77904 25687
rect 77852 25644 77904 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 22284 25483 22336 25492
rect 22284 25449 22293 25483
rect 22293 25449 22327 25483
rect 22327 25449 22336 25483
rect 22284 25440 22336 25449
rect 24400 25236 24452 25288
rect 30840 25100 30892 25152
rect 69664 25100 69716 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 24400 24828 24452 24880
rect 30840 24828 30892 24880
rect 22284 24760 22336 24812
rect 41512 24760 41564 24812
rect 1492 24667 1544 24676
rect 1492 24633 1501 24667
rect 1501 24633 1535 24667
rect 1535 24633 1544 24667
rect 1492 24624 1544 24633
rect 41696 24624 41748 24676
rect 60464 24624 60516 24676
rect 41604 24599 41656 24608
rect 41604 24565 41613 24599
rect 41613 24565 41647 24599
rect 41647 24565 41656 24599
rect 41604 24556 41656 24565
rect 69664 24556 69716 24608
rect 77852 24667 77904 24676
rect 77852 24633 77861 24667
rect 77861 24633 77895 24667
rect 77895 24633 77904 24667
rect 77852 24624 77904 24633
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 22284 24395 22336 24404
rect 22284 24361 22293 24395
rect 22293 24361 22327 24395
rect 22327 24361 22336 24395
rect 22284 24352 22336 24361
rect 41604 24352 41656 24404
rect 21824 24148 21876 24200
rect 23664 24080 23716 24132
rect 32036 24123 32088 24132
rect 32036 24089 32045 24123
rect 32045 24089 32079 24123
rect 32079 24089 32088 24123
rect 32036 24080 32088 24089
rect 41512 24123 41564 24132
rect 41512 24089 41521 24123
rect 41521 24089 41555 24123
rect 41555 24089 41564 24123
rect 41512 24080 41564 24089
rect 1492 24055 1544 24064
rect 1492 24021 1501 24055
rect 1501 24021 1535 24055
rect 1535 24021 1544 24055
rect 1492 24012 1544 24021
rect 41696 24055 41748 24064
rect 41696 24021 41705 24055
rect 41705 24021 41739 24055
rect 41739 24021 41748 24055
rect 41696 24012 41748 24021
rect 61200 24080 61252 24132
rect 69664 24012 69716 24064
rect 77300 24055 77352 24064
rect 77300 24021 77309 24055
rect 77309 24021 77343 24055
rect 77343 24021 77352 24055
rect 77300 24012 77352 24021
rect 78036 24055 78088 24064
rect 78036 24021 78045 24055
rect 78045 24021 78079 24055
rect 78079 24021 78088 24055
rect 78036 24012 78088 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 21824 23851 21876 23860
rect 21824 23817 21833 23851
rect 21833 23817 21867 23851
rect 21867 23817 21876 23851
rect 21824 23808 21876 23817
rect 30840 23851 30892 23860
rect 30840 23817 30849 23851
rect 30849 23817 30883 23851
rect 30883 23817 30892 23851
rect 30840 23808 30892 23817
rect 31576 23808 31628 23860
rect 22560 23672 22612 23724
rect 31392 23715 31444 23724
rect 31392 23681 31401 23715
rect 31401 23681 31435 23715
rect 31435 23681 31444 23715
rect 31392 23672 31444 23681
rect 31484 23672 31536 23724
rect 32220 23715 32272 23724
rect 32220 23681 32229 23715
rect 32229 23681 32263 23715
rect 32263 23681 32272 23715
rect 32220 23672 32272 23681
rect 37188 23672 37240 23724
rect 41696 23715 41748 23724
rect 41696 23681 41705 23715
rect 41705 23681 41739 23715
rect 41739 23681 41748 23715
rect 41696 23672 41748 23681
rect 77116 23672 77168 23724
rect 77300 23604 77352 23656
rect 19708 23536 19760 23588
rect 41604 23536 41656 23588
rect 1492 23511 1544 23520
rect 1492 23477 1501 23511
rect 1501 23477 1535 23511
rect 1535 23477 1544 23511
rect 1492 23468 1544 23477
rect 22560 23511 22612 23520
rect 22560 23477 22569 23511
rect 22569 23477 22603 23511
rect 22603 23477 22612 23511
rect 22560 23468 22612 23477
rect 41512 23468 41564 23520
rect 77116 23511 77168 23520
rect 77116 23477 77125 23511
rect 77125 23477 77159 23511
rect 77159 23477 77168 23511
rect 77116 23468 77168 23477
rect 77852 23511 77904 23520
rect 77852 23477 77861 23511
rect 77861 23477 77895 23511
rect 77895 23477 77904 23511
rect 77852 23468 77904 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 19708 23307 19760 23316
rect 19708 23273 19717 23307
rect 19717 23273 19751 23307
rect 19751 23273 19760 23307
rect 19708 23264 19760 23273
rect 24952 23264 25004 23316
rect 30288 23264 30340 23316
rect 31484 23264 31536 23316
rect 31576 23307 31628 23316
rect 31576 23273 31585 23307
rect 31585 23273 31619 23307
rect 31619 23273 31628 23307
rect 31576 23264 31628 23273
rect 77116 23128 77168 23180
rect 19984 22992 20036 23044
rect 1492 22967 1544 22976
rect 1492 22933 1501 22967
rect 1501 22933 1535 22967
rect 1535 22933 1544 22967
rect 1492 22924 1544 22933
rect 22560 23060 22612 23112
rect 22928 23060 22980 23112
rect 31668 23060 31720 23112
rect 32036 23103 32088 23112
rect 32036 23069 32045 23103
rect 32045 23069 32079 23103
rect 32079 23069 32088 23103
rect 32036 23060 32088 23069
rect 27160 22967 27212 22976
rect 27160 22933 27169 22967
rect 27169 22933 27203 22967
rect 27203 22933 27212 22967
rect 32220 22992 32272 23044
rect 27160 22924 27212 22933
rect 30288 22924 30340 22976
rect 31668 22924 31720 22976
rect 77300 22967 77352 22976
rect 77300 22933 77309 22967
rect 77309 22933 77343 22967
rect 77343 22933 77352 22967
rect 77300 22924 77352 22933
rect 78036 22967 78088 22976
rect 78036 22933 78045 22967
rect 78045 22933 78079 22967
rect 78079 22933 78088 22967
rect 78036 22924 78088 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 19984 22763 20036 22772
rect 19984 22729 19993 22763
rect 19993 22729 20027 22763
rect 20027 22729 20036 22763
rect 19984 22720 20036 22729
rect 32036 22720 32088 22772
rect 26976 22380 27028 22432
rect 77300 22448 77352 22500
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 19064 21972 19116 22024
rect 27344 21904 27396 21956
rect 1492 21879 1544 21888
rect 1492 21845 1501 21879
rect 1501 21845 1535 21879
rect 1535 21845 1544 21879
rect 1492 21836 1544 21845
rect 78036 21879 78088 21888
rect 78036 21845 78045 21879
rect 78045 21845 78079 21879
rect 78079 21845 78088 21879
rect 78036 21836 78088 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 19064 21675 19116 21684
rect 19064 21641 19073 21675
rect 19073 21641 19107 21675
rect 19107 21641 19116 21675
rect 19064 21632 19116 21641
rect 17868 21496 17920 21548
rect 1492 21335 1544 21344
rect 1492 21301 1501 21335
rect 1501 21301 1535 21335
rect 1535 21301 1544 21335
rect 1492 21292 1544 21301
rect 20352 21292 20404 21344
rect 77116 21335 77168 21344
rect 77116 21301 77125 21335
rect 77125 21301 77159 21335
rect 77159 21301 77168 21335
rect 77116 21292 77168 21301
rect 77852 21335 77904 21344
rect 77852 21301 77861 21335
rect 77861 21301 77895 21335
rect 77895 21301 77904 21335
rect 77852 21292 77904 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 17868 21131 17920 21140
rect 17868 21097 17877 21131
rect 17877 21097 17911 21131
rect 17911 21097 17920 21131
rect 17868 21088 17920 21097
rect 17960 20884 18012 20936
rect 19432 20884 19484 20936
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 32404 20884 32456 20936
rect 27068 20748 27120 20800
rect 77116 20748 77168 20800
rect 78036 20791 78088 20800
rect 78036 20757 78045 20791
rect 78045 20757 78079 20791
rect 78079 20757 78088 20791
rect 78036 20748 78088 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 17960 20544 18012 20596
rect 32404 20519 32456 20528
rect 32404 20485 32413 20519
rect 32413 20485 32447 20519
rect 32447 20485 32456 20519
rect 32404 20476 32456 20485
rect 17040 20408 17092 20460
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 31484 20408 31536 20460
rect 19340 20204 19392 20256
rect 31484 20247 31536 20256
rect 31484 20213 31493 20247
rect 31493 20213 31527 20247
rect 31527 20213 31536 20247
rect 31484 20204 31536 20213
rect 68008 20204 68060 20256
rect 77852 20247 77904 20256
rect 77852 20213 77861 20247
rect 77861 20213 77895 20247
rect 77895 20213 77904 20247
rect 77852 20204 77904 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 17040 20043 17092 20052
rect 17040 20009 17049 20043
rect 17049 20009 17083 20043
rect 17083 20009 17092 20043
rect 17040 20000 17092 20009
rect 17960 19660 18012 19712
rect 30932 19703 30984 19712
rect 30932 19669 30941 19703
rect 30941 19669 30975 19703
rect 30975 19669 30984 19703
rect 30932 19660 30984 19669
rect 68008 19660 68060 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 77852 19499 77904 19508
rect 77852 19465 77861 19499
rect 77861 19465 77895 19499
rect 77895 19465 77904 19499
rect 77852 19456 77904 19465
rect 1492 19227 1544 19236
rect 1492 19193 1501 19227
rect 1501 19193 1535 19227
rect 1535 19193 1544 19227
rect 1492 19184 1544 19193
rect 17960 19320 18012 19372
rect 18512 19320 18564 19372
rect 30932 19320 30984 19372
rect 31760 19320 31812 19372
rect 17776 19116 17828 19168
rect 31760 19116 31812 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 19340 18640 19392 18692
rect 30472 18640 30524 18692
rect 31392 18912 31444 18964
rect 30656 18776 30708 18828
rect 31484 18776 31536 18828
rect 30932 18708 30984 18760
rect 31760 18708 31812 18760
rect 16856 18615 16908 18624
rect 16856 18581 16865 18615
rect 16865 18581 16899 18615
rect 16899 18581 16908 18615
rect 16856 18572 16908 18581
rect 26332 18615 26384 18624
rect 26332 18581 26341 18615
rect 26341 18581 26375 18615
rect 26375 18581 26384 18615
rect 26332 18572 26384 18581
rect 27068 18572 27120 18624
rect 30564 18615 30616 18624
rect 30564 18581 30573 18615
rect 30573 18581 30607 18615
rect 30607 18581 30616 18615
rect 30564 18572 30616 18581
rect 78036 18615 78088 18624
rect 78036 18581 78045 18615
rect 78045 18581 78079 18615
rect 78079 18581 78088 18615
rect 78036 18572 78088 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 16856 18368 16908 18420
rect 17040 18368 17092 18420
rect 30564 18368 30616 18420
rect 12348 18232 12400 18284
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 20352 18028 20404 18080
rect 31760 18300 31812 18352
rect 26516 18232 26568 18284
rect 26976 18232 27028 18284
rect 27344 18275 27396 18284
rect 27344 18241 27353 18275
rect 27353 18241 27387 18275
rect 27387 18241 27396 18275
rect 27344 18232 27396 18241
rect 77116 18232 77168 18284
rect 27160 18207 27212 18216
rect 27160 18173 27169 18207
rect 27169 18173 27203 18207
rect 27203 18173 27212 18207
rect 27160 18164 27212 18173
rect 26332 18096 26384 18148
rect 27068 18071 27120 18080
rect 27068 18037 27077 18071
rect 27077 18037 27111 18071
rect 27111 18037 27120 18071
rect 27068 18028 27120 18037
rect 27712 18028 27764 18080
rect 77116 18071 77168 18080
rect 77116 18037 77125 18071
rect 77125 18037 77159 18071
rect 77159 18037 77168 18071
rect 77116 18028 77168 18037
rect 77852 18071 77904 18080
rect 77852 18037 77861 18071
rect 77861 18037 77895 18071
rect 77895 18037 77904 18071
rect 77852 18028 77904 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 12348 17824 12400 17876
rect 27712 17731 27764 17740
rect 27712 17697 27721 17731
rect 27721 17697 27755 17731
rect 27755 17697 27764 17731
rect 27712 17688 27764 17697
rect 14464 17620 14516 17672
rect 27344 17663 27396 17672
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 27344 17629 27353 17663
rect 27353 17629 27387 17663
rect 27387 17629 27396 17663
rect 27344 17620 27396 17629
rect 27528 17663 27580 17672
rect 27528 17629 27537 17663
rect 27537 17629 27571 17663
rect 27571 17629 27580 17663
rect 27528 17620 27580 17629
rect 15936 17484 15988 17536
rect 26424 17484 26476 17536
rect 26516 17527 26568 17536
rect 26516 17493 26525 17527
rect 26525 17493 26559 17527
rect 26559 17493 26568 17527
rect 26516 17484 26568 17493
rect 37188 17484 37240 17536
rect 77024 17484 77076 17536
rect 78036 17527 78088 17536
rect 78036 17493 78045 17527
rect 78045 17493 78079 17527
rect 78079 17493 78088 17527
rect 78036 17484 78088 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 14464 17323 14516 17332
rect 14464 17289 14473 17323
rect 14473 17289 14507 17323
rect 14507 17289 14516 17323
rect 14464 17280 14516 17289
rect 26424 17187 26476 17196
rect 15108 16940 15160 16992
rect 26424 17153 26433 17187
rect 26433 17153 26467 17187
rect 26467 17153 26476 17187
rect 26424 17144 26476 17153
rect 26240 16940 26292 16992
rect 28172 16983 28224 16992
rect 28172 16949 28181 16983
rect 28181 16949 28215 16983
rect 28215 16949 28224 16983
rect 28172 16940 28224 16949
rect 77116 16940 77168 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 26424 16736 26476 16788
rect 77024 16600 77076 16652
rect 12716 16532 12768 16584
rect 28172 16532 28224 16584
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 26240 16396 26292 16448
rect 78036 16439 78088 16448
rect 78036 16405 78045 16439
rect 78045 16405 78079 16439
rect 78079 16405 78088 16439
rect 78036 16396 78088 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 12716 16235 12768 16244
rect 12716 16201 12725 16235
rect 12725 16201 12759 16235
rect 12759 16201 12768 16235
rect 12716 16192 12768 16201
rect 26240 16192 26292 16244
rect 27528 16192 27580 16244
rect 14096 16056 14148 16108
rect 27620 16124 27672 16176
rect 28172 16124 28224 16176
rect 13820 15988 13872 16040
rect 26424 15988 26476 16040
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 14096 15895 14148 15904
rect 14096 15861 14105 15895
rect 14105 15861 14139 15895
rect 14139 15861 14148 15895
rect 14096 15852 14148 15861
rect 27712 15852 27764 15904
rect 77852 15895 77904 15904
rect 77852 15861 77861 15895
rect 77861 15861 77895 15895
rect 77895 15861 77904 15895
rect 77852 15852 77904 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 14096 15648 14148 15700
rect 27712 15691 27764 15700
rect 27712 15657 27721 15691
rect 27721 15657 27755 15691
rect 27755 15657 27764 15691
rect 27712 15648 27764 15657
rect 11520 15444 11572 15496
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 13820 15308 13872 15360
rect 14464 15308 14516 15360
rect 27620 15580 27672 15632
rect 27804 15376 27856 15428
rect 78036 15351 78088 15360
rect 78036 15317 78045 15351
rect 78045 15317 78079 15351
rect 78079 15317 78088 15351
rect 78036 15308 78088 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 11520 15147 11572 15156
rect 11520 15113 11529 15147
rect 11529 15113 11563 15147
rect 11563 15113 11572 15147
rect 11520 15104 11572 15113
rect 27804 15036 27856 15088
rect 11520 14968 11572 15020
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 27068 14968 27120 15020
rect 13360 14764 13412 14816
rect 68008 14764 68060 14816
rect 77852 14807 77904 14816
rect 77852 14773 77861 14807
rect 77861 14773 77895 14807
rect 77895 14773 77904 14807
rect 77852 14764 77904 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 11520 14603 11572 14612
rect 11520 14569 11529 14603
rect 11529 14569 11563 14603
rect 11563 14569 11572 14603
rect 11520 14560 11572 14569
rect 26976 14288 27028 14340
rect 12624 14220 12676 14272
rect 68008 14220 68060 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 12624 14016 12676 14068
rect 26976 14016 27028 14068
rect 27344 14059 27396 14068
rect 27344 14025 27353 14059
rect 27353 14025 27387 14059
rect 27387 14025 27396 14059
rect 27344 14016 27396 14025
rect 77852 14059 77904 14068
rect 77852 14025 77861 14059
rect 77861 14025 77895 14059
rect 77895 14025 77904 14059
rect 77852 14016 77904 14025
rect 13360 13880 13412 13932
rect 11888 13812 11940 13864
rect 27068 13923 27120 13932
rect 27068 13889 27077 13923
rect 27077 13889 27111 13923
rect 27111 13889 27120 13923
rect 27896 13923 27948 13932
rect 27068 13880 27120 13889
rect 27896 13889 27905 13923
rect 27905 13889 27939 13923
rect 27939 13889 27948 13923
rect 27896 13880 27948 13889
rect 1492 13787 1544 13796
rect 1492 13753 1501 13787
rect 1501 13753 1535 13787
rect 1535 13753 1544 13787
rect 1492 13744 1544 13753
rect 26976 13719 27028 13728
rect 26976 13685 26985 13719
rect 26985 13685 27019 13719
rect 27019 13685 27028 13719
rect 26976 13676 27028 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 26976 13472 27028 13524
rect 27896 13472 27948 13524
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 10784 13200 10836 13252
rect 41512 13175 41564 13184
rect 41512 13141 41521 13175
rect 41521 13141 41555 13175
rect 41555 13141 41564 13175
rect 41512 13132 41564 13141
rect 78036 13175 78088 13184
rect 78036 13141 78045 13175
rect 78045 13141 78079 13175
rect 78079 13141 78088 13175
rect 78036 13132 78088 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 9680 12792 9732 12844
rect 77116 12792 77168 12844
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 77116 12631 77168 12640
rect 77116 12597 77125 12631
rect 77125 12597 77159 12631
rect 77159 12597 77168 12631
rect 77116 12588 77168 12597
rect 77852 12631 77904 12640
rect 77852 12597 77861 12631
rect 77861 12597 77895 12631
rect 77895 12597 77904 12631
rect 77852 12588 77904 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 9036 12180 9088 12232
rect 10048 12180 10100 12232
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 77116 12044 77168 12096
rect 77300 12087 77352 12096
rect 77300 12053 77309 12087
rect 77309 12053 77343 12087
rect 77343 12053 77352 12087
rect 77300 12044 77352 12053
rect 78036 12087 78088 12096
rect 78036 12053 78045 12087
rect 78045 12053 78079 12087
rect 78079 12053 78088 12087
rect 78036 12044 78088 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9588 11704 9640 11756
rect 77300 11500 77352 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 1492 11271 1544 11280
rect 1492 11237 1501 11271
rect 1501 11237 1535 11271
rect 1535 11237 1544 11271
rect 1492 11228 1544 11237
rect 78036 11271 78088 11280
rect 78036 11237 78045 11271
rect 78045 11237 78079 11271
rect 78079 11237 78088 11271
rect 78036 11228 78088 11237
rect 8300 11092 8352 11144
rect 11704 11024 11756 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 7564 10616 7616 10668
rect 8944 10616 8996 10668
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 77116 10455 77168 10464
rect 77116 10421 77125 10455
rect 77125 10421 77159 10455
rect 77159 10421 77168 10455
rect 77116 10412 77168 10421
rect 77852 10455 77904 10464
rect 77852 10421 77861 10455
rect 77861 10421 77895 10455
rect 77895 10421 77904 10455
rect 77852 10412 77904 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 7564 10251 7616 10260
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 6736 10004 6788 10056
rect 8208 10004 8260 10056
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 77116 9936 77168 9988
rect 10968 9868 11020 9920
rect 78036 9911 78088 9920
rect 78036 9877 78045 9911
rect 78045 9877 78079 9911
rect 78079 9877 78088 9911
rect 78036 9868 78088 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 6736 9707 6788 9716
rect 6736 9673 6745 9707
rect 6745 9673 6779 9707
rect 6779 9673 6788 9707
rect 6736 9664 6788 9673
rect 10968 9664 11020 9716
rect 6000 9528 6052 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 69664 9324 69716 9376
rect 77852 9367 77904 9376
rect 77852 9333 77861 9367
rect 77861 9333 77895 9367
rect 77895 9333 77904 9367
rect 77852 9324 77904 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 6000 9163 6052 9172
rect 6000 9129 6009 9163
rect 6009 9129 6043 9163
rect 6043 9129 6052 9163
rect 6000 9120 6052 9129
rect 6184 8959 6236 8968
rect 6184 8925 6193 8959
rect 6193 8925 6227 8959
rect 6227 8925 6236 8959
rect 6184 8916 6236 8925
rect 69664 8780 69716 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 5264 8440 5316 8492
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 77116 8347 77168 8356
rect 77116 8313 77125 8347
rect 77125 8313 77159 8347
rect 77159 8313 77168 8347
rect 77116 8304 77168 8313
rect 77852 8347 77904 8356
rect 77852 8313 77861 8347
rect 77861 8313 77895 8347
rect 77895 8313 77904 8347
rect 77852 8304 77904 8313
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 4528 7828 4580 7880
rect 5632 7828 5684 7880
rect 77024 7760 77076 7812
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 77116 7692 77168 7744
rect 78036 7735 78088 7744
rect 78036 7701 78045 7735
rect 78045 7701 78079 7735
rect 78079 7701 78088 7735
rect 78036 7692 78088 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 3884 7352 3936 7404
rect 4712 7395 4764 7404
rect 4712 7361 4721 7395
rect 4721 7361 4755 7395
rect 4755 7361 4764 7395
rect 4712 7352 4764 7361
rect 77024 7216 77076 7268
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 76012 7148 76064 7200
rect 77852 7191 77904 7200
rect 77852 7157 77861 7191
rect 77861 7157 77895 7191
rect 77895 7157 77904 7191
rect 77852 7148 77904 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 3884 6987 3936 6996
rect 3884 6953 3893 6987
rect 3893 6953 3927 6987
rect 3927 6953 3936 6987
rect 3884 6944 3936 6953
rect 3240 6740 3292 6792
rect 4620 6740 4672 6792
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 76012 6604 76064 6656
rect 77300 6647 77352 6656
rect 77300 6613 77309 6647
rect 77309 6613 77343 6647
rect 77343 6613 77352 6647
rect 77300 6604 77352 6613
rect 78036 6647 78088 6656
rect 78036 6613 78045 6647
rect 78045 6613 78079 6647
rect 78079 6613 78088 6647
rect 78036 6604 78088 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 3240 6443 3292 6452
rect 3240 6409 3249 6443
rect 3249 6409 3283 6443
rect 3283 6409 3292 6443
rect 3240 6400 3292 6409
rect 3792 6264 3844 6316
rect 77300 6060 77352 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 6644 5652 6696 5704
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 78036 5559 78088 5568
rect 78036 5525 78045 5559
rect 78045 5525 78079 5559
rect 78079 5525 78088 5559
rect 78036 5516 78088 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 1676 5312 1728 5364
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 2044 5176 2096 5228
rect 3056 5176 3108 5228
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 69664 4972 69716 5024
rect 77852 5015 77904 5024
rect 77852 4981 77861 5015
rect 77861 4981 77895 5015
rect 77895 4981 77904 5015
rect 77852 4972 77904 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 2044 4811 2096 4820
rect 2044 4777 2053 4811
rect 2053 4777 2087 4811
rect 2087 4777 2096 4811
rect 2044 4768 2096 4777
rect 2320 4564 2372 4616
rect 69664 4428 69716 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 53840 3723 53892 3732
rect 53840 3689 53849 3723
rect 53849 3689 53883 3723
rect 53883 3689 53892 3723
rect 53840 3680 53892 3689
rect 64328 3723 64380 3732
rect 64328 3689 64337 3723
rect 64337 3689 64371 3723
rect 64371 3689 64380 3723
rect 64328 3680 64380 3689
rect 27528 3544 27580 3596
rect 63868 3544 63920 3596
rect 69664 3544 69716 3596
rect 27068 3476 27120 3528
rect 29276 3408 29328 3460
rect 66168 3408 66220 3460
rect 70584 3408 70636 3460
rect 28448 3383 28500 3392
rect 28448 3349 28457 3383
rect 28457 3349 28491 3383
rect 28491 3349 28500 3383
rect 28448 3340 28500 3349
rect 30012 3383 30064 3392
rect 30012 3349 30021 3383
rect 30021 3349 30055 3383
rect 30055 3349 30064 3383
rect 30012 3340 30064 3349
rect 32220 3383 32272 3392
rect 32220 3349 32229 3383
rect 32229 3349 32263 3383
rect 32263 3349 32272 3383
rect 32220 3340 32272 3349
rect 32956 3383 33008 3392
rect 32956 3349 32965 3383
rect 32965 3349 32999 3383
rect 32999 3349 33008 3383
rect 32956 3340 33008 3349
rect 33692 3383 33744 3392
rect 33692 3349 33701 3383
rect 33701 3349 33735 3383
rect 33735 3349 33744 3383
rect 33692 3340 33744 3349
rect 43720 3383 43772 3392
rect 43720 3349 43729 3383
rect 43729 3349 43763 3383
rect 43763 3349 43772 3383
rect 43720 3340 43772 3349
rect 74724 3383 74776 3392
rect 74724 3349 74733 3383
rect 74733 3349 74767 3383
rect 74767 3349 74776 3383
rect 74724 3340 74776 3349
rect 77852 3340 77904 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 3792 3179 3844 3188
rect 3792 3145 3801 3179
rect 3801 3145 3835 3179
rect 3835 3145 3844 3179
rect 3792 3136 3844 3145
rect 8944 3179 8996 3188
rect 8944 3145 8953 3179
rect 8953 3145 8987 3179
rect 8987 3145 8996 3179
rect 8944 3136 8996 3145
rect 14096 3179 14148 3188
rect 14096 3145 14105 3179
rect 14105 3145 14139 3179
rect 14139 3145 14148 3179
rect 14096 3136 14148 3145
rect 24400 3179 24452 3188
rect 24400 3145 24409 3179
rect 24409 3145 24443 3179
rect 24443 3145 24452 3179
rect 24400 3136 24452 3145
rect 32496 3179 32548 3188
rect 32496 3145 32505 3179
rect 32505 3145 32539 3179
rect 32539 3145 32548 3179
rect 32496 3136 32548 3145
rect 33232 3179 33284 3188
rect 33232 3145 33241 3179
rect 33241 3145 33275 3179
rect 33275 3145 33284 3179
rect 33232 3136 33284 3145
rect 34704 3179 34756 3188
rect 34704 3145 34713 3179
rect 34713 3145 34747 3179
rect 34747 3145 34756 3179
rect 34704 3136 34756 3145
rect 39856 3179 39908 3188
rect 39856 3145 39865 3179
rect 39865 3145 39899 3179
rect 39899 3145 39908 3179
rect 39856 3136 39908 3145
rect 44272 3179 44324 3188
rect 44272 3145 44281 3179
rect 44281 3145 44315 3179
rect 44315 3145 44324 3179
rect 44272 3136 44324 3145
rect 49976 3179 50028 3188
rect 49976 3145 49985 3179
rect 49985 3145 50019 3179
rect 50019 3145 50028 3179
rect 49976 3136 50028 3145
rect 50620 3179 50672 3188
rect 50620 3145 50629 3179
rect 50629 3145 50663 3179
rect 50663 3145 50672 3179
rect 50620 3136 50672 3145
rect 51264 3179 51316 3188
rect 51264 3145 51273 3179
rect 51273 3145 51307 3179
rect 51307 3145 51316 3179
rect 51264 3136 51316 3145
rect 51816 3179 51868 3188
rect 51816 3145 51825 3179
rect 51825 3145 51859 3179
rect 51859 3145 51868 3179
rect 51816 3136 51868 3145
rect 52368 3136 52420 3188
rect 53288 3179 53340 3188
rect 53288 3145 53297 3179
rect 53297 3145 53331 3179
rect 53331 3145 53340 3179
rect 53288 3136 53340 3145
rect 55404 3136 55456 3188
rect 56600 3136 56652 3188
rect 57152 3179 57204 3188
rect 57152 3145 57161 3179
rect 57161 3145 57195 3179
rect 57195 3145 57204 3179
rect 57152 3136 57204 3145
rect 58440 3179 58492 3188
rect 58440 3145 58449 3179
rect 58449 3145 58483 3179
rect 58483 3145 58492 3179
rect 58440 3136 58492 3145
rect 58992 3179 59044 3188
rect 58992 3145 59001 3179
rect 59001 3145 59035 3179
rect 59035 3145 59044 3179
rect 58992 3136 59044 3145
rect 60280 3179 60332 3188
rect 60280 3145 60289 3179
rect 60289 3145 60323 3179
rect 60323 3145 60332 3179
rect 60280 3136 60332 3145
rect 60648 3136 60700 3188
rect 63316 3136 63368 3188
rect 19340 3111 19392 3120
rect 19340 3077 19349 3111
rect 19349 3077 19383 3111
rect 19383 3077 19392 3111
rect 19340 3068 19392 3077
rect 3516 3000 3568 3052
rect 8668 3000 8720 3052
rect 13820 3000 13872 3052
rect 18972 3000 19024 3052
rect 24124 3000 24176 3052
rect 26056 3000 26108 3052
rect 27988 3000 28040 3052
rect 29368 3043 29420 3052
rect 29368 3009 29377 3043
rect 29377 3009 29411 3043
rect 29411 3009 29420 3043
rect 29368 3000 29420 3009
rect 30380 3043 30432 3052
rect 30380 3009 30389 3043
rect 30389 3009 30423 3043
rect 30423 3009 30432 3043
rect 30380 3000 30432 3009
rect 32220 3000 32272 3052
rect 32956 3000 33008 3052
rect 34428 3000 34480 3052
rect 39580 3000 39632 3052
rect 43996 3000 44048 3052
rect 52092 3068 52144 3120
rect 57060 3068 57112 3120
rect 57888 3068 57940 3120
rect 60556 3068 60608 3120
rect 62396 3068 62448 3120
rect 63408 3068 63460 3120
rect 65248 3136 65300 3188
rect 66168 3136 66220 3188
rect 69296 3179 69348 3188
rect 69296 3145 69305 3179
rect 69305 3145 69339 3179
rect 69339 3145 69348 3179
rect 69296 3136 69348 3145
rect 70584 3179 70636 3188
rect 70584 3145 70593 3179
rect 70593 3145 70627 3179
rect 70627 3145 70636 3179
rect 70584 3136 70636 3145
rect 72056 3179 72108 3188
rect 72056 3145 72065 3179
rect 72065 3145 72099 3179
rect 72099 3145 72108 3179
rect 72056 3136 72108 3145
rect 75920 3136 75972 3188
rect 65064 3068 65116 3120
rect 68192 3111 68244 3120
rect 68192 3077 68201 3111
rect 68201 3077 68235 3111
rect 68235 3077 68244 3111
rect 68192 3068 68244 3077
rect 65156 3000 65208 3052
rect 68928 3000 68980 3052
rect 25596 2932 25648 2984
rect 27804 2932 27856 2984
rect 28448 2932 28500 2984
rect 29276 2932 29328 2984
rect 30012 2932 30064 2984
rect 59912 2932 59964 2984
rect 61936 2975 61988 2984
rect 61936 2941 61945 2975
rect 61945 2941 61979 2975
rect 61979 2941 61988 2975
rect 61936 2932 61988 2941
rect 62488 2932 62540 2984
rect 65432 2975 65484 2984
rect 65432 2941 65441 2975
rect 65441 2941 65475 2975
rect 65475 2941 65484 2975
rect 65432 2932 65484 2941
rect 65524 2932 65576 2984
rect 74908 3000 74960 3052
rect 77852 3000 77904 3052
rect 62304 2864 62356 2916
rect 66352 2864 66404 2916
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 4988 2796 5040 2848
rect 5724 2839 5776 2848
rect 5724 2805 5733 2839
rect 5733 2805 5767 2839
rect 5767 2805 5776 2839
rect 5724 2796 5776 2805
rect 6460 2839 6512 2848
rect 6460 2805 6469 2839
rect 6469 2805 6503 2839
rect 6503 2805 6512 2839
rect 6460 2796 6512 2805
rect 7196 2839 7248 2848
rect 7196 2805 7205 2839
rect 7205 2805 7239 2839
rect 7239 2805 7248 2839
rect 7196 2796 7248 2805
rect 7932 2796 7984 2848
rect 9404 2796 9456 2848
rect 10140 2796 10192 2848
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 11612 2839 11664 2848
rect 11612 2805 11621 2839
rect 11621 2805 11655 2839
rect 11655 2805 11664 2839
rect 11612 2796 11664 2805
rect 12348 2839 12400 2848
rect 12348 2805 12357 2839
rect 12357 2805 12391 2839
rect 12391 2805 12400 2839
rect 12348 2796 12400 2805
rect 13084 2796 13136 2848
rect 14556 2796 14608 2848
rect 15292 2796 15344 2848
rect 16028 2839 16080 2848
rect 16028 2805 16037 2839
rect 16037 2805 16071 2839
rect 16071 2805 16080 2839
rect 16028 2796 16080 2805
rect 16764 2839 16816 2848
rect 16764 2805 16773 2839
rect 16773 2805 16807 2839
rect 16807 2805 16816 2839
rect 16764 2796 16816 2805
rect 17500 2839 17552 2848
rect 17500 2805 17509 2839
rect 17509 2805 17543 2839
rect 17543 2805 17552 2839
rect 17500 2796 17552 2805
rect 18236 2796 18288 2848
rect 19984 2839 20036 2848
rect 19984 2805 19993 2839
rect 19993 2805 20027 2839
rect 20027 2805 20036 2839
rect 19984 2796 20036 2805
rect 20444 2796 20496 2848
rect 21180 2839 21232 2848
rect 21180 2805 21189 2839
rect 21189 2805 21223 2839
rect 21223 2805 21232 2839
rect 21180 2796 21232 2805
rect 21916 2839 21968 2848
rect 21916 2805 21925 2839
rect 21925 2805 21959 2839
rect 21959 2805 21968 2839
rect 21916 2796 21968 2805
rect 22652 2839 22704 2848
rect 22652 2805 22661 2839
rect 22661 2805 22695 2839
rect 22695 2805 22704 2839
rect 22652 2796 22704 2805
rect 23388 2796 23440 2848
rect 24860 2796 24912 2848
rect 31484 2839 31536 2848
rect 31484 2805 31493 2839
rect 31493 2805 31527 2839
rect 31527 2805 31536 2839
rect 31484 2796 31536 2805
rect 35348 2839 35400 2848
rect 35348 2805 35357 2839
rect 35357 2805 35391 2839
rect 35391 2805 35400 2839
rect 35348 2796 35400 2805
rect 35900 2796 35952 2848
rect 36636 2839 36688 2848
rect 36636 2805 36645 2839
rect 36645 2805 36679 2839
rect 36679 2805 36688 2839
rect 36636 2796 36688 2805
rect 37372 2839 37424 2848
rect 37372 2805 37381 2839
rect 37381 2805 37415 2839
rect 37415 2805 37424 2839
rect 37372 2796 37424 2805
rect 38108 2839 38160 2848
rect 38108 2805 38117 2839
rect 38117 2805 38151 2839
rect 38151 2805 38160 2839
rect 38108 2796 38160 2805
rect 38844 2796 38896 2848
rect 41052 2839 41104 2848
rect 41052 2805 41061 2839
rect 41061 2805 41095 2839
rect 41095 2805 41104 2839
rect 41052 2796 41104 2805
rect 42432 2839 42484 2848
rect 42432 2805 42441 2839
rect 42441 2805 42475 2839
rect 42475 2805 42484 2839
rect 42432 2796 42484 2805
rect 42800 2796 42852 2848
rect 44732 2796 44784 2848
rect 45652 2839 45704 2848
rect 45652 2805 45661 2839
rect 45661 2805 45695 2839
rect 45695 2805 45704 2839
rect 45652 2796 45704 2805
rect 46204 2796 46256 2848
rect 47584 2839 47636 2848
rect 47584 2805 47593 2839
rect 47593 2805 47627 2839
rect 47627 2805 47636 2839
rect 47584 2796 47636 2805
rect 47676 2796 47728 2848
rect 48412 2796 48464 2848
rect 48780 2839 48832 2848
rect 48780 2805 48789 2839
rect 48789 2805 48823 2839
rect 48823 2805 48832 2839
rect 48780 2796 48832 2805
rect 49148 2796 49200 2848
rect 54300 2796 54352 2848
rect 59452 2796 59504 2848
rect 59820 2796 59872 2848
rect 63040 2839 63092 2848
rect 63040 2805 63049 2839
rect 63049 2805 63083 2839
rect 63083 2805 63092 2839
rect 63040 2796 63092 2805
rect 64604 2796 64656 2848
rect 66076 2796 66128 2848
rect 71504 2864 71556 2916
rect 77116 2907 77168 2916
rect 77116 2873 77125 2907
rect 77125 2873 77159 2907
rect 77159 2873 77168 2907
rect 77116 2864 77168 2873
rect 77392 2864 77444 2916
rect 69756 2796 69808 2848
rect 73344 2839 73396 2848
rect 73344 2805 73353 2839
rect 73353 2805 73387 2839
rect 73387 2805 73396 2839
rect 73344 2796 73396 2805
rect 73896 2839 73948 2848
rect 73896 2805 73905 2839
rect 73905 2805 73939 2839
rect 73939 2805 73948 2839
rect 73896 2796 73948 2805
rect 75736 2839 75788 2848
rect 75736 2805 75745 2839
rect 75745 2805 75779 2839
rect 75779 2805 75788 2839
rect 75736 2796 75788 2805
rect 76380 2796 76432 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 4620 2592 4672 2644
rect 4712 2592 4764 2644
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 6184 2592 6236 2644
rect 6920 2592 6972 2644
rect 8208 2635 8260 2644
rect 8208 2601 8217 2635
rect 8217 2601 8251 2635
rect 8251 2601 8260 2635
rect 8208 2592 8260 2601
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 11888 2635 11940 2644
rect 11888 2601 11897 2635
rect 11897 2601 11931 2635
rect 11931 2601 11940 2635
rect 11888 2592 11940 2601
rect 12624 2635 12676 2644
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 13360 2635 13412 2644
rect 13360 2601 13369 2635
rect 13369 2601 13403 2635
rect 13403 2601 13412 2635
rect 13360 2592 13412 2601
rect 14464 2635 14516 2644
rect 14464 2601 14473 2635
rect 14473 2601 14507 2635
rect 14507 2601 14516 2635
rect 14464 2592 14516 2601
rect 15936 2635 15988 2644
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 17040 2635 17092 2644
rect 17040 2601 17049 2635
rect 17049 2601 17083 2635
rect 17083 2601 17092 2635
rect 17040 2592 17092 2601
rect 17776 2635 17828 2644
rect 17776 2601 17785 2635
rect 17785 2601 17819 2635
rect 17819 2601 17828 2635
rect 17776 2592 17828 2601
rect 18512 2635 18564 2644
rect 18512 2601 18521 2635
rect 18521 2601 18555 2635
rect 18555 2601 18564 2635
rect 18512 2592 18564 2601
rect 20352 2635 20404 2644
rect 20352 2601 20361 2635
rect 20361 2601 20395 2635
rect 20395 2601 20404 2635
rect 20352 2592 20404 2601
rect 22928 2635 22980 2644
rect 22928 2601 22937 2635
rect 22937 2601 22971 2635
rect 22971 2601 22980 2635
rect 22928 2592 22980 2601
rect 23664 2635 23716 2644
rect 23664 2601 23673 2635
rect 23673 2601 23707 2635
rect 23707 2601 23716 2635
rect 23664 2592 23716 2601
rect 24952 2635 25004 2644
rect 24952 2601 24961 2635
rect 24961 2601 24995 2635
rect 24995 2601 25004 2635
rect 24952 2592 25004 2601
rect 33968 2635 34020 2644
rect 33968 2601 33977 2635
rect 33977 2601 34011 2635
rect 34011 2601 34020 2635
rect 33968 2592 34020 2601
rect 36268 2592 36320 2644
rect 36544 2635 36596 2644
rect 36544 2601 36553 2635
rect 36553 2601 36587 2635
rect 36587 2601 36596 2635
rect 36544 2592 36596 2601
rect 37648 2635 37700 2644
rect 37648 2601 37657 2635
rect 37657 2601 37691 2635
rect 37691 2601 37700 2635
rect 37648 2592 37700 2601
rect 38384 2635 38436 2644
rect 38384 2601 38393 2635
rect 38393 2601 38427 2635
rect 38427 2601 38436 2635
rect 38384 2592 38436 2601
rect 39120 2635 39172 2644
rect 39120 2601 39129 2635
rect 39129 2601 39163 2635
rect 39163 2601 39172 2635
rect 39120 2592 39172 2601
rect 40592 2635 40644 2644
rect 40592 2601 40601 2635
rect 40601 2601 40635 2635
rect 40635 2601 40644 2635
rect 40592 2592 40644 2601
rect 42616 2635 42668 2644
rect 42616 2601 42625 2635
rect 42625 2601 42659 2635
rect 42659 2601 42668 2635
rect 42616 2592 42668 2601
rect 43352 2635 43404 2644
rect 43352 2601 43361 2635
rect 43361 2601 43395 2635
rect 43395 2601 43404 2635
rect 43352 2592 43404 2601
rect 45192 2635 45244 2644
rect 45192 2601 45201 2635
rect 45201 2601 45235 2635
rect 45235 2601 45244 2635
rect 45192 2592 45244 2601
rect 45928 2635 45980 2644
rect 45928 2601 45937 2635
rect 45937 2601 45971 2635
rect 45971 2601 45980 2635
rect 45928 2592 45980 2601
rect 46664 2635 46716 2644
rect 46664 2601 46673 2635
rect 46673 2601 46707 2635
rect 46707 2601 46716 2635
rect 46664 2592 46716 2601
rect 47768 2635 47820 2644
rect 47768 2601 47777 2635
rect 47777 2601 47811 2635
rect 47811 2601 47820 2635
rect 47768 2592 47820 2601
rect 49240 2635 49292 2644
rect 49240 2601 49249 2635
rect 49249 2601 49283 2635
rect 49283 2601 49292 2635
rect 49240 2592 49292 2601
rect 73528 2635 73580 2644
rect 73528 2601 73537 2635
rect 73537 2601 73571 2635
rect 73571 2601 73580 2635
rect 73528 2592 73580 2601
rect 74264 2635 74316 2644
rect 74264 2601 74273 2635
rect 74273 2601 74307 2635
rect 74307 2601 74316 2635
rect 74264 2592 74316 2601
rect 75000 2635 75052 2644
rect 75000 2601 75009 2635
rect 75009 2601 75043 2635
rect 75043 2601 75052 2635
rect 75000 2592 75052 2601
rect 76288 2592 76340 2644
rect 15108 2567 15160 2576
rect 15108 2533 15117 2567
rect 15117 2533 15151 2567
rect 15151 2533 15160 2567
rect 15108 2524 15160 2533
rect 19432 2524 19484 2576
rect 26332 2524 26384 2576
rect 34796 2524 34848 2576
rect 41420 2567 41472 2576
rect 41420 2533 41429 2567
rect 41429 2533 41463 2567
rect 41463 2533 41472 2567
rect 41420 2524 41472 2533
rect 44180 2567 44232 2576
rect 44180 2533 44189 2567
rect 44189 2533 44223 2567
rect 44223 2533 44232 2567
rect 44180 2524 44232 2533
rect 47492 2524 47544 2576
rect 52828 2524 52880 2576
rect 57980 2524 58032 2576
rect 63868 2524 63920 2576
rect 69020 2524 69072 2576
rect 26148 2499 26200 2508
rect 26148 2465 26157 2499
rect 26157 2465 26191 2499
rect 26191 2465 26200 2499
rect 26148 2456 26200 2465
rect 28724 2499 28776 2508
rect 28724 2465 28733 2499
rect 28733 2465 28767 2499
rect 28767 2465 28776 2499
rect 28724 2456 28776 2465
rect 31024 2499 31076 2508
rect 31024 2465 31033 2499
rect 31033 2465 31067 2499
rect 31067 2465 31076 2499
rect 31024 2456 31076 2465
rect 31944 2456 31996 2508
rect 53288 2456 53340 2508
rect 2044 2388 2096 2440
rect 2780 2388 2832 2440
rect 4252 2388 4304 2440
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 5724 2388 5776 2440
rect 6460 2388 6512 2440
rect 7196 2388 7248 2440
rect 7932 2388 7984 2440
rect 9404 2431 9456 2440
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 10140 2388 10192 2440
rect 10876 2388 10928 2440
rect 22100 2431 22152 2440
rect 22100 2397 22109 2431
rect 22109 2397 22143 2431
rect 22143 2397 22152 2431
rect 22100 2388 22152 2397
rect 23480 2388 23532 2440
rect 26332 2388 26384 2440
rect 28540 2388 28592 2440
rect 30748 2431 30800 2440
rect 30748 2397 30757 2431
rect 30757 2397 30791 2431
rect 30791 2397 30800 2431
rect 30748 2388 30800 2397
rect 31484 2388 31536 2440
rect 45652 2388 45704 2440
rect 48412 2431 48464 2440
rect 48412 2397 48421 2431
rect 48421 2397 48455 2431
rect 48455 2397 48464 2431
rect 48412 2388 48464 2397
rect 50620 2388 50672 2440
rect 51264 2388 51316 2440
rect 51816 2388 51868 2440
rect 52368 2388 52420 2440
rect 53840 2388 53892 2440
rect 60556 2456 60608 2508
rect 55404 2388 55456 2440
rect 56600 2388 56652 2440
rect 57152 2388 57204 2440
rect 57888 2431 57940 2440
rect 57888 2397 57897 2431
rect 57897 2397 57931 2431
rect 57931 2397 57940 2431
rect 57888 2388 57940 2397
rect 58440 2388 58492 2440
rect 58992 2388 59044 2440
rect 60648 2388 60700 2440
rect 66168 2456 66220 2508
rect 61936 2431 61988 2440
rect 61936 2397 61945 2431
rect 61945 2397 61979 2431
rect 61979 2397 61988 2431
rect 61936 2388 61988 2397
rect 63040 2431 63092 2440
rect 63040 2397 63049 2431
rect 63049 2397 63083 2431
rect 63083 2397 63092 2431
rect 63040 2388 63092 2397
rect 63408 2388 63460 2440
rect 64328 2388 64380 2440
rect 65432 2388 65484 2440
rect 66352 2431 66404 2440
rect 66352 2397 66361 2431
rect 66361 2397 66395 2431
rect 66395 2397 66404 2431
rect 66352 2388 66404 2397
rect 68192 2431 68244 2440
rect 68192 2397 68201 2431
rect 68201 2397 68235 2431
rect 68235 2397 68244 2431
rect 68192 2388 68244 2397
rect 68928 2431 68980 2440
rect 68928 2397 68937 2431
rect 68937 2397 68971 2431
rect 68971 2397 68980 2431
rect 68928 2388 68980 2397
rect 69664 2431 69716 2440
rect 69664 2397 69673 2431
rect 69673 2397 69707 2431
rect 69707 2397 69716 2431
rect 69664 2388 69716 2397
rect 70584 2388 70636 2440
rect 71504 2431 71556 2440
rect 71504 2397 71513 2431
rect 71513 2397 71547 2431
rect 71547 2397 71556 2431
rect 71504 2388 71556 2397
rect 72056 2388 72108 2440
rect 72700 2388 72752 2440
rect 73344 2431 73396 2440
rect 73344 2397 73353 2431
rect 73353 2397 73387 2431
rect 73387 2397 73396 2431
rect 73344 2388 73396 2397
rect 73436 2388 73488 2440
rect 73896 2388 73948 2440
rect 74724 2388 74776 2440
rect 75920 2431 75972 2440
rect 75920 2397 75929 2431
rect 75929 2397 75963 2431
rect 75963 2397 75972 2431
rect 75920 2388 75972 2397
rect 76380 2388 76432 2440
rect 77392 2431 77444 2440
rect 77392 2397 77401 2431
rect 77401 2397 77435 2431
rect 77435 2397 77444 2431
rect 77392 2388 77444 2397
rect 11612 2320 11664 2372
rect 12440 2320 12492 2372
rect 13084 2320 13136 2372
rect 14556 2363 14608 2372
rect 14556 2329 14565 2363
rect 14565 2329 14599 2363
rect 14599 2329 14608 2363
rect 14556 2320 14608 2329
rect 15292 2363 15344 2372
rect 15292 2329 15301 2363
rect 15301 2329 15335 2363
rect 15335 2329 15344 2363
rect 15292 2320 15344 2329
rect 16028 2363 16080 2372
rect 16028 2329 16037 2363
rect 16037 2329 16071 2363
rect 16071 2329 16080 2363
rect 16028 2320 16080 2329
rect 16764 2320 16816 2372
rect 17500 2320 17552 2372
rect 18236 2320 18288 2372
rect 19984 2320 20036 2372
rect 20444 2363 20496 2372
rect 20444 2329 20453 2363
rect 20453 2329 20487 2363
rect 20487 2329 20496 2363
rect 20444 2320 20496 2329
rect 21180 2363 21232 2372
rect 21180 2329 21189 2363
rect 21189 2329 21223 2363
rect 21223 2329 21232 2363
rect 21180 2320 21232 2329
rect 22652 2320 22704 2372
rect 24860 2320 24912 2372
rect 33692 2320 33744 2372
rect 35164 2363 35216 2372
rect 35164 2329 35173 2363
rect 35173 2329 35207 2363
rect 35207 2329 35216 2363
rect 35164 2320 35216 2329
rect 35900 2363 35952 2372
rect 35900 2329 35909 2363
rect 35909 2329 35943 2363
rect 35943 2329 35952 2363
rect 36636 2363 36688 2372
rect 35900 2320 35952 2329
rect 36636 2329 36645 2363
rect 36645 2329 36679 2363
rect 36679 2329 36688 2363
rect 36636 2320 36688 2329
rect 37372 2320 37424 2372
rect 38108 2320 38160 2372
rect 38844 2320 38896 2372
rect 40316 2320 40368 2372
rect 41052 2320 41104 2372
rect 41788 2320 41840 2372
rect 42432 2320 42484 2372
rect 42800 2320 42852 2372
rect 43352 2320 43404 2372
rect 43720 2320 43772 2372
rect 44732 2320 44784 2372
rect 46204 2320 46256 2372
rect 46940 2320 46992 2372
rect 47584 2320 47636 2372
rect 48780 2320 48832 2372
rect 67364 2320 67416 2372
rect 26516 2252 26568 2304
rect 48412 2252 48464 2304
rect 49884 2252 49936 2304
rect 50620 2252 50672 2304
rect 51356 2252 51408 2304
rect 52092 2252 52144 2304
rect 53564 2252 53616 2304
rect 55036 2252 55088 2304
rect 55772 2252 55824 2304
rect 56508 2252 56560 2304
rect 57244 2252 57296 2304
rect 58716 2252 58768 2304
rect 60188 2252 60240 2304
rect 60924 2252 60976 2304
rect 61660 2252 61712 2304
rect 62396 2252 62448 2304
rect 63408 2252 63460 2304
rect 65340 2252 65392 2304
rect 66076 2252 66128 2304
rect 66812 2252 66864 2304
rect 67548 2252 67600 2304
rect 68560 2252 68612 2304
rect 70492 2252 70544 2304
rect 71228 2252 71280 2304
rect 71964 2252 72016 2304
rect 77116 2252 77168 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
<< metal2 >>
rect 4214 77820 4522 77829
rect 4214 77818 4220 77820
rect 4276 77818 4300 77820
rect 4356 77818 4380 77820
rect 4436 77818 4460 77820
rect 4516 77818 4522 77820
rect 4276 77766 4278 77818
rect 4458 77766 4460 77818
rect 4214 77764 4220 77766
rect 4276 77764 4300 77766
rect 4356 77764 4380 77766
rect 4436 77764 4460 77766
rect 4516 77764 4522 77766
rect 4214 77755 4522 77764
rect 34934 77820 35242 77829
rect 34934 77818 34940 77820
rect 34996 77818 35020 77820
rect 35076 77818 35100 77820
rect 35156 77818 35180 77820
rect 35236 77818 35242 77820
rect 34996 77766 34998 77818
rect 35178 77766 35180 77818
rect 34934 77764 34940 77766
rect 34996 77764 35020 77766
rect 35076 77764 35100 77766
rect 35156 77764 35180 77766
rect 35236 77764 35242 77766
rect 34934 77755 35242 77764
rect 65654 77820 65962 77829
rect 65654 77818 65660 77820
rect 65716 77818 65740 77820
rect 65796 77818 65820 77820
rect 65876 77818 65900 77820
rect 65956 77818 65962 77820
rect 65716 77766 65718 77818
rect 65898 77766 65900 77818
rect 65654 77764 65660 77766
rect 65716 77764 65740 77766
rect 65796 77764 65820 77766
rect 65876 77764 65900 77766
rect 65956 77764 65962 77766
rect 65654 77755 65962 77764
rect 19574 77276 19882 77285
rect 19574 77274 19580 77276
rect 19636 77274 19660 77276
rect 19716 77274 19740 77276
rect 19796 77274 19820 77276
rect 19876 77274 19882 77276
rect 19636 77222 19638 77274
rect 19818 77222 19820 77274
rect 19574 77220 19580 77222
rect 19636 77220 19660 77222
rect 19716 77220 19740 77222
rect 19796 77220 19820 77222
rect 19876 77220 19882 77222
rect 19574 77211 19882 77220
rect 50294 77276 50602 77285
rect 50294 77274 50300 77276
rect 50356 77274 50380 77276
rect 50436 77274 50460 77276
rect 50516 77274 50540 77276
rect 50596 77274 50602 77276
rect 50356 77222 50358 77274
rect 50538 77222 50540 77274
rect 50294 77220 50300 77222
rect 50356 77220 50380 77222
rect 50436 77220 50460 77222
rect 50516 77220 50540 77222
rect 50596 77220 50602 77222
rect 50294 77211 50602 77220
rect 4214 76732 4522 76741
rect 4214 76730 4220 76732
rect 4276 76730 4300 76732
rect 4356 76730 4380 76732
rect 4436 76730 4460 76732
rect 4516 76730 4522 76732
rect 4276 76678 4278 76730
rect 4458 76678 4460 76730
rect 4214 76676 4220 76678
rect 4276 76676 4300 76678
rect 4356 76676 4380 76678
rect 4436 76676 4460 76678
rect 4516 76676 4522 76678
rect 4214 76667 4522 76676
rect 34934 76732 35242 76741
rect 34934 76730 34940 76732
rect 34996 76730 35020 76732
rect 35076 76730 35100 76732
rect 35156 76730 35180 76732
rect 35236 76730 35242 76732
rect 34996 76678 34998 76730
rect 35178 76678 35180 76730
rect 34934 76676 34940 76678
rect 34996 76676 35020 76678
rect 35076 76676 35100 76678
rect 35156 76676 35180 76678
rect 35236 76676 35242 76678
rect 34934 76667 35242 76676
rect 65654 76732 65962 76741
rect 65654 76730 65660 76732
rect 65716 76730 65740 76732
rect 65796 76730 65820 76732
rect 65876 76730 65900 76732
rect 65956 76730 65962 76732
rect 65716 76678 65718 76730
rect 65898 76678 65900 76730
rect 65654 76676 65660 76678
rect 65716 76676 65740 76678
rect 65796 76676 65820 76678
rect 65876 76676 65900 76678
rect 65956 76676 65962 76678
rect 65654 76667 65962 76676
rect 19574 76188 19882 76197
rect 19574 76186 19580 76188
rect 19636 76186 19660 76188
rect 19716 76186 19740 76188
rect 19796 76186 19820 76188
rect 19876 76186 19882 76188
rect 19636 76134 19638 76186
rect 19818 76134 19820 76186
rect 19574 76132 19580 76134
rect 19636 76132 19660 76134
rect 19716 76132 19740 76134
rect 19796 76132 19820 76134
rect 19876 76132 19882 76134
rect 19574 76123 19882 76132
rect 50294 76188 50602 76197
rect 50294 76186 50300 76188
rect 50356 76186 50380 76188
rect 50436 76186 50460 76188
rect 50516 76186 50540 76188
rect 50596 76186 50602 76188
rect 50356 76134 50358 76186
rect 50538 76134 50540 76186
rect 50294 76132 50300 76134
rect 50356 76132 50380 76134
rect 50436 76132 50460 76134
rect 50516 76132 50540 76134
rect 50596 76132 50602 76134
rect 50294 76123 50602 76132
rect 4214 75644 4522 75653
rect 4214 75642 4220 75644
rect 4276 75642 4300 75644
rect 4356 75642 4380 75644
rect 4436 75642 4460 75644
rect 4516 75642 4522 75644
rect 4276 75590 4278 75642
rect 4458 75590 4460 75642
rect 4214 75588 4220 75590
rect 4276 75588 4300 75590
rect 4356 75588 4380 75590
rect 4436 75588 4460 75590
rect 4516 75588 4522 75590
rect 4214 75579 4522 75588
rect 34934 75644 35242 75653
rect 34934 75642 34940 75644
rect 34996 75642 35020 75644
rect 35076 75642 35100 75644
rect 35156 75642 35180 75644
rect 35236 75642 35242 75644
rect 34996 75590 34998 75642
rect 35178 75590 35180 75642
rect 34934 75588 34940 75590
rect 34996 75588 35020 75590
rect 35076 75588 35100 75590
rect 35156 75588 35180 75590
rect 35236 75588 35242 75590
rect 34934 75579 35242 75588
rect 65654 75644 65962 75653
rect 65654 75642 65660 75644
rect 65716 75642 65740 75644
rect 65796 75642 65820 75644
rect 65876 75642 65900 75644
rect 65956 75642 65962 75644
rect 65716 75590 65718 75642
rect 65898 75590 65900 75642
rect 65654 75588 65660 75590
rect 65716 75588 65740 75590
rect 65796 75588 65820 75590
rect 65876 75588 65900 75590
rect 65956 75588 65962 75590
rect 65654 75579 65962 75588
rect 1676 75336 1728 75342
rect 1674 75304 1676 75313
rect 1728 75304 1730 75313
rect 1674 75239 1730 75248
rect 1492 75200 1544 75206
rect 1492 75142 1544 75148
rect 76564 75200 76616 75206
rect 76564 75142 76616 75148
rect 78036 75200 78088 75206
rect 78036 75142 78088 75148
rect 1504 75041 1532 75142
rect 19574 75100 19882 75109
rect 19574 75098 19580 75100
rect 19636 75098 19660 75100
rect 19716 75098 19740 75100
rect 19796 75098 19820 75100
rect 19876 75098 19882 75100
rect 19636 75046 19638 75098
rect 19818 75046 19820 75098
rect 19574 75044 19580 75046
rect 19636 75044 19660 75046
rect 19716 75044 19740 75046
rect 19796 75044 19820 75046
rect 19876 75044 19882 75046
rect 1490 75032 1546 75041
rect 19574 75035 19882 75044
rect 50294 75100 50602 75109
rect 50294 75098 50300 75100
rect 50356 75098 50380 75100
rect 50436 75098 50460 75100
rect 50516 75098 50540 75100
rect 50596 75098 50602 75100
rect 50356 75046 50358 75098
rect 50538 75046 50540 75098
rect 50294 75044 50300 75046
rect 50356 75044 50380 75046
rect 50436 75044 50460 75046
rect 50516 75044 50540 75046
rect 50596 75044 50602 75046
rect 50294 75035 50602 75044
rect 1490 74967 1546 74976
rect 1400 74860 1452 74866
rect 1400 74802 1452 74808
rect 1412 74390 1440 74802
rect 2412 74656 2464 74662
rect 2412 74598 2464 74604
rect 2424 74534 2452 74598
rect 4214 74556 4522 74565
rect 4214 74554 4220 74556
rect 4276 74554 4300 74556
rect 4356 74554 4380 74556
rect 4436 74554 4460 74556
rect 4516 74554 4522 74556
rect 2424 74506 2544 74534
rect 1400 74384 1452 74390
rect 1398 74352 1400 74361
rect 1452 74352 1454 74361
rect 1398 74287 1454 74296
rect 1412 74261 1440 74287
rect 1490 73672 1546 73681
rect 1490 73607 1492 73616
rect 1544 73607 1546 73616
rect 1492 73578 1544 73584
rect 1492 73024 1544 73030
rect 1490 72992 1492 73001
rect 2320 73024 2372 73030
rect 1544 72992 1546 73001
rect 2320 72966 2372 72972
rect 1490 72927 1546 72936
rect 1492 72480 1544 72486
rect 1492 72422 1544 72428
rect 1504 72321 1532 72422
rect 1490 72312 1546 72321
rect 1490 72247 1546 72256
rect 1492 71936 1544 71942
rect 1492 71878 1544 71884
rect 2228 71936 2280 71942
rect 2228 71878 2280 71884
rect 1504 71641 1532 71878
rect 1490 71632 1546 71641
rect 1490 71567 1546 71576
rect 1490 70952 1546 70961
rect 1490 70887 1546 70896
rect 1504 70854 1532 70887
rect 1492 70848 1544 70854
rect 1492 70790 1544 70796
rect 2240 70582 2268 71878
rect 2332 71398 2360 72966
rect 2412 72480 2464 72486
rect 2412 72422 2464 72428
rect 2320 71392 2372 71398
rect 2320 71334 2372 71340
rect 2424 70922 2452 72422
rect 2412 70916 2464 70922
rect 2412 70858 2464 70864
rect 2320 70848 2372 70854
rect 2320 70790 2372 70796
rect 2228 70576 2280 70582
rect 2228 70518 2280 70524
rect 2228 70440 2280 70446
rect 2228 70382 2280 70388
rect 1492 70304 1544 70310
rect 1490 70272 1492 70281
rect 1544 70272 1546 70281
rect 1490 70207 1546 70216
rect 1400 69896 1452 69902
rect 1400 69838 1452 69844
rect 1412 69601 1440 69838
rect 1768 69760 1820 69766
rect 1768 69702 1820 69708
rect 1398 69592 1454 69601
rect 1398 69527 1454 69536
rect 1400 69420 1452 69426
rect 1400 69362 1452 69368
rect 1412 68921 1440 69362
rect 1676 69216 1728 69222
rect 1676 69158 1728 69164
rect 1398 68912 1454 68921
rect 1398 68847 1454 68856
rect 1400 68672 1452 68678
rect 1400 68614 1452 68620
rect 1412 68338 1440 68614
rect 1400 68332 1452 68338
rect 1400 68274 1452 68280
rect 1412 68241 1440 68274
rect 1398 68232 1454 68241
rect 1398 68167 1454 68176
rect 1400 67720 1452 67726
rect 1400 67662 1452 67668
rect 1412 67561 1440 67662
rect 1398 67552 1454 67561
rect 1398 67487 1454 67496
rect 1400 67244 1452 67250
rect 1400 67186 1452 67192
rect 1412 66881 1440 67186
rect 1584 67040 1636 67046
rect 1584 66982 1636 66988
rect 1398 66872 1454 66881
rect 1596 66842 1624 66982
rect 1398 66807 1454 66816
rect 1584 66836 1636 66842
rect 1584 66778 1636 66784
rect 1400 66632 1452 66638
rect 1400 66574 1452 66580
rect 1412 66201 1440 66574
rect 1584 66496 1636 66502
rect 1584 66438 1636 66444
rect 1398 66192 1454 66201
rect 1398 66127 1454 66136
rect 1400 65952 1452 65958
rect 1400 65894 1452 65900
rect 1412 65550 1440 65894
rect 1400 65544 1452 65550
rect 1398 65512 1400 65521
rect 1452 65512 1454 65521
rect 1398 65447 1454 65456
rect 1400 65068 1452 65074
rect 1400 65010 1452 65016
rect 1412 64841 1440 65010
rect 1398 64832 1454 64841
rect 1398 64767 1454 64776
rect 1400 64456 1452 64462
rect 1400 64398 1452 64404
rect 1412 64161 1440 64398
rect 1492 64320 1544 64326
rect 1492 64262 1544 64268
rect 1398 64152 1454 64161
rect 1398 64087 1454 64096
rect 1400 63980 1452 63986
rect 1400 63922 1452 63928
rect 1412 63481 1440 63922
rect 1398 63472 1454 63481
rect 1398 63407 1454 63416
rect 1400 63232 1452 63238
rect 1400 63174 1452 63180
rect 1412 62898 1440 63174
rect 1400 62892 1452 62898
rect 1400 62834 1452 62840
rect 1412 62801 1440 62834
rect 1398 62792 1454 62801
rect 1398 62727 1454 62736
rect 1400 62280 1452 62286
rect 1400 62222 1452 62228
rect 1412 62121 1440 62222
rect 1398 62112 1454 62121
rect 1398 62047 1454 62056
rect 1400 61804 1452 61810
rect 1400 61746 1452 61752
rect 1412 61441 1440 61746
rect 1398 61432 1454 61441
rect 1398 61367 1454 61376
rect 1400 61192 1452 61198
rect 1400 61134 1452 61140
rect 1412 60761 1440 61134
rect 1398 60752 1454 60761
rect 1398 60687 1454 60696
rect 1400 60512 1452 60518
rect 1400 60454 1452 60460
rect 1412 60110 1440 60454
rect 1400 60104 1452 60110
rect 1398 60072 1400 60081
rect 1452 60072 1454 60081
rect 1398 60007 1454 60016
rect 1400 59628 1452 59634
rect 1400 59570 1452 59576
rect 1412 59401 1440 59570
rect 1398 59392 1454 59401
rect 1398 59327 1454 59336
rect 1400 59016 1452 59022
rect 1400 58958 1452 58964
rect 1412 58721 1440 58958
rect 1398 58712 1454 58721
rect 1398 58647 1454 58656
rect 1400 58540 1452 58546
rect 1400 58482 1452 58488
rect 1412 58041 1440 58482
rect 1398 58032 1454 58041
rect 1398 57967 1454 57976
rect 1400 57792 1452 57798
rect 1400 57734 1452 57740
rect 1412 57458 1440 57734
rect 1504 57594 1532 64262
rect 1596 61402 1624 66438
rect 1584 61396 1636 61402
rect 1584 61338 1636 61344
rect 1688 60217 1716 69158
rect 1780 62218 1808 69702
rect 2240 68678 2268 70382
rect 2332 69834 2360 70790
rect 2320 69828 2372 69834
rect 2320 69770 2372 69776
rect 2228 68672 2280 68678
rect 2228 68614 2280 68620
rect 1860 67856 1912 67862
rect 1860 67798 1912 67804
rect 1768 62212 1820 62218
rect 1768 62154 1820 62160
rect 1674 60208 1730 60217
rect 1674 60143 1730 60152
rect 1872 59673 1900 67798
rect 2320 65204 2372 65210
rect 2320 65146 2372 65152
rect 2228 63776 2280 63782
rect 2228 63718 2280 63724
rect 2136 62688 2188 62694
rect 2136 62630 2188 62636
rect 1952 62144 2004 62150
rect 1952 62086 2004 62092
rect 1858 59664 1914 59673
rect 1858 59599 1914 59608
rect 1584 58880 1636 58886
rect 1584 58822 1636 58828
rect 1596 58614 1624 58822
rect 1584 58608 1636 58614
rect 1584 58550 1636 58556
rect 1492 57588 1544 57594
rect 1492 57530 1544 57536
rect 1400 57452 1452 57458
rect 1400 57394 1452 57400
rect 1412 57361 1440 57394
rect 1398 57352 1454 57361
rect 1398 57287 1454 57296
rect 1584 57248 1636 57254
rect 1584 57190 1636 57196
rect 1400 56840 1452 56846
rect 1400 56782 1452 56788
rect 1412 56681 1440 56782
rect 1398 56672 1454 56681
rect 1398 56607 1454 56616
rect 1596 56506 1624 57190
rect 1964 56914 1992 62086
rect 2044 61056 2096 61062
rect 2044 60998 2096 61004
rect 1952 56908 2004 56914
rect 1952 56850 2004 56856
rect 2056 56778 2084 60998
rect 2148 58410 2176 62630
rect 2240 59498 2268 63718
rect 2332 59566 2360 65146
rect 2412 61600 2464 61606
rect 2412 61542 2464 61548
rect 2320 59560 2372 59566
rect 2320 59502 2372 59508
rect 2228 59492 2280 59498
rect 2228 59434 2280 59440
rect 2424 59022 2452 61542
rect 2412 59016 2464 59022
rect 2412 58958 2464 58964
rect 2136 58404 2188 58410
rect 2136 58346 2188 58352
rect 2044 56772 2096 56778
rect 2044 56714 2096 56720
rect 1584 56500 1636 56506
rect 1584 56442 1636 56448
rect 1400 56364 1452 56370
rect 1400 56306 1452 56312
rect 1412 56001 1440 56306
rect 1398 55992 1454 56001
rect 1398 55927 1454 55936
rect 1492 55684 1544 55690
rect 1492 55626 1544 55632
rect 1504 55321 1532 55626
rect 1490 55312 1546 55321
rect 1490 55247 1546 55256
rect 1492 55072 1544 55078
rect 1492 55014 1544 55020
rect 1504 54670 1532 55014
rect 1492 54664 1544 54670
rect 1490 54632 1492 54641
rect 1544 54632 1546 54641
rect 1490 54567 1546 54576
rect 1492 54188 1544 54194
rect 1492 54130 1544 54136
rect 1504 53961 1532 54130
rect 1676 54052 1728 54058
rect 1676 53994 1728 54000
rect 1490 53952 1546 53961
rect 1490 53887 1546 53896
rect 1492 53508 1544 53514
rect 1492 53450 1544 53456
rect 1504 53281 1532 53450
rect 1490 53272 1546 53281
rect 1490 53207 1546 53216
rect 1688 53174 1716 53994
rect 1676 53168 1728 53174
rect 1676 53110 1728 53116
rect 1492 53100 1544 53106
rect 1492 53042 1544 53048
rect 1504 52601 1532 53042
rect 1490 52592 1546 52601
rect 1490 52527 1546 52536
rect 1492 52352 1544 52358
rect 1492 52294 1544 52300
rect 1504 52018 1532 52294
rect 1492 52012 1544 52018
rect 1492 51954 1544 51960
rect 1504 51921 1532 51954
rect 1490 51912 1546 51921
rect 1490 51847 1546 51856
rect 1584 51808 1636 51814
rect 1584 51750 1636 51756
rect 1596 51610 1624 51750
rect 1584 51604 1636 51610
rect 1584 51546 1636 51552
rect 1492 51332 1544 51338
rect 1492 51274 1544 51280
rect 1504 51241 1532 51274
rect 1490 51232 1546 51241
rect 1490 51167 1546 51176
rect 1492 50924 1544 50930
rect 1492 50866 1544 50872
rect 1504 50561 1532 50866
rect 1490 50552 1546 50561
rect 1490 50487 1546 50496
rect 2516 50386 2544 74506
rect 4276 74502 4278 74554
rect 4458 74502 4460 74554
rect 4214 74500 4220 74502
rect 4276 74500 4300 74502
rect 4356 74500 4380 74502
rect 4436 74500 4460 74502
rect 4516 74500 4522 74502
rect 4214 74491 4522 74500
rect 34934 74556 35242 74565
rect 34934 74554 34940 74556
rect 34996 74554 35020 74556
rect 35076 74554 35100 74556
rect 35156 74554 35180 74556
rect 35236 74554 35242 74556
rect 34996 74502 34998 74554
rect 35178 74502 35180 74554
rect 34934 74500 34940 74502
rect 34996 74500 35020 74502
rect 35076 74500 35100 74502
rect 35156 74500 35180 74502
rect 35236 74500 35242 74502
rect 34934 74491 35242 74500
rect 65654 74556 65962 74565
rect 65654 74554 65660 74556
rect 65716 74554 65740 74556
rect 65796 74554 65820 74556
rect 65876 74554 65900 74556
rect 65956 74554 65962 74556
rect 65716 74502 65718 74554
rect 65898 74502 65900 74554
rect 65654 74500 65660 74502
rect 65716 74500 65740 74502
rect 65796 74500 65820 74502
rect 65876 74500 65900 74502
rect 65956 74500 65962 74502
rect 65654 74491 65962 74500
rect 19574 74012 19882 74021
rect 19574 74010 19580 74012
rect 19636 74010 19660 74012
rect 19716 74010 19740 74012
rect 19796 74010 19820 74012
rect 19876 74010 19882 74012
rect 19636 73958 19638 74010
rect 19818 73958 19820 74010
rect 19574 73956 19580 73958
rect 19636 73956 19660 73958
rect 19716 73956 19740 73958
rect 19796 73956 19820 73958
rect 19876 73956 19882 73958
rect 19574 73947 19882 73956
rect 50294 74012 50602 74021
rect 50294 74010 50300 74012
rect 50356 74010 50380 74012
rect 50436 74010 50460 74012
rect 50516 74010 50540 74012
rect 50596 74010 50602 74012
rect 50356 73958 50358 74010
rect 50538 73958 50540 74010
rect 50294 73956 50300 73958
rect 50356 73956 50380 73958
rect 50436 73956 50460 73958
rect 50516 73956 50540 73958
rect 50596 73956 50602 73958
rect 50294 73947 50602 73956
rect 2688 73568 2740 73574
rect 2688 73510 2740 73516
rect 2700 61606 2728 73510
rect 4214 73468 4522 73477
rect 4214 73466 4220 73468
rect 4276 73466 4300 73468
rect 4356 73466 4380 73468
rect 4436 73466 4460 73468
rect 4516 73466 4522 73468
rect 4276 73414 4278 73466
rect 4458 73414 4460 73466
rect 4214 73412 4220 73414
rect 4276 73412 4300 73414
rect 4356 73412 4380 73414
rect 4436 73412 4460 73414
rect 4516 73412 4522 73414
rect 4214 73403 4522 73412
rect 34934 73468 35242 73477
rect 34934 73466 34940 73468
rect 34996 73466 35020 73468
rect 35076 73466 35100 73468
rect 35156 73466 35180 73468
rect 35236 73466 35242 73468
rect 34996 73414 34998 73466
rect 35178 73414 35180 73466
rect 34934 73412 34940 73414
rect 34996 73412 35020 73414
rect 35076 73412 35100 73414
rect 35156 73412 35180 73414
rect 35236 73412 35242 73414
rect 34934 73403 35242 73412
rect 65654 73468 65962 73477
rect 65654 73466 65660 73468
rect 65716 73466 65740 73468
rect 65796 73466 65820 73468
rect 65876 73466 65900 73468
rect 65956 73466 65962 73468
rect 65716 73414 65718 73466
rect 65898 73414 65900 73466
rect 65654 73412 65660 73414
rect 65716 73412 65740 73414
rect 65796 73412 65820 73414
rect 65876 73412 65900 73414
rect 65956 73412 65962 73414
rect 65654 73403 65962 73412
rect 76196 73160 76248 73166
rect 76196 73102 76248 73108
rect 19574 72924 19882 72933
rect 19574 72922 19580 72924
rect 19636 72922 19660 72924
rect 19716 72922 19740 72924
rect 19796 72922 19820 72924
rect 19876 72922 19882 72924
rect 19636 72870 19638 72922
rect 19818 72870 19820 72922
rect 19574 72868 19580 72870
rect 19636 72868 19660 72870
rect 19716 72868 19740 72870
rect 19796 72868 19820 72870
rect 19876 72868 19882 72870
rect 19574 72859 19882 72868
rect 50294 72924 50602 72933
rect 50294 72922 50300 72924
rect 50356 72922 50380 72924
rect 50436 72922 50460 72924
rect 50516 72922 50540 72924
rect 50596 72922 50602 72924
rect 50356 72870 50358 72922
rect 50538 72870 50540 72922
rect 50294 72868 50300 72870
rect 50356 72868 50380 72870
rect 50436 72868 50460 72870
rect 50516 72868 50540 72870
rect 50596 72868 50602 72870
rect 50294 72859 50602 72868
rect 76104 72684 76156 72690
rect 76104 72626 76156 72632
rect 4214 72380 4522 72389
rect 4214 72378 4220 72380
rect 4276 72378 4300 72380
rect 4356 72378 4380 72380
rect 4436 72378 4460 72380
rect 4516 72378 4522 72380
rect 4276 72326 4278 72378
rect 4458 72326 4460 72378
rect 4214 72324 4220 72326
rect 4276 72324 4300 72326
rect 4356 72324 4380 72326
rect 4436 72324 4460 72326
rect 4516 72324 4522 72326
rect 4214 72315 4522 72324
rect 34934 72380 35242 72389
rect 34934 72378 34940 72380
rect 34996 72378 35020 72380
rect 35076 72378 35100 72380
rect 35156 72378 35180 72380
rect 35236 72378 35242 72380
rect 34996 72326 34998 72378
rect 35178 72326 35180 72378
rect 34934 72324 34940 72326
rect 34996 72324 35020 72326
rect 35076 72324 35100 72326
rect 35156 72324 35180 72326
rect 35236 72324 35242 72326
rect 34934 72315 35242 72324
rect 65654 72380 65962 72389
rect 65654 72378 65660 72380
rect 65716 72378 65740 72380
rect 65796 72378 65820 72380
rect 65876 72378 65900 72380
rect 65956 72378 65962 72380
rect 65716 72326 65718 72378
rect 65898 72326 65900 72378
rect 65654 72324 65660 72326
rect 65716 72324 65740 72326
rect 65796 72324 65820 72326
rect 65876 72324 65900 72326
rect 65956 72324 65962 72326
rect 65654 72315 65962 72324
rect 75920 72072 75972 72078
rect 75920 72014 75972 72020
rect 19574 71836 19882 71845
rect 19574 71834 19580 71836
rect 19636 71834 19660 71836
rect 19716 71834 19740 71836
rect 19796 71834 19820 71836
rect 19876 71834 19882 71836
rect 19636 71782 19638 71834
rect 19818 71782 19820 71834
rect 19574 71780 19580 71782
rect 19636 71780 19660 71782
rect 19716 71780 19740 71782
rect 19796 71780 19820 71782
rect 19876 71780 19882 71782
rect 19574 71771 19882 71780
rect 50294 71836 50602 71845
rect 50294 71834 50300 71836
rect 50356 71834 50380 71836
rect 50436 71834 50460 71836
rect 50516 71834 50540 71836
rect 50596 71834 50602 71836
rect 50356 71782 50358 71834
rect 50538 71782 50540 71834
rect 50294 71780 50300 71782
rect 50356 71780 50380 71782
rect 50436 71780 50460 71782
rect 50516 71780 50540 71782
rect 50596 71780 50602 71782
rect 50294 71771 50602 71780
rect 4214 71292 4522 71301
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71227 4522 71236
rect 34934 71292 35242 71301
rect 34934 71290 34940 71292
rect 34996 71290 35020 71292
rect 35076 71290 35100 71292
rect 35156 71290 35180 71292
rect 35236 71290 35242 71292
rect 34996 71238 34998 71290
rect 35178 71238 35180 71290
rect 34934 71236 34940 71238
rect 34996 71236 35020 71238
rect 35076 71236 35100 71238
rect 35156 71236 35180 71238
rect 35236 71236 35242 71238
rect 34934 71227 35242 71236
rect 65654 71292 65962 71301
rect 65654 71290 65660 71292
rect 65716 71290 65740 71292
rect 65796 71290 65820 71292
rect 65876 71290 65900 71292
rect 65956 71290 65962 71292
rect 65716 71238 65718 71290
rect 65898 71238 65900 71290
rect 65654 71236 65660 71238
rect 65716 71236 65740 71238
rect 65796 71236 65820 71238
rect 65876 71236 65900 71238
rect 65956 71236 65962 71238
rect 65654 71227 65962 71236
rect 75828 70916 75880 70922
rect 75828 70858 75880 70864
rect 19574 70748 19882 70757
rect 19574 70746 19580 70748
rect 19636 70746 19660 70748
rect 19716 70746 19740 70748
rect 19796 70746 19820 70748
rect 19876 70746 19882 70748
rect 19636 70694 19638 70746
rect 19818 70694 19820 70746
rect 19574 70692 19580 70694
rect 19636 70692 19660 70694
rect 19716 70692 19740 70694
rect 19796 70692 19820 70694
rect 19876 70692 19882 70694
rect 19574 70683 19882 70692
rect 50294 70748 50602 70757
rect 50294 70746 50300 70748
rect 50356 70746 50380 70748
rect 50436 70746 50460 70748
rect 50516 70746 50540 70748
rect 50596 70746 50602 70748
rect 50356 70694 50358 70746
rect 50538 70694 50540 70746
rect 50294 70692 50300 70694
rect 50356 70692 50380 70694
rect 50436 70692 50460 70694
rect 50516 70692 50540 70694
rect 50596 70692 50602 70694
rect 50294 70683 50602 70692
rect 75000 70508 75052 70514
rect 75000 70450 75052 70456
rect 73344 70440 73396 70446
rect 73344 70382 73396 70388
rect 4214 70204 4522 70213
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 4214 70139 4522 70148
rect 34934 70204 35242 70213
rect 34934 70202 34940 70204
rect 34996 70202 35020 70204
rect 35076 70202 35100 70204
rect 35156 70202 35180 70204
rect 35236 70202 35242 70204
rect 34996 70150 34998 70202
rect 35178 70150 35180 70202
rect 34934 70148 34940 70150
rect 34996 70148 35020 70150
rect 35076 70148 35100 70150
rect 35156 70148 35180 70150
rect 35236 70148 35242 70150
rect 34934 70139 35242 70148
rect 65654 70204 65962 70213
rect 65654 70202 65660 70204
rect 65716 70202 65740 70204
rect 65796 70202 65820 70204
rect 65876 70202 65900 70204
rect 65956 70202 65962 70204
rect 65716 70150 65718 70202
rect 65898 70150 65900 70202
rect 65654 70148 65660 70150
rect 65716 70148 65740 70150
rect 65796 70148 65820 70150
rect 65876 70148 65900 70150
rect 65956 70148 65962 70150
rect 65654 70139 65962 70148
rect 19574 69660 19882 69669
rect 19574 69658 19580 69660
rect 19636 69658 19660 69660
rect 19716 69658 19740 69660
rect 19796 69658 19820 69660
rect 19876 69658 19882 69660
rect 19636 69606 19638 69658
rect 19818 69606 19820 69658
rect 19574 69604 19580 69606
rect 19636 69604 19660 69606
rect 19716 69604 19740 69606
rect 19796 69604 19820 69606
rect 19876 69604 19882 69606
rect 19574 69595 19882 69604
rect 50294 69660 50602 69669
rect 50294 69658 50300 69660
rect 50356 69658 50380 69660
rect 50436 69658 50460 69660
rect 50516 69658 50540 69660
rect 50596 69658 50602 69660
rect 50356 69606 50358 69658
rect 50538 69606 50540 69658
rect 50294 69604 50300 69606
rect 50356 69604 50380 69606
rect 50436 69604 50460 69606
rect 50516 69604 50540 69606
rect 50596 69604 50602 69606
rect 50294 69595 50602 69604
rect 65984 69556 66036 69562
rect 65984 69498 66036 69504
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 34934 69116 35242 69125
rect 34934 69114 34940 69116
rect 34996 69114 35020 69116
rect 35076 69114 35100 69116
rect 35156 69114 35180 69116
rect 35236 69114 35242 69116
rect 34996 69062 34998 69114
rect 35178 69062 35180 69114
rect 34934 69060 34940 69062
rect 34996 69060 35020 69062
rect 35076 69060 35100 69062
rect 35156 69060 35180 69062
rect 35236 69060 35242 69062
rect 34934 69051 35242 69060
rect 65654 69116 65962 69125
rect 65654 69114 65660 69116
rect 65716 69114 65740 69116
rect 65796 69114 65820 69116
rect 65876 69114 65900 69116
rect 65956 69114 65962 69116
rect 65716 69062 65718 69114
rect 65898 69062 65900 69114
rect 65654 69060 65660 69062
rect 65716 69060 65740 69062
rect 65796 69060 65820 69062
rect 65876 69060 65900 69062
rect 65956 69060 65962 69062
rect 65654 69051 65962 69060
rect 19574 68572 19882 68581
rect 19574 68570 19580 68572
rect 19636 68570 19660 68572
rect 19716 68570 19740 68572
rect 19796 68570 19820 68572
rect 19876 68570 19882 68572
rect 19636 68518 19638 68570
rect 19818 68518 19820 68570
rect 19574 68516 19580 68518
rect 19636 68516 19660 68518
rect 19716 68516 19740 68518
rect 19796 68516 19820 68518
rect 19876 68516 19882 68518
rect 19574 68507 19882 68516
rect 50294 68572 50602 68581
rect 50294 68570 50300 68572
rect 50356 68570 50380 68572
rect 50436 68570 50460 68572
rect 50516 68570 50540 68572
rect 50596 68570 50602 68572
rect 50356 68518 50358 68570
rect 50538 68518 50540 68570
rect 50294 68516 50300 68518
rect 50356 68516 50380 68518
rect 50436 68516 50460 68518
rect 50516 68516 50540 68518
rect 50596 68516 50602 68518
rect 50294 68507 50602 68516
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 34934 68028 35242 68037
rect 34934 68026 34940 68028
rect 34996 68026 35020 68028
rect 35076 68026 35100 68028
rect 35156 68026 35180 68028
rect 35236 68026 35242 68028
rect 34996 67974 34998 68026
rect 35178 67974 35180 68026
rect 34934 67972 34940 67974
rect 34996 67972 35020 67974
rect 35076 67972 35100 67974
rect 35156 67972 35180 67974
rect 35236 67972 35242 67974
rect 34934 67963 35242 67972
rect 65654 68028 65962 68037
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67963 65962 67972
rect 19574 67484 19882 67493
rect 19574 67482 19580 67484
rect 19636 67482 19660 67484
rect 19716 67482 19740 67484
rect 19796 67482 19820 67484
rect 19876 67482 19882 67484
rect 19636 67430 19638 67482
rect 19818 67430 19820 67482
rect 19574 67428 19580 67430
rect 19636 67428 19660 67430
rect 19716 67428 19740 67430
rect 19796 67428 19820 67430
rect 19876 67428 19882 67430
rect 19574 67419 19882 67428
rect 50294 67484 50602 67493
rect 50294 67482 50300 67484
rect 50356 67482 50380 67484
rect 50436 67482 50460 67484
rect 50516 67482 50540 67484
rect 50596 67482 50602 67484
rect 50356 67430 50358 67482
rect 50538 67430 50540 67482
rect 50294 67428 50300 67430
rect 50356 67428 50380 67430
rect 50436 67428 50460 67430
rect 50516 67428 50540 67430
rect 50596 67428 50602 67430
rect 50294 67419 50602 67428
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 34934 66940 35242 66949
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66875 35242 66884
rect 65654 66940 65962 66949
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66875 65962 66884
rect 63132 66836 63184 66842
rect 63132 66778 63184 66784
rect 19574 66396 19882 66405
rect 19574 66394 19580 66396
rect 19636 66394 19660 66396
rect 19716 66394 19740 66396
rect 19796 66394 19820 66396
rect 19876 66394 19882 66396
rect 19636 66342 19638 66394
rect 19818 66342 19820 66394
rect 19574 66340 19580 66342
rect 19636 66340 19660 66342
rect 19716 66340 19740 66342
rect 19796 66340 19820 66342
rect 19876 66340 19882 66342
rect 19574 66331 19882 66340
rect 50294 66396 50602 66405
rect 50294 66394 50300 66396
rect 50356 66394 50380 66396
rect 50436 66394 50460 66396
rect 50516 66394 50540 66396
rect 50596 66394 50602 66396
rect 50356 66342 50358 66394
rect 50538 66342 50540 66394
rect 50294 66340 50300 66342
rect 50356 66340 50380 66342
rect 50436 66340 50460 66342
rect 50516 66340 50540 66342
rect 50596 66340 50602 66342
rect 50294 66331 50602 66340
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 34934 65852 35242 65861
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65787 35242 65796
rect 19574 65308 19882 65317
rect 19574 65306 19580 65308
rect 19636 65306 19660 65308
rect 19716 65306 19740 65308
rect 19796 65306 19820 65308
rect 19876 65306 19882 65308
rect 19636 65254 19638 65306
rect 19818 65254 19820 65306
rect 19574 65252 19580 65254
rect 19636 65252 19660 65254
rect 19716 65252 19740 65254
rect 19796 65252 19820 65254
rect 19876 65252 19882 65254
rect 19574 65243 19882 65252
rect 50294 65308 50602 65317
rect 50294 65306 50300 65308
rect 50356 65306 50380 65308
rect 50436 65306 50460 65308
rect 50516 65306 50540 65308
rect 50596 65306 50602 65308
rect 50356 65254 50358 65306
rect 50538 65254 50540 65306
rect 50294 65252 50300 65254
rect 50356 65252 50380 65254
rect 50436 65252 50460 65254
rect 50516 65252 50540 65254
rect 50596 65252 50602 65254
rect 50294 65243 50602 65252
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 34934 64764 35242 64773
rect 34934 64762 34940 64764
rect 34996 64762 35020 64764
rect 35076 64762 35100 64764
rect 35156 64762 35180 64764
rect 35236 64762 35242 64764
rect 34996 64710 34998 64762
rect 35178 64710 35180 64762
rect 34934 64708 34940 64710
rect 34996 64708 35020 64710
rect 35076 64708 35100 64710
rect 35156 64708 35180 64710
rect 35236 64708 35242 64710
rect 34934 64699 35242 64708
rect 19574 64220 19882 64229
rect 19574 64218 19580 64220
rect 19636 64218 19660 64220
rect 19716 64218 19740 64220
rect 19796 64218 19820 64220
rect 19876 64218 19882 64220
rect 19636 64166 19638 64218
rect 19818 64166 19820 64218
rect 19574 64164 19580 64166
rect 19636 64164 19660 64166
rect 19716 64164 19740 64166
rect 19796 64164 19820 64166
rect 19876 64164 19882 64166
rect 19574 64155 19882 64164
rect 50294 64220 50602 64229
rect 50294 64218 50300 64220
rect 50356 64218 50380 64220
rect 50436 64218 50460 64220
rect 50516 64218 50540 64220
rect 50596 64218 50602 64220
rect 50356 64166 50358 64218
rect 50538 64166 50540 64218
rect 50294 64164 50300 64166
rect 50356 64164 50380 64166
rect 50436 64164 50460 64166
rect 50516 64164 50540 64166
rect 50596 64164 50602 64166
rect 50294 64155 50602 64164
rect 62672 63776 62724 63782
rect 62672 63718 62724 63724
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 34934 63676 35242 63685
rect 34934 63674 34940 63676
rect 34996 63674 35020 63676
rect 35076 63674 35100 63676
rect 35156 63674 35180 63676
rect 35236 63674 35242 63676
rect 34996 63622 34998 63674
rect 35178 63622 35180 63674
rect 34934 63620 34940 63622
rect 34996 63620 35020 63622
rect 35076 63620 35100 63622
rect 35156 63620 35180 63622
rect 35236 63620 35242 63622
rect 34934 63611 35242 63620
rect 19574 63132 19882 63141
rect 19574 63130 19580 63132
rect 19636 63130 19660 63132
rect 19716 63130 19740 63132
rect 19796 63130 19820 63132
rect 19876 63130 19882 63132
rect 19636 63078 19638 63130
rect 19818 63078 19820 63130
rect 19574 63076 19580 63078
rect 19636 63076 19660 63078
rect 19716 63076 19740 63078
rect 19796 63076 19820 63078
rect 19876 63076 19882 63078
rect 19574 63067 19882 63076
rect 50294 63132 50602 63141
rect 50294 63130 50300 63132
rect 50356 63130 50380 63132
rect 50436 63130 50460 63132
rect 50516 63130 50540 63132
rect 50596 63130 50602 63132
rect 50356 63078 50358 63130
rect 50538 63078 50540 63130
rect 50294 63076 50300 63078
rect 50356 63076 50380 63078
rect 50436 63076 50460 63078
rect 50516 63076 50540 63078
rect 50596 63076 50602 63078
rect 50294 63067 50602 63076
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 34934 62588 35242 62597
rect 34934 62586 34940 62588
rect 34996 62586 35020 62588
rect 35076 62586 35100 62588
rect 35156 62586 35180 62588
rect 35236 62586 35242 62588
rect 34996 62534 34998 62586
rect 35178 62534 35180 62586
rect 34934 62532 34940 62534
rect 34996 62532 35020 62534
rect 35076 62532 35100 62534
rect 35156 62532 35180 62534
rect 35236 62532 35242 62534
rect 34934 62523 35242 62532
rect 19574 62044 19882 62053
rect 19574 62042 19580 62044
rect 19636 62042 19660 62044
rect 19716 62042 19740 62044
rect 19796 62042 19820 62044
rect 19876 62042 19882 62044
rect 19636 61990 19638 62042
rect 19818 61990 19820 62042
rect 19574 61988 19580 61990
rect 19636 61988 19660 61990
rect 19716 61988 19740 61990
rect 19796 61988 19820 61990
rect 19876 61988 19882 61990
rect 19574 61979 19882 61988
rect 50294 62044 50602 62053
rect 50294 62042 50300 62044
rect 50356 62042 50380 62044
rect 50436 62042 50460 62044
rect 50516 62042 50540 62044
rect 50596 62042 50602 62044
rect 50356 61990 50358 62042
rect 50538 61990 50540 62042
rect 50294 61988 50300 61990
rect 50356 61988 50380 61990
rect 50436 61988 50460 61990
rect 50516 61988 50540 61990
rect 50596 61988 50602 61990
rect 50294 61979 50602 61988
rect 61660 61668 61712 61674
rect 61660 61610 61712 61616
rect 2688 61600 2740 61606
rect 2688 61542 2740 61548
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 34934 61500 35242 61509
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61435 35242 61444
rect 61672 61402 61700 61610
rect 61660 61396 61712 61402
rect 61660 61338 61712 61344
rect 19574 60956 19882 60965
rect 19574 60954 19580 60956
rect 19636 60954 19660 60956
rect 19716 60954 19740 60956
rect 19796 60954 19820 60956
rect 19876 60954 19882 60956
rect 19636 60902 19638 60954
rect 19818 60902 19820 60954
rect 19574 60900 19580 60902
rect 19636 60900 19660 60902
rect 19716 60900 19740 60902
rect 19796 60900 19820 60902
rect 19876 60900 19882 60902
rect 19574 60891 19882 60900
rect 50294 60956 50602 60965
rect 50294 60954 50300 60956
rect 50356 60954 50380 60956
rect 50436 60954 50460 60956
rect 50516 60954 50540 60956
rect 50596 60954 50602 60956
rect 50356 60902 50358 60954
rect 50538 60902 50540 60954
rect 50294 60900 50300 60902
rect 50356 60900 50380 60902
rect 50436 60900 50460 60902
rect 50516 60900 50540 60902
rect 50596 60900 50602 60902
rect 50294 60891 50602 60900
rect 60004 60784 60056 60790
rect 60004 60726 60056 60732
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 34934 60412 35242 60421
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60347 35242 60356
rect 59544 60240 59596 60246
rect 59544 60182 59596 60188
rect 2596 59968 2648 59974
rect 2596 59910 2648 59916
rect 2608 57866 2636 59910
rect 19574 59868 19882 59877
rect 19574 59866 19580 59868
rect 19636 59866 19660 59868
rect 19716 59866 19740 59868
rect 19796 59866 19820 59868
rect 19876 59866 19882 59868
rect 19636 59814 19638 59866
rect 19818 59814 19820 59866
rect 19574 59812 19580 59814
rect 19636 59812 19660 59814
rect 19716 59812 19740 59814
rect 19796 59812 19820 59814
rect 19876 59812 19882 59814
rect 19574 59803 19882 59812
rect 50294 59868 50602 59877
rect 50294 59866 50300 59868
rect 50356 59866 50380 59868
rect 50436 59866 50460 59868
rect 50516 59866 50540 59868
rect 50596 59866 50602 59868
rect 50356 59814 50358 59866
rect 50538 59814 50540 59866
rect 50294 59812 50300 59814
rect 50356 59812 50380 59814
rect 50436 59812 50460 59814
rect 50516 59812 50540 59814
rect 50596 59812 50602 59814
rect 50294 59803 50602 59812
rect 2688 59424 2740 59430
rect 2688 59366 2740 59372
rect 2700 58682 2728 59366
rect 4214 59324 4522 59333
rect 4214 59322 4220 59324
rect 4276 59322 4300 59324
rect 4356 59322 4380 59324
rect 4436 59322 4460 59324
rect 4516 59322 4522 59324
rect 4276 59270 4278 59322
rect 4458 59270 4460 59322
rect 4214 59268 4220 59270
rect 4276 59268 4300 59270
rect 4356 59268 4380 59270
rect 4436 59268 4460 59270
rect 4516 59268 4522 59270
rect 4214 59259 4522 59268
rect 34934 59324 35242 59333
rect 34934 59322 34940 59324
rect 34996 59322 35020 59324
rect 35076 59322 35100 59324
rect 35156 59322 35180 59324
rect 35236 59322 35242 59324
rect 34996 59270 34998 59322
rect 35178 59270 35180 59322
rect 34934 59268 34940 59270
rect 34996 59268 35020 59270
rect 35076 59268 35100 59270
rect 35156 59268 35180 59270
rect 35236 59268 35242 59270
rect 34934 59259 35242 59268
rect 19574 58780 19882 58789
rect 19574 58778 19580 58780
rect 19636 58778 19660 58780
rect 19716 58778 19740 58780
rect 19796 58778 19820 58780
rect 19876 58778 19882 58780
rect 19636 58726 19638 58778
rect 19818 58726 19820 58778
rect 19574 58724 19580 58726
rect 19636 58724 19660 58726
rect 19716 58724 19740 58726
rect 19796 58724 19820 58726
rect 19876 58724 19882 58726
rect 19574 58715 19882 58724
rect 50294 58780 50602 58789
rect 50294 58778 50300 58780
rect 50356 58778 50380 58780
rect 50436 58778 50460 58780
rect 50516 58778 50540 58780
rect 50596 58778 50602 58780
rect 50356 58726 50358 58778
rect 50538 58726 50540 58778
rect 50294 58724 50300 58726
rect 50356 58724 50380 58726
rect 50436 58724 50460 58726
rect 50516 58724 50540 58726
rect 50596 58724 50602 58726
rect 50294 58715 50602 58724
rect 59556 58682 59584 60182
rect 59820 58880 59872 58886
rect 59820 58822 59872 58828
rect 2688 58676 2740 58682
rect 2688 58618 2740 58624
rect 59544 58676 59596 58682
rect 59544 58618 59596 58624
rect 2688 58336 2740 58342
rect 2688 58278 2740 58284
rect 2596 57860 2648 57866
rect 2596 57802 2648 57808
rect 2700 57254 2728 58278
rect 4214 58236 4522 58245
rect 4214 58234 4220 58236
rect 4276 58234 4300 58236
rect 4356 58234 4380 58236
rect 4436 58234 4460 58236
rect 4516 58234 4522 58236
rect 4276 58182 4278 58234
rect 4458 58182 4460 58234
rect 4214 58180 4220 58182
rect 4276 58180 4300 58182
rect 4356 58180 4380 58182
rect 4436 58180 4460 58182
rect 4516 58180 4522 58182
rect 4214 58171 4522 58180
rect 34934 58236 35242 58245
rect 34934 58234 34940 58236
rect 34996 58234 35020 58236
rect 35076 58234 35100 58236
rect 35156 58234 35180 58236
rect 35236 58234 35242 58236
rect 34996 58182 34998 58234
rect 35178 58182 35180 58234
rect 34934 58180 34940 58182
rect 34996 58180 35020 58182
rect 35076 58180 35100 58182
rect 35156 58180 35180 58182
rect 35236 58180 35242 58182
rect 34934 58171 35242 58180
rect 59556 57934 59584 58618
rect 59832 58546 59860 58822
rect 59820 58540 59872 58546
rect 59820 58482 59872 58488
rect 59544 57928 59596 57934
rect 59544 57870 59596 57876
rect 59728 57928 59780 57934
rect 59728 57870 59780 57876
rect 59544 57792 59596 57798
rect 59544 57734 59596 57740
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 59556 57458 59584 57734
rect 59636 57520 59688 57526
rect 59636 57462 59688 57468
rect 59544 57452 59596 57458
rect 59464 57412 59544 57440
rect 2688 57248 2740 57254
rect 2688 57190 2740 57196
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 59084 56908 59136 56914
rect 59084 56850 59136 56856
rect 2688 56704 2740 56710
rect 2688 56646 2740 56652
rect 2700 55758 2728 56646
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 57704 56500 57756 56506
rect 57704 56442 57756 56448
rect 55956 56228 56008 56234
rect 55956 56170 56008 56176
rect 56784 56228 56836 56234
rect 56784 56170 56836 56176
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 55968 55962 55996 56170
rect 55956 55956 56008 55962
rect 55956 55898 56008 55904
rect 56796 55758 56824 56170
rect 57152 56160 57204 56166
rect 57152 56102 57204 56108
rect 57164 55962 57192 56102
rect 57152 55956 57204 55962
rect 57152 55898 57204 55904
rect 57060 55888 57112 55894
rect 57060 55830 57112 55836
rect 2688 55752 2740 55758
rect 2688 55694 2740 55700
rect 56784 55752 56836 55758
rect 56784 55694 56836 55700
rect 56876 55752 56928 55758
rect 56876 55694 56928 55700
rect 56888 55622 56916 55694
rect 55680 55616 55732 55622
rect 55680 55558 55732 55564
rect 56600 55616 56652 55622
rect 56876 55616 56928 55622
rect 56600 55558 56652 55564
rect 56704 55564 56876 55570
rect 56704 55558 56928 55564
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 55692 55418 55720 55558
rect 55680 55412 55732 55418
rect 55680 55354 55732 55360
rect 56612 55146 56640 55558
rect 56704 55542 56916 55558
rect 56704 55282 56732 55542
rect 56888 55493 56916 55542
rect 56692 55276 56744 55282
rect 56692 55218 56744 55224
rect 56600 55140 56652 55146
rect 56600 55082 56652 55088
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 53104 54732 53156 54738
rect 53104 54674 53156 54680
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 2688 53440 2740 53446
rect 2688 53382 2740 53388
rect 2700 51882 2728 53382
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 52828 53100 52880 53106
rect 52828 53042 52880 53048
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 52840 52698 52868 53042
rect 52828 52692 52880 52698
rect 52828 52634 52880 52640
rect 51816 52556 51868 52562
rect 51816 52498 51868 52504
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 51828 52086 51856 52498
rect 52184 52420 52236 52426
rect 52184 52362 52236 52368
rect 51816 52080 51868 52086
rect 51816 52022 51868 52028
rect 52196 52018 52224 52362
rect 51724 52012 51776 52018
rect 51724 51954 51776 51960
rect 52184 52012 52236 52018
rect 52184 51954 52236 51960
rect 2688 51876 2740 51882
rect 2688 51818 2740 51824
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 51736 51474 51764 51954
rect 52092 51808 52144 51814
rect 52092 51750 52144 51756
rect 51724 51468 51776 51474
rect 51724 51410 51776 51416
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50252 50720 50304 50726
rect 50252 50662 50304 50668
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 50264 50522 50292 50662
rect 50252 50516 50304 50522
rect 50252 50458 50304 50464
rect 51816 50448 51868 50454
rect 51816 50390 51868 50396
rect 2504 50380 2556 50386
rect 2504 50322 2556 50328
rect 51172 50312 51224 50318
rect 51172 50254 51224 50260
rect 1492 50244 1544 50250
rect 1492 50186 1544 50192
rect 50988 50244 51040 50250
rect 50988 50186 51040 50192
rect 1504 49881 1532 50186
rect 49792 50176 49844 50182
rect 49792 50118 49844 50124
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 49804 49978 49832 50118
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 51000 49978 51028 50186
rect 49792 49972 49844 49978
rect 49792 49914 49844 49920
rect 50344 49972 50396 49978
rect 50344 49914 50396 49920
rect 50988 49972 51040 49978
rect 50988 49914 51040 49920
rect 1490 49872 1546 49881
rect 1490 49807 1546 49816
rect 1492 49632 1544 49638
rect 1492 49574 1544 49580
rect 1504 49230 1532 49574
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 50356 49230 50384 49914
rect 51184 49842 51212 50254
rect 50712 49836 50764 49842
rect 50712 49778 50764 49784
rect 51172 49836 51224 49842
rect 51172 49778 51224 49784
rect 50620 49360 50672 49366
rect 50620 49302 50672 49308
rect 1492 49224 1544 49230
rect 1490 49192 1492 49201
rect 50344 49224 50396 49230
rect 1544 49192 1546 49201
rect 1490 49127 1546 49136
rect 50172 49172 50344 49178
rect 50172 49166 50396 49172
rect 50172 49150 50384 49166
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 50172 48890 50200 49150
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50160 48884 50212 48890
rect 50160 48826 50212 48832
rect 1492 48748 1544 48754
rect 1492 48690 1544 48696
rect 1504 48521 1532 48690
rect 49976 48544 50028 48550
rect 1490 48512 1546 48521
rect 49976 48486 50028 48492
rect 1490 48447 1546 48456
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 47768 48068 47820 48074
rect 47768 48010 47820 48016
rect 1492 48000 1544 48006
rect 1492 47942 1544 47948
rect 1504 47841 1532 47942
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 1490 47832 1546 47841
rect 19574 47835 19882 47844
rect 47780 47802 47808 48010
rect 48320 48000 48372 48006
rect 48320 47942 48372 47948
rect 1490 47767 1546 47776
rect 47768 47796 47820 47802
rect 47768 47738 47820 47744
rect 48332 47666 48360 47942
rect 47124 47660 47176 47666
rect 47124 47602 47176 47608
rect 48320 47660 48372 47666
rect 48320 47602 48372 47608
rect 49240 47660 49292 47666
rect 49240 47602 49292 47608
rect 1492 47456 1544 47462
rect 1492 47398 1544 47404
rect 1504 47161 1532 47398
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 47136 47258 47164 47602
rect 49252 47462 49280 47602
rect 49240 47456 49292 47462
rect 49240 47398 49292 47404
rect 47124 47252 47176 47258
rect 47124 47194 47176 47200
rect 1490 47152 1546 47161
rect 1490 47087 1546 47096
rect 47676 47048 47728 47054
rect 47676 46990 47728 46996
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 47688 46714 47716 46990
rect 47676 46708 47728 46714
rect 47676 46650 47728 46656
rect 46388 46572 46440 46578
rect 46388 46514 46440 46520
rect 1490 46472 1546 46481
rect 1490 46407 1492 46416
rect 1544 46407 1546 46416
rect 1492 46378 1544 46384
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 46400 46170 46428 46514
rect 46940 46368 46992 46374
rect 46940 46310 46992 46316
rect 46388 46164 46440 46170
rect 46388 46106 46440 46112
rect 46848 46028 46900 46034
rect 46848 45970 46900 45976
rect 1492 45824 1544 45830
rect 1490 45792 1492 45801
rect 2228 45824 2280 45830
rect 1544 45792 1546 45801
rect 2228 45766 2280 45772
rect 1490 45727 1546 45736
rect 2240 45354 2268 45766
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 46860 45558 46888 45970
rect 46952 45966 46980 46310
rect 46940 45960 46992 45966
rect 46940 45902 46992 45908
rect 46848 45552 46900 45558
rect 47688 45554 47716 46650
rect 47768 45960 47820 45966
rect 47768 45902 47820 45908
rect 46848 45494 46900 45500
rect 47596 45526 47716 45554
rect 44916 45484 44968 45490
rect 44916 45426 44968 45432
rect 46664 45484 46716 45490
rect 46664 45426 46716 45432
rect 2228 45348 2280 45354
rect 2228 45290 2280 45296
rect 1492 45280 1544 45286
rect 1492 45222 1544 45228
rect 1504 45121 1532 45222
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 1490 45112 1546 45121
rect 4214 45115 4522 45124
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 44928 45082 44956 45426
rect 1490 45047 1546 45056
rect 44916 45076 44968 45082
rect 44916 45018 44968 45024
rect 44272 44872 44324 44878
rect 44272 44814 44324 44820
rect 1492 44736 1544 44742
rect 1492 44678 1544 44684
rect 1504 44441 1532 44678
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 44284 44538 44312 44814
rect 45928 44804 45980 44810
rect 45928 44746 45980 44752
rect 44272 44532 44324 44538
rect 44272 44474 44324 44480
rect 1490 44432 1546 44441
rect 1490 44367 1546 44376
rect 45192 44396 45244 44402
rect 45192 44338 45244 44344
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 43536 43784 43588 43790
rect 1490 43752 1546 43761
rect 43536 43726 43588 43732
rect 1490 43687 1546 43696
rect 1504 43654 1532 43687
rect 1492 43648 1544 43654
rect 1492 43590 1544 43596
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 43548 43450 43576 43726
rect 44272 43648 44324 43654
rect 44272 43590 44324 43596
rect 43536 43444 43588 43450
rect 43536 43386 43588 43392
rect 44284 43314 44312 43590
rect 44272 43308 44324 43314
rect 44272 43250 44324 43256
rect 1492 43104 1544 43110
rect 1490 43072 1492 43081
rect 2320 43104 2372 43110
rect 1544 43072 1546 43081
rect 2320 43046 2372 43052
rect 1490 43007 1546 43016
rect 2332 42702 2360 43046
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 2320 42696 2372 42702
rect 2320 42638 2372 42644
rect 42524 42628 42576 42634
rect 42524 42570 42576 42576
rect 1492 42560 1544 42566
rect 1492 42502 1544 42508
rect 1504 42401 1532 42502
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 1490 42392 1546 42401
rect 19574 42395 19882 42404
rect 42536 42362 42564 42570
rect 44180 42560 44232 42566
rect 44180 42502 44232 42508
rect 1490 42327 1546 42336
rect 42524 42356 42576 42362
rect 42524 42298 42576 42304
rect 43352 42220 43404 42226
rect 43352 42162 43404 42168
rect 41328 42084 41380 42090
rect 41328 42026 41380 42032
rect 1492 42016 1544 42022
rect 1492 41958 1544 41964
rect 1504 41721 1532 41958
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 41340 41750 41368 42026
rect 41328 41744 41380 41750
rect 1490 41712 1546 41721
rect 41328 41686 41380 41692
rect 1490 41647 1546 41656
rect 42616 41608 42668 41614
rect 42616 41550 42668 41556
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 1490 41032 1546 41041
rect 1490 40967 1492 40976
rect 1544 40967 1546 40976
rect 40684 40996 40736 41002
rect 1492 40938 1544 40944
rect 40684 40938 40736 40944
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 40696 40730 40724 40938
rect 42628 40934 42656 41550
rect 43364 41478 43392 42162
rect 43352 41472 43404 41478
rect 43352 41414 43404 41420
rect 41420 40928 41472 40934
rect 41420 40870 41472 40876
rect 42616 40928 42668 40934
rect 42616 40870 42668 40876
rect 40684 40724 40736 40730
rect 40684 40666 40736 40672
rect 41432 40458 41460 40870
rect 41420 40452 41472 40458
rect 41420 40394 41472 40400
rect 1492 40384 1544 40390
rect 1490 40352 1492 40361
rect 2320 40384 2372 40390
rect 1544 40352 1546 40361
rect 2320 40326 2372 40332
rect 41052 40384 41104 40390
rect 41052 40326 41104 40332
rect 1490 40287 1546 40296
rect 2332 39982 2360 40326
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 41064 40050 41092 40326
rect 40592 40044 40644 40050
rect 40592 39986 40644 39992
rect 41052 40044 41104 40050
rect 41052 39986 41104 39992
rect 2320 39976 2372 39982
rect 2320 39918 2372 39924
rect 39120 39908 39172 39914
rect 39120 39850 39172 39856
rect 1492 39840 1544 39846
rect 1492 39782 1544 39788
rect 1504 39681 1532 39782
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 1490 39672 1546 39681
rect 4214 39675 4522 39684
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 39132 39642 39160 39850
rect 1490 39607 1546 39616
rect 39120 39636 39172 39642
rect 39120 39578 39172 39584
rect 38384 39364 38436 39370
rect 38384 39306 38436 39312
rect 39856 39364 39908 39370
rect 39856 39306 39908 39312
rect 1492 39296 1544 39302
rect 1492 39238 1544 39244
rect 1504 39001 1532 39238
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 38396 39098 38424 39306
rect 38384 39092 38436 39098
rect 38384 39034 38436 39040
rect 1490 38992 1546 39001
rect 1490 38927 1546 38936
rect 39120 38956 39172 38962
rect 39120 38898 39172 38904
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 1490 38312 1546 38321
rect 1490 38247 1546 38256
rect 37740 38276 37792 38282
rect 1504 38214 1532 38247
rect 37740 38218 37792 38224
rect 1492 38208 1544 38214
rect 1492 38150 1544 38156
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 37752 38010 37780 38218
rect 39132 38214 39160 38898
rect 39868 38758 39896 39306
rect 40604 39302 40632 39986
rect 41432 39846 41460 40394
rect 41420 39840 41472 39846
rect 41420 39782 41472 39788
rect 40592 39296 40644 39302
rect 40592 39238 40644 39244
rect 39856 38752 39908 38758
rect 39856 38694 39908 38700
rect 38384 38208 38436 38214
rect 38384 38150 38436 38156
rect 39120 38208 39172 38214
rect 39120 38150 39172 38156
rect 37740 38004 37792 38010
rect 37740 37946 37792 37952
rect 38396 37874 38424 38150
rect 38384 37868 38436 37874
rect 38384 37810 38436 37816
rect 37004 37732 37056 37738
rect 37004 37674 37056 37680
rect 1492 37664 1544 37670
rect 1490 37632 1492 37641
rect 1544 37632 1546 37641
rect 1490 37567 1546 37576
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 37016 37466 37044 37674
rect 37004 37460 37056 37466
rect 37004 37402 37056 37408
rect 38396 37398 38424 37810
rect 38384 37392 38436 37398
rect 38384 37334 38436 37340
rect 36268 37188 36320 37194
rect 36268 37130 36320 37136
rect 37648 37188 37700 37194
rect 37648 37130 37700 37136
rect 38016 37188 38068 37194
rect 38016 37130 38068 37136
rect 1492 37120 1544 37126
rect 1492 37062 1544 37068
rect 1504 36961 1532 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 1490 36952 1546 36961
rect 19574 36955 19882 36964
rect 36280 36922 36308 37130
rect 1490 36887 1546 36896
rect 36268 36916 36320 36922
rect 36268 36858 36320 36864
rect 35624 36780 35676 36786
rect 35624 36722 35676 36728
rect 36636 36780 36688 36786
rect 36636 36722 36688 36728
rect 37188 36780 37240 36786
rect 37188 36722 37240 36728
rect 1492 36576 1544 36582
rect 1492 36518 1544 36524
rect 1504 36281 1532 36518
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35636 36378 35664 36722
rect 35624 36372 35676 36378
rect 35624 36314 35676 36320
rect 1490 36272 1546 36281
rect 1490 36207 1546 36216
rect 36268 36100 36320 36106
rect 36268 36042 36320 36048
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 1490 35592 1546 35601
rect 1490 35527 1492 35536
rect 1544 35527 1546 35536
rect 34704 35556 34756 35562
rect 1492 35498 1544 35504
rect 34704 35498 34756 35504
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34716 35290 34744 35498
rect 36280 35494 36308 36042
rect 35716 35488 35768 35494
rect 35716 35430 35768 35436
rect 36268 35488 36320 35494
rect 36268 35430 36320 35436
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34704 35284 34756 35290
rect 34704 35226 34756 35232
rect 34152 35080 34204 35086
rect 34152 35022 34204 35028
rect 1492 34944 1544 34950
rect 1490 34912 1492 34921
rect 1544 34912 1546 34921
rect 1490 34847 1546 34856
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 34164 34746 34192 35022
rect 35728 35018 35756 35430
rect 34796 35012 34848 35018
rect 34796 34954 34848 34960
rect 35716 35012 35768 35018
rect 35716 34954 35768 34960
rect 34152 34740 34204 34746
rect 34152 34682 34204 34688
rect 34704 34604 34756 34610
rect 34704 34546 34756 34552
rect 2320 34536 2372 34542
rect 2320 34478 2372 34484
rect 1492 34400 1544 34406
rect 1492 34342 1544 34348
rect 1504 34241 1532 34342
rect 1490 34232 1546 34241
rect 1490 34167 1546 34176
rect 2332 33998 2360 34478
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 2320 33992 2372 33998
rect 2320 33934 2372 33940
rect 32680 33924 32732 33930
rect 32680 33866 32732 33872
rect 1492 33856 1544 33862
rect 1492 33798 1544 33804
rect 1504 33561 1532 33798
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 32692 33658 32720 33866
rect 34716 33862 34744 34546
rect 33968 33856 34020 33862
rect 33968 33798 34020 33804
rect 34704 33856 34756 33862
rect 34704 33798 34756 33804
rect 32680 33652 32732 33658
rect 32680 33594 32732 33600
rect 1490 33552 1546 33561
rect 1490 33487 1546 33496
rect 33232 33516 33284 33522
rect 33232 33458 33284 33464
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 1490 32872 1546 32881
rect 1490 32807 1546 32816
rect 32220 32836 32272 32842
rect 1504 32774 1532 32807
rect 32220 32778 32272 32784
rect 1492 32768 1544 32774
rect 1492 32710 1544 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 32232 32570 32260 32778
rect 33244 32774 33272 33458
rect 32956 32768 33008 32774
rect 32956 32710 33008 32716
rect 33232 32768 33284 32774
rect 33232 32710 33284 32716
rect 32220 32564 32272 32570
rect 32220 32506 32272 32512
rect 32968 32434 32996 32710
rect 31208 32428 31260 32434
rect 31208 32370 31260 32376
rect 32956 32428 33008 32434
rect 32956 32370 33008 32376
rect 1492 32224 1544 32230
rect 1490 32192 1492 32201
rect 1544 32192 1546 32201
rect 1490 32127 1546 32136
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 31220 32026 31248 32370
rect 31208 32020 31260 32026
rect 31208 31962 31260 31968
rect 32404 31952 32456 31958
rect 32404 31894 32456 31900
rect 2320 31816 2372 31822
rect 2320 31758 2372 31764
rect 1492 31680 1544 31686
rect 1492 31622 1544 31628
rect 1504 31521 1532 31622
rect 1490 31512 1546 31521
rect 1490 31447 1546 31456
rect 2332 31278 2360 31758
rect 31944 31748 31996 31754
rect 31944 31690 31996 31696
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 31668 31340 31720 31346
rect 31668 31282 31720 31288
rect 2320 31272 2372 31278
rect 2320 31214 2372 31220
rect 29736 31204 29788 31210
rect 29736 31146 29788 31152
rect 1492 31136 1544 31142
rect 1492 31078 1544 31084
rect 1504 30841 1532 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 29748 30938 29776 31146
rect 29736 30932 29788 30938
rect 29736 30874 29788 30880
rect 1490 30832 1546 30841
rect 1490 30767 1546 30776
rect 30380 30660 30432 30666
rect 30380 30602 30432 30608
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 1490 30152 1546 30161
rect 1490 30087 1492 30096
rect 1544 30087 1546 30096
rect 28816 30116 28868 30122
rect 1492 30058 1544 30064
rect 28816 30058 28868 30064
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 28828 29850 28856 30058
rect 30392 30054 30420 30602
rect 31680 30598 31708 31282
rect 31956 31142 31984 31690
rect 32416 31414 32444 31894
rect 32968 31822 32996 32370
rect 32588 31816 32640 31822
rect 32588 31758 32640 31764
rect 32956 31816 33008 31822
rect 32956 31758 33008 31764
rect 32404 31408 32456 31414
rect 32404 31350 32456 31356
rect 31944 31136 31996 31142
rect 31944 31078 31996 31084
rect 31024 30592 31076 30598
rect 31024 30534 31076 30540
rect 31668 30592 31720 30598
rect 31668 30534 31720 30540
rect 29368 30048 29420 30054
rect 29368 29990 29420 29996
rect 30380 30048 30432 30054
rect 30380 29990 30432 29996
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 28264 29640 28316 29646
rect 28264 29582 28316 29588
rect 1492 29504 1544 29510
rect 1490 29472 1492 29481
rect 1544 29472 1546 29481
rect 1490 29407 1546 29416
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 28276 29306 28304 29582
rect 29380 29510 29408 29990
rect 29368 29504 29420 29510
rect 29368 29446 29420 29452
rect 28264 29300 28316 29306
rect 28264 29242 28316 29248
rect 26148 29096 26200 29102
rect 26148 29038 26200 29044
rect 1492 29028 1544 29034
rect 1492 28970 1544 28976
rect 1504 28801 1532 28970
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 1490 28792 1546 28801
rect 4214 28795 4522 28804
rect 1490 28727 1546 28736
rect 26160 28694 26188 29038
rect 28724 29028 28776 29034
rect 28724 28970 28776 28976
rect 26148 28688 26200 28694
rect 26148 28630 26200 28636
rect 27068 28552 27120 28558
rect 27068 28494 27120 28500
rect 1492 28416 1544 28422
rect 1492 28358 1544 28364
rect 1504 28121 1532 28358
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 27080 28218 27108 28494
rect 27988 28416 28040 28422
rect 27988 28358 28040 28364
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 1490 28112 1546 28121
rect 1490 28047 1546 28056
rect 27436 28076 27488 28082
rect 27436 28018 27488 28024
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 26056 27464 26108 27470
rect 1490 27432 1546 27441
rect 26056 27406 26108 27412
rect 1490 27367 1546 27376
rect 1504 27334 1532 27367
rect 1492 27328 1544 27334
rect 1492 27270 1544 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 26068 27130 26096 27406
rect 27448 27334 27476 28018
rect 26148 27328 26200 27334
rect 26148 27270 26200 27276
rect 27436 27328 27488 27334
rect 27436 27270 27488 27276
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 26160 26994 26188 27270
rect 25228 26988 25280 26994
rect 25228 26930 25280 26936
rect 26148 26988 26200 26994
rect 26148 26930 26200 26936
rect 1492 26784 1544 26790
rect 1490 26752 1492 26761
rect 1544 26752 1546 26761
rect 1490 26687 1546 26696
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 25240 26586 25268 26930
rect 25228 26580 25280 26586
rect 25228 26522 25280 26528
rect 26160 26450 26188 26930
rect 26148 26444 26200 26450
rect 26148 26386 26200 26392
rect 22836 26376 22888 26382
rect 22836 26318 22888 26324
rect 1492 26240 1544 26246
rect 1492 26182 1544 26188
rect 1504 26081 1532 26182
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 1490 26072 1546 26081
rect 19574 26075 19882 26084
rect 1490 26007 1546 26016
rect 22848 25974 22876 26318
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 22836 25968 22888 25974
rect 22836 25910 22888 25916
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 22284 25764 22336 25770
rect 22284 25706 22336 25712
rect 1492 25696 1544 25702
rect 1492 25638 1544 25644
rect 1504 25401 1532 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 22296 25498 22324 25706
rect 22284 25492 22336 25498
rect 22284 25434 22336 25440
rect 1490 25392 1546 25401
rect 1490 25327 1546 25336
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 24412 24886 24440 25230
rect 24400 24880 24452 24886
rect 24400 24822 24452 24828
rect 22284 24812 22336 24818
rect 22284 24754 22336 24760
rect 1490 24712 1546 24721
rect 1490 24647 1492 24656
rect 1544 24647 1546 24656
rect 1492 24618 1544 24624
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 22296 24410 22324 24754
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 1492 24064 1544 24070
rect 1490 24032 1492 24041
rect 1544 24032 1546 24041
rect 1490 23967 1546 23976
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 21836 23866 21864 24142
rect 23664 24132 23716 24138
rect 23664 24074 23716 24080
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 1492 23520 1544 23526
rect 1492 23462 1544 23468
rect 1504 23361 1532 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 1490 23352 1546 23361
rect 4214 23355 4522 23364
rect 19720 23322 19748 23530
rect 22572 23526 22600 23666
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 1490 23287 1546 23296
rect 19708 23316 19760 23322
rect 19708 23258 19760 23264
rect 22572 23118 22600 23462
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 1492 22976 1544 22982
rect 1492 22918 1544 22924
rect 1504 22681 1532 22918
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22778 20024 22986
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 1490 22672 1546 22681
rect 1490 22607 1546 22616
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 19064 22024 19116 22030
rect 1490 21992 1546 22001
rect 19064 21966 19116 21972
rect 1490 21927 1546 21936
rect 1504 21894 1532 21927
rect 1492 21888 1544 21894
rect 1492 21830 1544 21836
rect 19076 21690 19104 21966
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 1492 21344 1544 21350
rect 1490 21312 1492 21321
rect 1544 21312 1546 21321
rect 1490 21247 1546 21256
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 17880 21146 17908 21490
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 20641 1532 20742
rect 1490 20632 1546 20641
rect 17972 20602 18000 20878
rect 1490 20567 1546 20576
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1504 19961 1532 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 17052 20058 17080 20402
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 1490 19952 1546 19961
rect 1490 19887 1546 19896
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17972 19378 18000 19654
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 1490 19272 1546 19281
rect 1490 19207 1492 19216
rect 1544 19207 1546 19216
rect 1492 19178 1544 19184
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 1492 18624 1544 18630
rect 1490 18592 1492 18601
rect 16856 18624 16908 18630
rect 1544 18592 1546 18601
rect 16856 18566 16908 18572
rect 1490 18527 1546 18536
rect 16868 18426 16896 18566
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17921 1532 18022
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 1490 17912 1546 17921
rect 4214 17915 4522 17924
rect 12360 17882 12388 18226
rect 1490 17847 1546 17856
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 14476 17338 14504 17614
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 12716 16584 12768 16590
rect 1490 16552 1546 16561
rect 12716 16526 12768 16532
rect 1490 16487 1546 16496
rect 1504 16454 1532 16487
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 12728 16250 12756 16526
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 1492 15904 1544 15910
rect 1490 15872 1492 15881
rect 1544 15872 1546 15881
rect 1490 15807 1546 15816
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 11532 15162 11560 15438
rect 13832 15366 13860 15982
rect 14108 15910 14136 16050
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14108 15706 14136 15846
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 1490 15127 1546 15136
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14521 1532 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 11532 14618 11560 14962
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 1490 14512 1546 14521
rect 1490 14447 1546 14456
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 14074 12664 14214
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 11888 13864 11940 13870
rect 1490 13832 1546 13841
rect 11888 13806 11940 13812
rect 1490 13767 1492 13776
rect 1544 13767 1546 13776
rect 1492 13738 1544 13744
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 1492 13184 1544 13190
rect 1490 13152 1492 13161
rect 1544 13152 1546 13161
rect 1490 13087 1546 13096
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12481 1532 12582
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 1490 12472 1546 12481
rect 4214 12475 4522 12484
rect 9692 12442 9720 12786
rect 1490 12407 1546 12416
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11801 1532 12038
rect 9048 11898 9076 12174
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 1490 11792 1546 11801
rect 1490 11727 1546 11736
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 1492 11280 1544 11286
rect 1492 11222 1544 11228
rect 1504 11121 1532 11222
rect 8300 11144 8352 11150
rect 1490 11112 1546 11121
rect 8300 11086 8352 11092
rect 1490 11047 1546 11056
rect 8312 10810 8340 11086
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 1492 10464 1544 10470
rect 1490 10432 1492 10441
rect 1544 10432 1546 10441
rect 1490 10367 1546 10376
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 7576 10266 7604 10610
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9761 1532 9862
rect 1490 9752 1546 9761
rect 6748 9722 6776 9998
rect 1490 9687 1546 9696
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1504 9081 1532 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 6012 9178 6040 9522
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 1490 8392 1546 8401
rect 1490 8327 1492 8336
rect 1544 8327 1546 8336
rect 1492 8298 1544 8304
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 5276 8090 5304 8434
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 1492 7744 1544 7750
rect 1490 7712 1492 7721
rect 1544 7712 1546 7721
rect 1490 7647 1546 7656
rect 4540 7546 4568 7822
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 7041 1532 7142
rect 1490 7032 1546 7041
rect 3896 7002 3924 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1490 6967 1546 6976
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6361 1532 6598
rect 3252 6458 3280 6734
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 1490 6352 1546 6361
rect 1490 6287 1546 6296
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 1676 5704 1728 5710
rect 1490 5672 1546 5681
rect 1676 5646 1728 5652
rect 1490 5607 1546 5616
rect 1504 5574 1532 5607
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1688 5370 1716 5646
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 1492 5024 1544 5030
rect 1490 4992 1492 5001
rect 1544 4992 1546 5001
rect 1490 4927 1546 4936
rect 2056 4826 2084 5170
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2332 2650 2360 4558
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2792 2446 2820 2790
rect 3068 2650 3096 5170
rect 3804 3194 3832 6258
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2056 800 2084 2382
rect 2792 800 2820 2382
rect 3528 800 3556 2994
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 6734
rect 4724 2650 4752 7346
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5000 2446 5028 2790
rect 5644 2650 5672 7822
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5736 2446 5764 2790
rect 6196 2650 6224 8910
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6656 5370 6684 5646
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6472 2446 6500 2790
rect 6932 2650 6960 9522
rect 7196 2848 7248 2854
rect 7196 2790 7248 2796
rect 7932 2848 7984 2854
rect 7932 2790 7984 2796
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7208 2446 7236 2790
rect 7944 2446 7972 2790
rect 8220 2650 8248 9998
rect 8956 3194 8984 10610
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 4264 800 4292 2382
rect 5000 800 5028 2382
rect 5736 800 5764 2382
rect 6472 800 6500 2382
rect 7208 800 7236 2382
rect 7944 800 7972 2382
rect 8680 800 8708 2994
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9416 2446 9444 2790
rect 9600 2650 9628 11698
rect 10060 2650 10088 12174
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10152 2446 10180 2790
rect 10796 2650 10824 13194
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 11716 10810 11744 11018
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10980 9722 11008 9862
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10888 2446 10916 2790
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 9416 800 9444 2382
rect 10152 800 10180 2382
rect 10888 800 10916 2382
rect 11624 2378 11652 2790
rect 11900 2650 11928 13806
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11612 2372 11664 2378
rect 11612 2314 11664 2320
rect 12360 2360 12388 2790
rect 12636 2650 12664 14010
rect 13372 13938 13400 14758
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 13096 2378 13124 2790
rect 13372 2650 13400 13874
rect 14108 3194 14136 15642
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13360 2644 13412 2650
rect 13360 2586 13412 2592
rect 12440 2372 12492 2378
rect 12360 2332 12440 2360
rect 11624 800 11652 2314
rect 12360 800 12388 2332
rect 12440 2314 12492 2320
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 13096 800 13124 2314
rect 13832 800 13860 2994
rect 14476 2650 14504 15302
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14568 2378 14596 2790
rect 15120 2582 15148 16934
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15304 2378 15332 2790
rect 15948 2650 15976 17478
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16040 2378 16068 2790
rect 16776 2378 16804 2790
rect 17052 2650 17080 18362
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 17512 2378 17540 2790
rect 17788 2650 17816 19110
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 18248 2378 18276 2790
rect 18524 2650 18552 19314
rect 19352 18698 19380 20198
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19352 3126 19380 18634
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 16028 2372 16080 2378
rect 16028 2314 16080 2320
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 17500 2372 17552 2378
rect 17500 2314 17552 2320
rect 18236 2372 18288 2378
rect 18236 2314 18288 2320
rect 14568 800 14596 2314
rect 15304 800 15332 2314
rect 16040 800 16068 2314
rect 16776 800 16804 2314
rect 17512 800 17540 2314
rect 18248 800 18276 2314
rect 18984 800 19012 2994
rect 19444 2582 19472 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20364 18086 20392 21286
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19996 2378 20024 2790
rect 20364 2650 20392 18022
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 20352 2644 20404 2650
rect 20352 2586 20404 2592
rect 20456 2378 20484 2790
rect 21192 2378 21220 2790
rect 21928 2428 21956 2790
rect 22100 2440 22152 2446
rect 21928 2400 22100 2428
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 20444 2372 20496 2378
rect 20444 2314 20496 2320
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19720 870 19840 898
rect 19720 800 19748 870
rect 2042 0 2098 800
rect 2778 0 2834 800
rect 3514 0 3570 800
rect 4250 0 4306 800
rect 4986 0 5042 800
rect 5722 0 5778 800
rect 6458 0 6514 800
rect 7194 0 7250 800
rect 7930 0 7986 800
rect 8666 0 8722 800
rect 9402 0 9458 800
rect 10138 0 10194 800
rect 10874 0 10930 800
rect 11610 0 11666 800
rect 12346 0 12402 800
rect 13082 0 13138 800
rect 13818 0 13874 800
rect 14554 0 14610 800
rect 15290 0 15346 800
rect 16026 0 16082 800
rect 16762 0 16818 800
rect 17498 0 17554 800
rect 18234 0 18290 800
rect 18970 0 19026 800
rect 19706 0 19762 800
rect 19812 762 19840 870
rect 19996 762 20024 2314
rect 20456 800 20484 2314
rect 21192 800 21220 2314
rect 21928 800 21956 2400
rect 22100 2382 22152 2388
rect 22664 2378 22692 2790
rect 22940 2650 22968 23054
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 23400 2428 23428 2790
rect 23676 2650 23704 24074
rect 24412 3194 24440 24822
rect 24964 23322 24992 25842
rect 26068 25702 26096 26182
rect 26056 25696 26108 25702
rect 26056 25638 26108 25644
rect 24952 23316 25004 23322
rect 24952 23258 25004 23264
rect 24400 3188 24452 3194
rect 24400 3130 24452 3136
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23480 2440 23532 2446
rect 23400 2400 23480 2428
rect 22652 2372 22704 2378
rect 22652 2314 22704 2320
rect 22664 800 22692 2314
rect 23400 800 23428 2400
rect 23480 2382 23532 2388
rect 24136 800 24164 2994
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 24872 2378 24900 2790
rect 24964 2650 24992 23258
rect 26068 3058 26096 25638
rect 26056 3052 26108 3058
rect 26056 2994 26108 3000
rect 25596 2984 25648 2990
rect 25596 2926 25648 2932
rect 24952 2644 25004 2650
rect 24952 2586 25004 2592
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 24872 800 24900 2314
rect 25608 800 25636 2926
rect 26160 2514 26188 26386
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 26976 22432 27028 22438
rect 26976 22374 27028 22380
rect 26332 18624 26384 18630
rect 26332 18566 26384 18572
rect 26344 18154 26372 18566
rect 26988 18290 27016 22374
rect 27068 20800 27120 20806
rect 27068 20742 27120 20748
rect 27080 18630 27108 20742
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 26516 18284 26568 18290
rect 26516 18226 26568 18232
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 26332 18148 26384 18154
rect 26332 18090 26384 18096
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 26252 16454 26280 16934
rect 26240 16448 26292 16454
rect 26240 16390 26292 16396
rect 26252 16250 26280 16390
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26344 2582 26372 18090
rect 26528 17542 26556 18226
rect 27080 18086 27108 18566
rect 27172 18222 27200 22918
rect 27344 21956 27396 21962
rect 27344 21898 27396 21904
rect 27356 18290 27384 21898
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 27344 17672 27396 17678
rect 27344 17614 27396 17620
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26516 17536 26568 17542
rect 26516 17478 26568 17484
rect 26436 17202 26464 17478
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26436 16794 26464 17138
rect 26424 16788 26476 16794
rect 26424 16730 26476 16736
rect 26436 16046 26464 16730
rect 26424 16040 26476 16046
rect 26424 15982 26476 15988
rect 26332 2576 26384 2582
rect 26332 2518 26384 2524
rect 26148 2508 26200 2514
rect 26148 2450 26200 2456
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 26344 800 26372 2382
rect 26528 2310 26556 17478
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 26976 14340 27028 14346
rect 26976 14282 27028 14288
rect 26988 14074 27016 14282
rect 26976 14068 27028 14074
rect 26976 14010 27028 14016
rect 26988 13734 27016 14010
rect 27080 13938 27108 14962
rect 27356 14074 27384 17614
rect 27344 14068 27396 14074
rect 27344 14010 27396 14016
rect 27068 13932 27120 13938
rect 27068 13874 27120 13880
rect 26976 13728 27028 13734
rect 26976 13670 27028 13676
rect 26988 13530 27016 13670
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 27448 6914 27476 27270
rect 27712 18080 27764 18086
rect 27712 18022 27764 18028
rect 27724 17746 27752 18022
rect 27712 17740 27764 17746
rect 27712 17682 27764 17688
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27540 16250 27568 17614
rect 27528 16244 27580 16250
rect 27528 16186 27580 16192
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 27632 15638 27660 16118
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 27724 15706 27752 15846
rect 27712 15700 27764 15706
rect 27712 15642 27764 15648
rect 27620 15632 27672 15638
rect 27620 15574 27672 15580
rect 27804 15428 27856 15434
rect 27804 15370 27856 15376
rect 27816 15094 27844 15370
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 27896 13932 27948 13938
rect 27896 13874 27948 13880
rect 27908 13530 27936 13874
rect 27896 13524 27948 13530
rect 27896 13466 27948 13472
rect 27448 6886 27568 6914
rect 27540 3602 27568 6886
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27068 3528 27120 3534
rect 27068 3470 27120 3476
rect 26516 2304 26568 2310
rect 26516 2246 26568 2252
rect 27080 800 27108 3470
rect 28000 3058 28028 28358
rect 28172 16992 28224 16998
rect 28172 16934 28224 16940
rect 28184 16590 28212 16934
rect 28172 16584 28224 16590
rect 28172 16526 28224 16532
rect 28184 16182 28212 16526
rect 28172 16176 28224 16182
rect 28172 16118 28224 16124
rect 28448 3392 28500 3398
rect 28448 3334 28500 3340
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 28460 2990 28488 3334
rect 27804 2984 27856 2990
rect 27804 2926 27856 2932
rect 28448 2984 28500 2990
rect 28448 2926 28500 2932
rect 27816 800 27844 2926
rect 28736 2514 28764 28970
rect 29276 3460 29328 3466
rect 29276 3402 29328 3408
rect 29288 2990 29316 3402
rect 29380 3058 29408 29446
rect 30288 23316 30340 23322
rect 30288 23258 30340 23264
rect 30300 22982 30328 23258
rect 30288 22976 30340 22982
rect 30288 22918 30340 22924
rect 30012 3392 30064 3398
rect 30012 3334 30064 3340
rect 29368 3052 29420 3058
rect 29368 2994 29420 3000
rect 30024 2990 30052 3334
rect 30392 3058 30420 29990
rect 30840 25152 30892 25158
rect 30840 25094 30892 25100
rect 30852 24886 30880 25094
rect 30840 24880 30892 24886
rect 30840 24822 30892 24828
rect 30852 23866 30880 24822
rect 30840 23860 30892 23866
rect 30840 23802 30892 23808
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 30944 19378 30972 19654
rect 30932 19372 30984 19378
rect 30932 19314 30984 19320
rect 30656 18828 30708 18834
rect 30656 18770 30708 18776
rect 30668 18714 30696 18770
rect 30944 18766 30972 19314
rect 30484 18698 30696 18714
rect 30932 18760 30984 18766
rect 30932 18702 30984 18708
rect 30472 18692 30696 18698
rect 30524 18686 30696 18692
rect 30472 18634 30524 18640
rect 30564 18624 30616 18630
rect 30564 18566 30616 18572
rect 30576 18426 30604 18566
rect 30564 18420 30616 18426
rect 30564 18362 30616 18368
rect 30380 3052 30432 3058
rect 30380 2994 30432 3000
rect 29276 2984 29328 2990
rect 29276 2926 29328 2932
rect 30012 2984 30064 2990
rect 30012 2926 30064 2932
rect 28724 2508 28776 2514
rect 28724 2450 28776 2456
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 28552 800 28580 2382
rect 29288 800 29316 2926
rect 30024 800 30052 2926
rect 31036 2514 31064 30534
rect 31668 25968 31720 25974
rect 31668 25910 31720 25916
rect 31576 23860 31628 23866
rect 31576 23802 31628 23808
rect 31392 23724 31444 23730
rect 31392 23666 31444 23672
rect 31484 23724 31536 23730
rect 31484 23666 31536 23672
rect 31404 18970 31432 23666
rect 31496 23322 31524 23666
rect 31588 23322 31616 23802
rect 31484 23316 31536 23322
rect 31484 23258 31536 23264
rect 31576 23316 31628 23322
rect 31576 23258 31628 23264
rect 31680 23118 31708 25910
rect 31668 23112 31720 23118
rect 31668 23054 31720 23060
rect 31680 22982 31708 23054
rect 31668 22976 31720 22982
rect 31668 22918 31720 22924
rect 31484 20460 31536 20466
rect 31484 20402 31536 20408
rect 31496 20262 31524 20402
rect 31484 20256 31536 20262
rect 31484 20198 31536 20204
rect 31392 18964 31444 18970
rect 31392 18906 31444 18912
rect 31496 18834 31524 20198
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31772 19174 31800 19314
rect 31760 19168 31812 19174
rect 31760 19110 31812 19116
rect 31484 18828 31536 18834
rect 31484 18770 31536 18776
rect 31772 18766 31800 19110
rect 31760 18760 31812 18766
rect 31760 18702 31812 18708
rect 31772 18358 31800 18702
rect 31760 18352 31812 18358
rect 31760 18294 31812 18300
rect 31484 2848 31536 2854
rect 31484 2790 31536 2796
rect 31024 2508 31076 2514
rect 31024 2450 31076 2456
rect 31496 2446 31524 2790
rect 31956 2514 31984 31078
rect 32600 26234 32628 31758
rect 32508 26206 32628 26234
rect 32680 26240 32732 26246
rect 32036 24132 32088 24138
rect 32036 24074 32088 24080
rect 32048 23118 32076 24074
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 32036 23112 32088 23118
rect 32036 23054 32088 23060
rect 32048 22778 32076 23054
rect 32232 23050 32260 23666
rect 32220 23044 32272 23050
rect 32220 22986 32272 22992
rect 32036 22772 32088 22778
rect 32036 22714 32088 22720
rect 32404 20936 32456 20942
rect 32404 20878 32456 20884
rect 32416 20534 32444 20878
rect 32404 20528 32456 20534
rect 32404 20470 32456 20476
rect 32220 3392 32272 3398
rect 32220 3334 32272 3340
rect 32232 3058 32260 3334
rect 32508 3194 32536 26206
rect 32680 26182 32732 26188
rect 32692 25974 32720 26182
rect 32680 25968 32732 25974
rect 32680 25910 32732 25916
rect 32956 3392 33008 3398
rect 32956 3334 33008 3340
rect 32496 3188 32548 3194
rect 32496 3130 32548 3136
rect 32968 3058 32996 3334
rect 33244 3194 33272 32710
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33232 3188 33284 3194
rect 33232 3130 33284 3136
rect 32220 3052 32272 3058
rect 32220 2994 32272 3000
rect 32956 3052 33008 3058
rect 32956 2994 33008 3000
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 31484 2440 31536 2446
rect 31484 2382 31536 2388
rect 30760 800 30788 2382
rect 31496 800 31524 2382
rect 32232 800 32260 2994
rect 32968 800 32996 2994
rect 33704 2378 33732 3334
rect 33980 2650 34008 33798
rect 34716 3194 34744 33798
rect 34704 3188 34756 3194
rect 34704 3130 34756 3136
rect 34428 3052 34480 3058
rect 34428 2994 34480 3000
rect 33968 2644 34020 2650
rect 33968 2586 34020 2592
rect 33692 2372 33744 2378
rect 33692 2314 33744 2320
rect 33704 800 33732 2314
rect 34440 800 34468 2994
rect 34808 2582 34836 34954
rect 35728 34746 35756 34954
rect 35716 34740 35768 34746
rect 35716 34682 35768 34688
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 35900 2848 35952 2854
rect 35900 2790 35952 2796
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2576 34848 2582
rect 34796 2518 34848 2524
rect 35164 2372 35216 2378
rect 35360 2360 35388 2790
rect 35912 2378 35940 2790
rect 36280 2650 36308 35430
rect 36648 26234 36676 36722
rect 37200 36378 37228 36722
rect 37188 36372 37240 36378
rect 37188 36314 37240 36320
rect 36556 26206 36676 26234
rect 36556 2650 36584 26206
rect 37188 23724 37240 23730
rect 37188 23666 37240 23672
rect 37200 17542 37228 23666
rect 37188 17536 37240 17542
rect 37188 17478 37240 17484
rect 36636 2848 36688 2854
rect 36636 2790 36688 2796
rect 37372 2848 37424 2854
rect 37372 2790 37424 2796
rect 36268 2644 36320 2650
rect 36268 2586 36320 2592
rect 36544 2644 36596 2650
rect 36544 2586 36596 2592
rect 36648 2378 36676 2790
rect 37384 2378 37412 2790
rect 37660 2650 37688 37130
rect 38028 36922 38056 37130
rect 38016 36916 38068 36922
rect 38016 36858 38068 36864
rect 38108 2848 38160 2854
rect 38108 2790 38160 2796
rect 37648 2644 37700 2650
rect 37648 2586 37700 2592
rect 38120 2378 38148 2790
rect 38396 2650 38424 37334
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 38384 2644 38436 2650
rect 38384 2586 38436 2592
rect 38856 2378 38884 2790
rect 39132 2650 39160 38150
rect 39868 3194 39896 38694
rect 39856 3188 39908 3194
rect 39856 3130 39908 3136
rect 39580 3052 39632 3058
rect 39580 2994 39632 3000
rect 39120 2644 39172 2650
rect 39120 2586 39172 2592
rect 35216 2332 35388 2360
rect 35900 2372 35952 2378
rect 35164 2314 35216 2320
rect 35900 2314 35952 2320
rect 36636 2372 36688 2378
rect 36636 2314 36688 2320
rect 37372 2372 37424 2378
rect 37372 2314 37424 2320
rect 38108 2372 38160 2378
rect 38108 2314 38160 2320
rect 38844 2372 38896 2378
rect 38844 2314 38896 2320
rect 35176 800 35204 2314
rect 35912 800 35940 2314
rect 36648 800 36676 2314
rect 37384 800 37412 2314
rect 38120 800 38148 2314
rect 38856 800 38884 2314
rect 39592 800 39620 2994
rect 40604 2650 40632 39238
rect 41052 2848 41104 2854
rect 41052 2790 41104 2796
rect 40592 2644 40644 2650
rect 40592 2586 40644 2592
rect 41064 2378 41092 2790
rect 41432 2582 41460 39782
rect 41512 24812 41564 24818
rect 41512 24754 41564 24760
rect 41524 24138 41552 24754
rect 41696 24676 41748 24682
rect 41696 24618 41748 24624
rect 41604 24608 41656 24614
rect 41604 24550 41656 24556
rect 41616 24410 41644 24550
rect 41604 24404 41656 24410
rect 41604 24346 41656 24352
rect 41512 24132 41564 24138
rect 41512 24074 41564 24080
rect 41524 23526 41552 24074
rect 41616 23594 41644 24346
rect 41708 24070 41736 24618
rect 41696 24064 41748 24070
rect 41696 24006 41748 24012
rect 41708 23730 41736 24006
rect 41696 23724 41748 23730
rect 41696 23666 41748 23672
rect 41604 23588 41656 23594
rect 41604 23530 41656 23536
rect 41512 23520 41564 23526
rect 41512 23462 41564 23468
rect 41524 13190 41552 23462
rect 41512 13184 41564 13190
rect 41512 13126 41564 13132
rect 42432 2848 42484 2854
rect 42432 2790 42484 2796
rect 41420 2576 41472 2582
rect 41420 2518 41472 2524
rect 42444 2378 42472 2790
rect 42628 2650 42656 40870
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 42616 2644 42668 2650
rect 42616 2586 42668 2592
rect 42812 2378 42840 2790
rect 43364 2650 43392 41414
rect 43720 3392 43772 3398
rect 43720 3334 43772 3340
rect 43352 2644 43404 2650
rect 43352 2586 43404 2592
rect 43732 2378 43760 3334
rect 43996 3052 44048 3058
rect 43996 2994 44048 3000
rect 40316 2372 40368 2378
rect 40316 2314 40368 2320
rect 41052 2372 41104 2378
rect 41052 2314 41104 2320
rect 41788 2372 41840 2378
rect 41788 2314 41840 2320
rect 42432 2372 42484 2378
rect 42432 2314 42484 2320
rect 42800 2372 42852 2378
rect 43352 2372 43404 2378
rect 42800 2314 42852 2320
rect 43272 2332 43352 2360
rect 40328 800 40356 2314
rect 41064 800 41092 2314
rect 41800 800 41828 2314
rect 42812 2258 42840 2314
rect 42536 2230 42840 2258
rect 42536 800 42564 2230
rect 43272 800 43300 2332
rect 43352 2314 43404 2320
rect 43720 2372 43772 2378
rect 43720 2314 43772 2320
rect 44008 800 44036 2994
rect 44192 2582 44220 42502
rect 44284 3194 44312 43250
rect 44272 3188 44324 3194
rect 44272 3130 44324 3136
rect 44732 2848 44784 2854
rect 44732 2790 44784 2796
rect 44180 2576 44232 2582
rect 44180 2518 44232 2524
rect 44744 2378 44772 2790
rect 45204 2650 45232 44338
rect 45940 44198 45968 44746
rect 45928 44192 45980 44198
rect 45928 44134 45980 44140
rect 45652 2848 45704 2854
rect 45652 2790 45704 2796
rect 45192 2644 45244 2650
rect 45192 2586 45244 2592
rect 45664 2446 45692 2790
rect 45940 2650 45968 44134
rect 46204 2848 46256 2854
rect 46204 2790 46256 2796
rect 45928 2644 45980 2650
rect 45928 2586 45980 2592
rect 45652 2440 45704 2446
rect 45652 2382 45704 2388
rect 44732 2372 44784 2378
rect 44732 2314 44784 2320
rect 44744 800 44772 2314
rect 45664 2258 45692 2382
rect 46216 2378 46244 2790
rect 46676 2650 46704 45426
rect 47596 6914 47624 45526
rect 47504 6886 47624 6914
rect 46664 2644 46716 2650
rect 46664 2586 46716 2592
rect 47504 2582 47532 6886
rect 47584 2848 47636 2854
rect 47584 2790 47636 2796
rect 47676 2848 47728 2854
rect 47676 2790 47728 2796
rect 47492 2576 47544 2582
rect 47492 2518 47544 2524
rect 47596 2378 47624 2790
rect 46204 2372 46256 2378
rect 46204 2314 46256 2320
rect 46940 2372 46992 2378
rect 46940 2314 46992 2320
rect 47584 2372 47636 2378
rect 47584 2314 47636 2320
rect 45480 2230 45692 2258
rect 45480 800 45508 2230
rect 46216 800 46244 2314
rect 46952 800 46980 2314
rect 47688 800 47716 2790
rect 47780 2650 47808 45902
rect 48412 2848 48464 2854
rect 48412 2790 48464 2796
rect 48780 2848 48832 2854
rect 48780 2790 48832 2796
rect 49148 2848 49200 2854
rect 49148 2790 49200 2796
rect 47768 2644 47820 2650
rect 47768 2586 47820 2592
rect 48424 2446 48452 2790
rect 48412 2440 48464 2446
rect 48412 2382 48464 2388
rect 48792 2378 48820 2790
rect 48780 2372 48832 2378
rect 48780 2314 48832 2320
rect 48412 2304 48464 2310
rect 48412 2246 48464 2252
rect 48424 800 48452 2246
rect 49160 800 49188 2790
rect 49252 2650 49280 47398
rect 49988 3194 50016 48486
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50632 3194 50660 49302
rect 50724 49230 50752 49778
rect 51264 49768 51316 49774
rect 51264 49710 51316 49716
rect 50712 49224 50764 49230
rect 50712 49166 50764 49172
rect 50724 48754 50752 49166
rect 50712 48748 50764 48754
rect 50712 48690 50764 48696
rect 51276 3194 51304 49710
rect 51828 3194 51856 50390
rect 49976 3188 50028 3194
rect 49976 3130 50028 3136
rect 50620 3188 50672 3194
rect 50620 3130 50672 3136
rect 51264 3188 51316 3194
rect 51264 3130 51316 3136
rect 51816 3188 51868 3194
rect 51816 3130 51868 3136
rect 49240 2644 49292 2650
rect 49240 2586 49292 2592
rect 50632 2446 50660 3130
rect 51276 2446 51304 3130
rect 51828 2446 51856 3130
rect 52104 3126 52132 51750
rect 52196 51406 52224 51954
rect 53116 51950 53144 54674
rect 56612 54670 56640 55082
rect 56704 54738 56732 55218
rect 56692 54732 56744 54738
rect 56692 54674 56744 54680
rect 56600 54664 56652 54670
rect 56600 54606 56652 54612
rect 53380 54596 53432 54602
rect 53380 54538 53432 54544
rect 53288 53508 53340 53514
rect 53288 53450 53340 53456
rect 53300 53174 53328 53450
rect 53288 53168 53340 53174
rect 53288 53110 53340 53116
rect 53196 53100 53248 53106
rect 53196 53042 53248 53048
rect 53208 52970 53236 53042
rect 53196 52964 53248 52970
rect 53196 52906 53248 52912
rect 53208 52018 53236 52906
rect 53288 52896 53340 52902
rect 53288 52838 53340 52844
rect 53196 52012 53248 52018
rect 53196 51954 53248 51960
rect 53104 51944 53156 51950
rect 53104 51886 53156 51892
rect 52368 51536 52420 51542
rect 52368 51478 52420 51484
rect 52184 51400 52236 51406
rect 52184 51342 52236 51348
rect 52380 3194 52408 51478
rect 53116 51474 53144 51886
rect 53104 51468 53156 51474
rect 53104 51410 53156 51416
rect 53012 51400 53064 51406
rect 53012 51342 53064 51348
rect 52736 50312 52788 50318
rect 52736 50254 52788 50260
rect 52748 50182 52776 50254
rect 53024 50250 53052 51342
rect 53012 50244 53064 50250
rect 53012 50186 53064 50192
rect 52736 50176 52788 50182
rect 52736 50118 52788 50124
rect 52748 49978 52776 50118
rect 52736 49972 52788 49978
rect 52736 49914 52788 49920
rect 53300 3194 53328 52838
rect 53392 52494 53420 54538
rect 55496 54528 55548 54534
rect 55496 54470 55548 54476
rect 55508 54330 55536 54470
rect 55496 54324 55548 54330
rect 55496 54266 55548 54272
rect 56612 54262 56640 54606
rect 56600 54256 56652 54262
rect 56600 54198 56652 54204
rect 56704 54194 56732 54674
rect 56692 54188 56744 54194
rect 56692 54130 56744 54136
rect 56600 53984 56652 53990
rect 56600 53926 56652 53932
rect 54116 53440 54168 53446
rect 54116 53382 54168 53388
rect 54128 53106 54156 53382
rect 53840 53100 53892 53106
rect 53840 53042 53892 53048
rect 54116 53100 54168 53106
rect 54116 53042 54168 53048
rect 53852 52494 53880 53042
rect 55220 52896 55272 52902
rect 55220 52838 55272 52844
rect 53380 52488 53432 52494
rect 53380 52430 53432 52436
rect 53840 52488 53892 52494
rect 53840 52430 53892 52436
rect 53392 50930 53420 52430
rect 53852 52018 53880 52430
rect 55036 52352 55088 52358
rect 55036 52294 55088 52300
rect 55048 52018 55076 52294
rect 53840 52012 53892 52018
rect 53840 51954 53892 51960
rect 55036 52012 55088 52018
rect 55036 51954 55088 51960
rect 53840 51808 53892 51814
rect 53840 51750 53892 51756
rect 53380 50924 53432 50930
rect 53380 50866 53432 50872
rect 53472 50856 53524 50862
rect 53472 50798 53524 50804
rect 53380 50448 53432 50454
rect 53380 50390 53432 50396
rect 52368 3188 52420 3194
rect 52368 3130 52420 3136
rect 53288 3188 53340 3194
rect 53288 3130 53340 3136
rect 52092 3120 52144 3126
rect 52092 3062 52144 3068
rect 52380 2446 52408 3130
rect 52828 2576 52880 2582
rect 52828 2518 52880 2524
rect 50620 2440 50672 2446
rect 50620 2382 50672 2388
rect 51264 2440 51316 2446
rect 51264 2382 51316 2388
rect 51816 2440 51868 2446
rect 51816 2382 51868 2388
rect 52368 2440 52420 2446
rect 52368 2382 52420 2388
rect 49884 2304 49936 2310
rect 49884 2246 49936 2252
rect 50620 2304 50672 2310
rect 50620 2246 50672 2252
rect 51356 2304 51408 2310
rect 51356 2246 51408 2252
rect 52092 2304 52144 2310
rect 52092 2246 52144 2252
rect 49896 800 49924 2246
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 800 50660 2246
rect 51368 800 51396 2246
rect 52104 800 52132 2246
rect 52840 800 52868 2518
rect 53300 2514 53328 3130
rect 53392 2961 53420 50390
rect 53484 50318 53512 50798
rect 53472 50312 53524 50318
rect 53472 50254 53524 50260
rect 53852 3738 53880 51750
rect 55048 51610 55076 51954
rect 55036 51604 55088 51610
rect 55036 51546 55088 51552
rect 55232 51074 55260 52838
rect 55232 51046 55444 51074
rect 53840 3732 53892 3738
rect 53840 3674 53892 3680
rect 53378 2952 53434 2961
rect 53378 2887 53434 2896
rect 53288 2508 53340 2514
rect 53288 2450 53340 2456
rect 53852 2446 53880 3674
rect 55416 3194 55444 51046
rect 56612 3194 56640 53926
rect 55404 3188 55456 3194
rect 55404 3130 55456 3136
rect 56600 3188 56652 3194
rect 56600 3130 56652 3136
rect 54300 2848 54352 2854
rect 54300 2790 54352 2796
rect 53840 2440 53892 2446
rect 53840 2382 53892 2388
rect 53564 2304 53616 2310
rect 53564 2246 53616 2252
rect 53576 800 53604 2246
rect 54312 800 54340 2790
rect 55416 2446 55444 3130
rect 56612 2446 56640 3130
rect 57072 3126 57100 55830
rect 57164 55350 57192 55898
rect 57152 55344 57204 55350
rect 57152 55286 57204 55292
rect 57716 55282 57744 56442
rect 57888 56432 57940 56438
rect 57888 56374 57940 56380
rect 57900 55758 57928 56374
rect 58440 55888 58492 55894
rect 58440 55830 58492 55836
rect 57888 55752 57940 55758
rect 57888 55694 57940 55700
rect 57796 55684 57848 55690
rect 57796 55626 57848 55632
rect 57808 55350 57836 55626
rect 57888 55616 57940 55622
rect 57888 55558 57940 55564
rect 57900 55418 57928 55558
rect 57888 55412 57940 55418
rect 57888 55354 57940 55360
rect 57796 55344 57848 55350
rect 57796 55286 57848 55292
rect 57704 55276 57756 55282
rect 57704 55218 57756 55224
rect 57152 55072 57204 55078
rect 57152 55014 57204 55020
rect 57164 3194 57192 55014
rect 58452 3194 58480 55830
rect 58992 55276 59044 55282
rect 58992 55218 59044 55224
rect 59004 3194 59032 55218
rect 59096 55214 59124 56850
rect 59464 56846 59492 57412
rect 59544 57394 59596 57400
rect 59648 57254 59676 57462
rect 59740 57458 59768 57870
rect 59820 57792 59872 57798
rect 59820 57734 59872 57740
rect 59728 57452 59780 57458
rect 59728 57394 59780 57400
rect 59636 57248 59688 57254
rect 59636 57190 59688 57196
rect 59740 56846 59768 57394
rect 59832 57066 59860 57734
rect 59832 57038 59952 57066
rect 59820 56976 59872 56982
rect 59820 56918 59872 56924
rect 59452 56840 59504 56846
rect 59452 56782 59504 56788
rect 59728 56840 59780 56846
rect 59728 56782 59780 56788
rect 59544 56772 59596 56778
rect 59544 56714 59596 56720
rect 59556 56506 59584 56714
rect 59544 56500 59596 56506
rect 59544 56442 59596 56448
rect 59740 56370 59768 56782
rect 59728 56364 59780 56370
rect 59728 56306 59780 56312
rect 59084 55208 59136 55214
rect 59084 55150 59136 55156
rect 59096 54874 59124 55150
rect 59084 54868 59136 54874
rect 59084 54810 59136 54816
rect 57152 3188 57204 3194
rect 57152 3130 57204 3136
rect 58440 3188 58492 3194
rect 58440 3130 58492 3136
rect 58992 3188 59044 3194
rect 58992 3130 59044 3136
rect 57060 3120 57112 3126
rect 57060 3062 57112 3068
rect 57164 2446 57192 3130
rect 57888 3120 57940 3126
rect 57888 3062 57940 3068
rect 57900 2446 57928 3062
rect 57980 2576 58032 2582
rect 57980 2518 58032 2524
rect 55404 2440 55456 2446
rect 55404 2382 55456 2388
rect 56600 2440 56652 2446
rect 56600 2382 56652 2388
rect 57152 2440 57204 2446
rect 57152 2382 57204 2388
rect 57888 2440 57940 2446
rect 57888 2382 57940 2388
rect 55036 2304 55088 2310
rect 55036 2246 55088 2252
rect 55772 2304 55824 2310
rect 55772 2246 55824 2252
rect 56508 2304 56560 2310
rect 56508 2246 56560 2252
rect 57244 2304 57296 2310
rect 57244 2246 57296 2252
rect 55048 800 55076 2246
rect 55784 800 55812 2246
rect 56520 800 56548 2246
rect 57256 800 57284 2246
rect 57992 800 58020 2518
rect 58452 2446 58480 3130
rect 59004 2446 59032 3130
rect 59832 2854 59860 56918
rect 59924 2990 59952 57038
rect 60016 56778 60044 60726
rect 62684 60314 62712 63718
rect 63144 61402 63172 66778
rect 65654 65852 65962 65861
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65787 65962 65796
rect 64512 65408 64564 65414
rect 64512 65350 64564 65356
rect 64420 62144 64472 62150
rect 64420 62086 64472 62092
rect 64052 61804 64104 61810
rect 64052 61746 64104 61752
rect 63132 61396 63184 61402
rect 63132 61338 63184 61344
rect 63224 61396 63276 61402
rect 63224 61338 63276 61344
rect 63040 60512 63092 60518
rect 63040 60454 63092 60460
rect 62672 60308 62724 60314
rect 62672 60250 62724 60256
rect 62120 59764 62172 59770
rect 62120 59706 62172 59712
rect 61844 59424 61896 59430
rect 61844 59366 61896 59372
rect 60280 59084 60332 59090
rect 60280 59026 60332 59032
rect 60292 58614 60320 59026
rect 61856 59022 61884 59366
rect 61660 59016 61712 59022
rect 61660 58958 61712 58964
rect 61844 59016 61896 59022
rect 61844 58958 61896 58964
rect 61292 58880 61344 58886
rect 61292 58822 61344 58828
rect 61304 58682 61332 58822
rect 61292 58676 61344 58682
rect 61292 58618 61344 58624
rect 60280 58608 60332 58614
rect 60280 58550 60332 58556
rect 60188 58540 60240 58546
rect 60188 58482 60240 58488
rect 60372 58540 60424 58546
rect 60372 58482 60424 58488
rect 60200 57866 60228 58482
rect 60384 57934 60412 58482
rect 61016 58404 61068 58410
rect 61016 58346 61068 58352
rect 60556 58336 60608 58342
rect 60556 58278 60608 58284
rect 60372 57928 60424 57934
rect 60372 57870 60424 57876
rect 60188 57860 60240 57866
rect 60188 57802 60240 57808
rect 60464 57860 60516 57866
rect 60464 57802 60516 57808
rect 60280 57248 60332 57254
rect 60280 57190 60332 57196
rect 60004 56772 60056 56778
rect 60004 56714 60056 56720
rect 60292 3194 60320 57190
rect 60476 56982 60504 57802
rect 60464 56976 60516 56982
rect 60464 56918 60516 56924
rect 60464 55752 60516 55758
rect 60464 55694 60516 55700
rect 60476 55282 60504 55694
rect 60464 55276 60516 55282
rect 60464 55218 60516 55224
rect 60476 24682 60504 55218
rect 60464 24676 60516 24682
rect 60464 24618 60516 24624
rect 60280 3188 60332 3194
rect 60280 3130 60332 3136
rect 60568 3126 60596 58278
rect 61028 58002 61056 58346
rect 61108 58336 61160 58342
rect 61108 58278 61160 58284
rect 61016 57996 61068 58002
rect 61016 57938 61068 57944
rect 61120 57934 61148 58278
rect 61304 58070 61332 58618
rect 61672 58546 61700 58958
rect 61936 58948 61988 58954
rect 61936 58890 61988 58896
rect 61948 58546 61976 58890
rect 62132 58614 62160 59706
rect 62488 59152 62540 59158
rect 62488 59094 62540 59100
rect 62212 59016 62264 59022
rect 62212 58958 62264 58964
rect 62120 58608 62172 58614
rect 62120 58550 62172 58556
rect 62224 58546 62252 58958
rect 61660 58540 61712 58546
rect 61660 58482 61712 58488
rect 61936 58540 61988 58546
rect 61936 58482 61988 58488
rect 62212 58540 62264 58546
rect 62212 58482 62264 58488
rect 61292 58064 61344 58070
rect 61292 58006 61344 58012
rect 61108 57928 61160 57934
rect 61108 57870 61160 57876
rect 61752 57928 61804 57934
rect 61752 57870 61804 57876
rect 61384 57860 61436 57866
rect 61384 57802 61436 57808
rect 60648 57792 60700 57798
rect 60648 57734 60700 57740
rect 60660 3194 60688 57734
rect 61396 57390 61424 57802
rect 61764 57458 61792 57870
rect 61948 57866 61976 58482
rect 62224 58138 62252 58482
rect 62396 58336 62448 58342
rect 62396 58278 62448 58284
rect 62212 58132 62264 58138
rect 62212 58074 62264 58080
rect 62120 57928 62172 57934
rect 62224 57916 62252 58074
rect 62172 57888 62252 57916
rect 62304 57928 62356 57934
rect 62120 57870 62172 57876
rect 62304 57870 62356 57876
rect 61936 57860 61988 57866
rect 61936 57802 61988 57808
rect 61752 57452 61804 57458
rect 61752 57394 61804 57400
rect 61384 57384 61436 57390
rect 61384 57326 61436 57332
rect 60832 57316 60884 57322
rect 60832 57258 60884 57264
rect 60740 56772 60792 56778
rect 60740 56714 60792 56720
rect 60752 56302 60780 56714
rect 60844 56710 60872 57258
rect 62132 56846 62160 57870
rect 62120 56840 62172 56846
rect 62120 56782 62172 56788
rect 60832 56704 60884 56710
rect 60832 56646 60884 56652
rect 60740 56296 60792 56302
rect 60740 56238 60792 56244
rect 60752 55894 60780 56238
rect 60844 56166 60872 56646
rect 61200 56296 61252 56302
rect 61200 56238 61252 56244
rect 60832 56160 60884 56166
rect 60832 56102 60884 56108
rect 60740 55888 60792 55894
rect 60740 55830 60792 55836
rect 60752 54670 60780 55830
rect 60844 54806 60872 56102
rect 61212 55282 61240 56238
rect 61200 55276 61252 55282
rect 61200 55218 61252 55224
rect 60832 54800 60884 54806
rect 60832 54742 60884 54748
rect 60740 54664 60792 54670
rect 60740 54606 60792 54612
rect 61212 24138 61240 55218
rect 61200 24132 61252 24138
rect 61200 24074 61252 24080
rect 60648 3188 60700 3194
rect 60648 3130 60700 3136
rect 60556 3120 60608 3126
rect 60556 3062 60608 3068
rect 59912 2984 59964 2990
rect 59912 2926 59964 2932
rect 59452 2848 59504 2854
rect 59452 2790 59504 2796
rect 59820 2848 59872 2854
rect 59820 2790 59872 2796
rect 58440 2440 58492 2446
rect 58440 2382 58492 2388
rect 58992 2440 59044 2446
rect 58992 2382 59044 2388
rect 58716 2304 58768 2310
rect 58716 2246 58768 2252
rect 58728 800 58756 2246
rect 59464 800 59492 2790
rect 60568 2514 60596 3062
rect 60556 2508 60608 2514
rect 60556 2450 60608 2456
rect 60660 2446 60688 3130
rect 61936 2984 61988 2990
rect 61936 2926 61988 2932
rect 61948 2446 61976 2926
rect 62316 2922 62344 57870
rect 62408 3126 62436 58278
rect 62396 3120 62448 3126
rect 62396 3062 62448 3068
rect 62500 2990 62528 59094
rect 62684 58954 62712 60250
rect 63052 58970 63080 60454
rect 63144 59634 63172 61338
rect 63236 59770 63264 61338
rect 63960 61192 64012 61198
rect 63774 61160 63830 61169
rect 63684 61124 63736 61130
rect 63960 61134 64012 61140
rect 63774 61095 63830 61104
rect 63684 61066 63736 61072
rect 63696 60722 63724 61066
rect 63788 61062 63816 61095
rect 63776 61056 63828 61062
rect 63776 60998 63828 61004
rect 63684 60716 63736 60722
rect 63684 60658 63736 60664
rect 63696 60110 63724 60658
rect 63972 60314 64000 61134
rect 64064 60858 64092 61746
rect 64328 61668 64380 61674
rect 64328 61610 64380 61616
rect 64052 60852 64104 60858
rect 64052 60794 64104 60800
rect 64340 60722 64368 61610
rect 64432 61198 64460 62086
rect 64524 61946 64552 65350
rect 65654 64764 65962 64773
rect 65654 64762 65660 64764
rect 65716 64762 65740 64764
rect 65796 64762 65820 64764
rect 65876 64762 65900 64764
rect 65956 64762 65962 64764
rect 65716 64710 65718 64762
rect 65898 64710 65900 64762
rect 65654 64708 65660 64710
rect 65716 64708 65740 64710
rect 65796 64708 65820 64710
rect 65876 64708 65900 64710
rect 65956 64708 65962 64710
rect 65654 64699 65962 64708
rect 65654 63676 65962 63685
rect 65654 63674 65660 63676
rect 65716 63674 65740 63676
rect 65796 63674 65820 63676
rect 65876 63674 65900 63676
rect 65956 63674 65962 63676
rect 65716 63622 65718 63674
rect 65898 63622 65900 63674
rect 65654 63620 65660 63622
rect 65716 63620 65740 63622
rect 65796 63620 65820 63622
rect 65876 63620 65900 63622
rect 65956 63620 65962 63622
rect 65654 63611 65962 63620
rect 65654 62588 65962 62597
rect 65654 62586 65660 62588
rect 65716 62586 65740 62588
rect 65796 62586 65820 62588
rect 65876 62586 65900 62588
rect 65956 62586 65962 62588
rect 65716 62534 65718 62586
rect 65898 62534 65900 62586
rect 65654 62532 65660 62534
rect 65716 62532 65740 62534
rect 65796 62532 65820 62534
rect 65876 62532 65900 62534
rect 65956 62532 65962 62534
rect 65654 62523 65962 62532
rect 65996 62490 66024 69498
rect 73356 69018 73384 70382
rect 74264 69760 74316 69766
rect 74264 69702 74316 69708
rect 73344 69012 73396 69018
rect 73344 68954 73396 68960
rect 73528 68672 73580 68678
rect 73528 68614 73580 68620
rect 66168 68128 66220 68134
rect 66168 68070 66220 68076
rect 66076 66292 66128 66298
rect 66076 66234 66128 66240
rect 65432 62484 65484 62490
rect 65432 62426 65484 62432
rect 65984 62484 66036 62490
rect 65984 62426 66036 62432
rect 64512 61940 64564 61946
rect 64512 61882 64564 61888
rect 64420 61192 64472 61198
rect 64420 61134 64472 61140
rect 64328 60716 64380 60722
rect 64328 60658 64380 60664
rect 63960 60308 64012 60314
rect 63960 60250 64012 60256
rect 64524 60110 64552 61882
rect 65340 61872 65392 61878
rect 65340 61814 65392 61820
rect 64972 61328 65024 61334
rect 64972 61270 65024 61276
rect 64604 60716 64656 60722
rect 64604 60658 64656 60664
rect 64788 60716 64840 60722
rect 64788 60658 64840 60664
rect 63592 60104 63644 60110
rect 63590 60072 63592 60081
rect 63684 60104 63736 60110
rect 63644 60072 63646 60081
rect 63684 60046 63736 60052
rect 64512 60104 64564 60110
rect 64512 60046 64564 60052
rect 63590 60007 63646 60016
rect 63224 59764 63276 59770
rect 63224 59706 63276 59712
rect 63132 59628 63184 59634
rect 63132 59570 63184 59576
rect 63696 59226 63724 60046
rect 64616 60042 64644 60658
rect 64800 60110 64828 60658
rect 64788 60104 64840 60110
rect 64788 60046 64840 60052
rect 64604 60036 64656 60042
rect 64604 59978 64656 59984
rect 63774 59936 63830 59945
rect 63774 59871 63830 59880
rect 63788 59634 63816 59871
rect 64616 59634 64644 59978
rect 64800 59945 64828 60046
rect 64786 59936 64842 59945
rect 64786 59871 64842 59880
rect 64800 59752 64828 59871
rect 64880 59764 64932 59770
rect 64800 59724 64880 59752
rect 64880 59706 64932 59712
rect 64696 59696 64748 59702
rect 64696 59638 64748 59644
rect 63776 59628 63828 59634
rect 63776 59570 63828 59576
rect 64420 59628 64472 59634
rect 64420 59570 64472 59576
rect 64604 59628 64656 59634
rect 64604 59570 64656 59576
rect 63684 59220 63736 59226
rect 63684 59162 63736 59168
rect 63132 59016 63184 59022
rect 63052 58964 63132 58970
rect 63052 58958 63184 58964
rect 62672 58948 62724 58954
rect 63052 58942 63172 58958
rect 62672 58890 62724 58896
rect 63040 57452 63092 57458
rect 63040 57394 63092 57400
rect 63052 57050 63080 57394
rect 63040 57044 63092 57050
rect 63040 56986 63092 56992
rect 63144 56302 63172 58942
rect 63788 58546 63816 59570
rect 64432 59498 64460 59570
rect 64616 59537 64644 59570
rect 64602 59528 64658 59537
rect 64420 59492 64472 59498
rect 64602 59463 64658 59472
rect 64420 59434 64472 59440
rect 63868 59424 63920 59430
rect 63868 59366 63920 59372
rect 63776 58540 63828 58546
rect 63776 58482 63828 58488
rect 63592 58336 63644 58342
rect 63592 58278 63644 58284
rect 63224 58132 63276 58138
rect 63224 58074 63276 58080
rect 63236 57934 63264 58074
rect 63604 58070 63632 58278
rect 63592 58064 63644 58070
rect 63592 58006 63644 58012
rect 63224 57928 63276 57934
rect 63592 57928 63644 57934
rect 63276 57888 63448 57916
rect 63224 57870 63276 57876
rect 63224 57792 63276 57798
rect 63224 57734 63276 57740
rect 63316 57792 63368 57798
rect 63316 57734 63368 57740
rect 63236 57458 63264 57734
rect 63224 57452 63276 57458
rect 63224 57394 63276 57400
rect 63132 56296 63184 56302
rect 63132 56238 63184 56244
rect 63328 3194 63356 57734
rect 63420 57458 63448 57888
rect 63592 57870 63644 57876
rect 63604 57798 63632 57870
rect 63592 57792 63644 57798
rect 63592 57734 63644 57740
rect 63408 57452 63460 57458
rect 63408 57394 63460 57400
rect 63880 3602 63908 59366
rect 64432 58682 64460 59434
rect 64616 59226 64644 59463
rect 64604 59220 64656 59226
rect 64604 59162 64656 59168
rect 64708 59158 64736 59638
rect 64696 59152 64748 59158
rect 64696 59094 64748 59100
rect 64420 58676 64472 58682
rect 64420 58618 64472 58624
rect 64880 58472 64932 58478
rect 64880 58414 64932 58420
rect 64328 57316 64380 57322
rect 64328 57258 64380 57264
rect 64340 3738 64368 57258
rect 64892 55758 64920 58414
rect 64880 55752 64932 55758
rect 64880 55694 64932 55700
rect 64328 3732 64380 3738
rect 64328 3674 64380 3680
rect 63868 3596 63920 3602
rect 63868 3538 63920 3544
rect 63316 3188 63368 3194
rect 63316 3130 63368 3136
rect 63408 3120 63460 3126
rect 63408 3062 63460 3068
rect 62488 2984 62540 2990
rect 62488 2926 62540 2932
rect 62304 2916 62356 2922
rect 62304 2858 62356 2864
rect 63040 2848 63092 2854
rect 63040 2790 63092 2796
rect 63052 2446 63080 2790
rect 63420 2446 63448 3062
rect 63868 2576 63920 2582
rect 63868 2518 63920 2524
rect 60648 2440 60700 2446
rect 60648 2382 60700 2388
rect 61936 2440 61988 2446
rect 61936 2382 61988 2388
rect 63040 2440 63092 2446
rect 63040 2382 63092 2388
rect 63408 2440 63460 2446
rect 63408 2382 63460 2388
rect 60188 2304 60240 2310
rect 60188 2246 60240 2252
rect 60924 2304 60976 2310
rect 60924 2246 60976 2252
rect 61660 2304 61712 2310
rect 61660 2246 61712 2252
rect 62396 2304 62448 2310
rect 62396 2246 62448 2252
rect 63408 2304 63460 2310
rect 63408 2246 63460 2252
rect 60200 800 60228 2246
rect 60936 800 60964 2246
rect 61672 800 61700 2246
rect 62408 800 62436 2246
rect 63144 870 63264 898
rect 63144 800 63172 870
rect 19812 734 20024 762
rect 20442 0 20498 800
rect 21178 0 21234 800
rect 21914 0 21970 800
rect 22650 0 22706 800
rect 23386 0 23442 800
rect 24122 0 24178 800
rect 24858 0 24914 800
rect 25594 0 25650 800
rect 26330 0 26386 800
rect 27066 0 27122 800
rect 27802 0 27858 800
rect 28538 0 28594 800
rect 29274 0 29330 800
rect 30010 0 30066 800
rect 30746 0 30802 800
rect 31482 0 31538 800
rect 32218 0 32274 800
rect 32954 0 33010 800
rect 33690 0 33746 800
rect 34426 0 34482 800
rect 35162 0 35218 800
rect 35898 0 35954 800
rect 36634 0 36690 800
rect 37370 0 37426 800
rect 38106 0 38162 800
rect 38842 0 38898 800
rect 39578 0 39634 800
rect 40314 0 40370 800
rect 41050 0 41106 800
rect 41786 0 41842 800
rect 42522 0 42578 800
rect 43258 0 43314 800
rect 43994 0 44050 800
rect 44730 0 44786 800
rect 45466 0 45522 800
rect 46202 0 46258 800
rect 46938 0 46994 800
rect 47674 0 47730 800
rect 48410 0 48466 800
rect 49146 0 49202 800
rect 49882 0 49938 800
rect 50618 0 50674 800
rect 51354 0 51410 800
rect 52090 0 52146 800
rect 52826 0 52882 800
rect 53562 0 53618 800
rect 54298 0 54354 800
rect 55034 0 55090 800
rect 55770 0 55826 800
rect 56506 0 56562 800
rect 57242 0 57298 800
rect 57978 0 58034 800
rect 58714 0 58770 800
rect 59450 0 59506 800
rect 60186 0 60242 800
rect 60922 0 60978 800
rect 61658 0 61714 800
rect 62394 0 62450 800
rect 63130 0 63186 800
rect 63236 762 63264 870
rect 63420 762 63448 2246
rect 63880 800 63908 2518
rect 64340 2446 64368 3674
rect 64984 3369 65012 61270
rect 65248 61192 65300 61198
rect 65248 61134 65300 61140
rect 65260 60722 65288 61134
rect 65248 60716 65300 60722
rect 65248 60658 65300 60664
rect 65352 60654 65380 61814
rect 65444 61130 65472 62426
rect 65524 61940 65576 61946
rect 65524 61882 65576 61888
rect 65536 61198 65564 61882
rect 66088 61878 66116 66234
rect 66180 61946 66208 68070
rect 66996 67856 67048 67862
rect 66996 67798 67048 67804
rect 66168 61940 66220 61946
rect 66168 61882 66220 61888
rect 66076 61872 66128 61878
rect 66076 61814 66128 61820
rect 66076 61600 66128 61606
rect 66076 61542 66128 61548
rect 65654 61500 65962 61509
rect 65654 61498 65660 61500
rect 65716 61498 65740 61500
rect 65796 61498 65820 61500
rect 65876 61498 65900 61500
rect 65956 61498 65962 61500
rect 65716 61446 65718 61498
rect 65898 61446 65900 61498
rect 65654 61444 65660 61446
rect 65716 61444 65740 61446
rect 65796 61444 65820 61446
rect 65876 61444 65900 61446
rect 65956 61444 65962 61446
rect 65654 61435 65962 61444
rect 65524 61192 65576 61198
rect 65524 61134 65576 61140
rect 65984 61192 66036 61198
rect 65984 61134 66036 61140
rect 65432 61124 65484 61130
rect 65432 61066 65484 61072
rect 65996 60722 66024 61134
rect 65432 60716 65484 60722
rect 65432 60658 65484 60664
rect 65984 60716 66036 60722
rect 65984 60658 66036 60664
rect 65340 60648 65392 60654
rect 65340 60590 65392 60596
rect 65156 60512 65208 60518
rect 65156 60454 65208 60460
rect 65064 60240 65116 60246
rect 65064 60182 65116 60188
rect 64970 3360 65026 3369
rect 64970 3295 65026 3304
rect 65076 3126 65104 60182
rect 65064 3120 65116 3126
rect 65064 3062 65116 3068
rect 65168 3058 65196 60454
rect 65248 60308 65300 60314
rect 65248 60250 65300 60256
rect 65260 59770 65288 60250
rect 65248 59764 65300 59770
rect 65248 59706 65300 59712
rect 65338 59664 65394 59673
rect 65338 59599 65394 59608
rect 65248 59560 65300 59566
rect 65248 59502 65300 59508
rect 65260 3194 65288 59502
rect 65352 59498 65380 59599
rect 65340 59492 65392 59498
rect 65340 59434 65392 59440
rect 65352 57934 65380 59434
rect 65444 59226 65472 60658
rect 65524 60648 65576 60654
rect 65524 60590 65576 60596
rect 65536 60518 65564 60590
rect 65524 60512 65576 60518
rect 65524 60454 65576 60460
rect 65536 60081 65564 60454
rect 65654 60412 65962 60421
rect 65654 60410 65660 60412
rect 65716 60410 65740 60412
rect 65796 60410 65820 60412
rect 65876 60410 65900 60412
rect 65956 60410 65962 60412
rect 65716 60358 65718 60410
rect 65898 60358 65900 60410
rect 65654 60356 65660 60358
rect 65716 60356 65740 60358
rect 65796 60356 65820 60358
rect 65876 60356 65900 60358
rect 65956 60356 65962 60358
rect 65654 60347 65962 60356
rect 65614 60208 65670 60217
rect 65614 60143 65670 60152
rect 65628 60110 65656 60143
rect 65996 60110 66024 60658
rect 66088 60518 66116 61542
rect 66168 61328 66220 61334
rect 66168 61270 66220 61276
rect 66076 60512 66128 60518
rect 66076 60454 66128 60460
rect 66076 60240 66128 60246
rect 66076 60182 66128 60188
rect 65616 60104 65668 60110
rect 65522 60072 65578 60081
rect 65616 60046 65668 60052
rect 65984 60104 66036 60110
rect 65984 60046 66036 60052
rect 65522 60007 65578 60016
rect 65708 60036 65760 60042
rect 65432 59220 65484 59226
rect 65432 59162 65484 59168
rect 65340 57928 65392 57934
rect 65340 57870 65392 57876
rect 65248 3188 65300 3194
rect 65248 3130 65300 3136
rect 65156 3052 65208 3058
rect 65156 2994 65208 3000
rect 65536 2990 65564 60007
rect 65708 59978 65760 59984
rect 65720 59650 65748 59978
rect 65720 59634 65840 59650
rect 65720 59628 65852 59634
rect 65720 59622 65800 59628
rect 65800 59570 65852 59576
rect 65706 59528 65762 59537
rect 65706 59463 65708 59472
rect 65760 59463 65762 59472
rect 65708 59434 65760 59440
rect 65984 59424 66036 59430
rect 65984 59366 66036 59372
rect 65654 59324 65962 59333
rect 65654 59322 65660 59324
rect 65716 59322 65740 59324
rect 65796 59322 65820 59324
rect 65876 59322 65900 59324
rect 65956 59322 65962 59324
rect 65716 59270 65718 59322
rect 65898 59270 65900 59322
rect 65654 59268 65660 59270
rect 65716 59268 65740 59270
rect 65796 59268 65820 59270
rect 65876 59268 65900 59270
rect 65956 59268 65962 59270
rect 65654 59259 65962 59268
rect 65616 59016 65668 59022
rect 65616 58958 65668 58964
rect 65628 58478 65656 58958
rect 65616 58472 65668 58478
rect 65616 58414 65668 58420
rect 65654 58236 65962 58245
rect 65654 58234 65660 58236
rect 65716 58234 65740 58236
rect 65796 58234 65820 58236
rect 65876 58234 65900 58236
rect 65956 58234 65962 58236
rect 65716 58182 65718 58234
rect 65898 58182 65900 58234
rect 65654 58180 65660 58182
rect 65716 58180 65740 58182
rect 65796 58180 65820 58182
rect 65876 58180 65900 58182
rect 65956 58180 65962 58182
rect 65654 58171 65962 58180
rect 65654 57148 65962 57157
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57083 65962 57092
rect 65654 56060 65962 56069
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55995 65962 56004
rect 65654 54972 65962 54981
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54907 65962 54916
rect 65654 53884 65962 53893
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53819 65962 53828
rect 65654 52796 65962 52805
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52731 65962 52740
rect 65654 51708 65962 51717
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51643 65962 51652
rect 65654 50620 65962 50629
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50555 65962 50564
rect 65654 49532 65962 49541
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49467 65962 49476
rect 65654 48444 65962 48453
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48379 65962 48388
rect 65654 47356 65962 47365
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47291 65962 47300
rect 65654 46268 65962 46277
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46203 65962 46212
rect 65654 45180 65962 45189
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45115 65962 45124
rect 65654 44092 65962 44101
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44027 65962 44036
rect 65654 43004 65962 43013
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42939 65962 42948
rect 65654 41916 65962 41925
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41851 65962 41860
rect 65654 40828 65962 40837
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40763 65962 40772
rect 65654 39740 65962 39749
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39675 65962 39684
rect 65654 38652 65962 38661
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38587 65962 38596
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 65996 3233 66024 59366
rect 65982 3224 66038 3233
rect 65982 3159 66038 3168
rect 65432 2984 65484 2990
rect 65432 2926 65484 2932
rect 65524 2984 65576 2990
rect 65524 2926 65576 2932
rect 64604 2848 64656 2854
rect 64604 2790 64656 2796
rect 64328 2440 64380 2446
rect 64328 2382 64380 2388
rect 64616 800 64644 2790
rect 65444 2446 65472 2926
rect 66088 2854 66116 60182
rect 66180 3466 66208 61270
rect 66720 61192 66772 61198
rect 66720 61134 66772 61140
rect 66732 60314 66760 61134
rect 66720 60308 66772 60314
rect 66720 60250 66772 60256
rect 67008 60042 67036 67798
rect 72332 67108 72384 67114
rect 72332 67050 72384 67056
rect 67364 60580 67416 60586
rect 67364 60522 67416 60528
rect 67376 60110 67404 60522
rect 68100 60240 68152 60246
rect 68098 60208 68100 60217
rect 68152 60208 68154 60217
rect 68098 60143 68154 60152
rect 67364 60104 67416 60110
rect 67364 60046 67416 60052
rect 66996 60036 67048 60042
rect 66996 59978 67048 59984
rect 67008 58682 67036 59978
rect 67180 59696 67232 59702
rect 67180 59638 67232 59644
rect 67192 59430 67220 59638
rect 67180 59424 67232 59430
rect 67180 59366 67232 59372
rect 67192 59158 67220 59366
rect 67180 59152 67232 59158
rect 67180 59094 67232 59100
rect 67376 58886 67404 60046
rect 72344 59566 72372 67050
rect 72424 65000 72476 65006
rect 72424 64942 72476 64948
rect 72436 59702 72464 64942
rect 72424 59696 72476 59702
rect 72424 59638 72476 59644
rect 72332 59560 72384 59566
rect 72332 59502 72384 59508
rect 67364 58880 67416 58886
rect 67364 58822 67416 58828
rect 66996 58676 67048 58682
rect 66996 58618 67048 58624
rect 66168 3460 66220 3466
rect 66168 3402 66220 3408
rect 66168 3188 66220 3194
rect 66168 3130 66220 3136
rect 66076 2848 66128 2854
rect 66076 2790 66128 2796
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 66180 2514 66208 3130
rect 66352 2916 66404 2922
rect 66352 2858 66404 2864
rect 66168 2508 66220 2514
rect 66168 2450 66220 2456
rect 66364 2446 66392 2858
rect 65432 2440 65484 2446
rect 65432 2382 65484 2388
rect 66352 2440 66404 2446
rect 66352 2382 66404 2388
rect 67376 2378 67404 58822
rect 69664 47456 69716 47462
rect 69664 47398 69716 47404
rect 69676 46986 69704 47398
rect 69664 46980 69716 46986
rect 69664 46922 69716 46928
rect 69664 46368 69716 46374
rect 69664 46310 69716 46316
rect 69676 45830 69704 46310
rect 69664 45824 69716 45830
rect 69664 45766 69716 45772
rect 69664 45280 69716 45286
rect 69664 45222 69716 45228
rect 69676 44742 69704 45222
rect 69664 44736 69716 44742
rect 69664 44678 69716 44684
rect 69664 42016 69716 42022
rect 69664 41958 69716 41964
rect 69676 41478 69704 41958
rect 69664 41472 69716 41478
rect 69664 41414 69716 41420
rect 69664 39840 69716 39846
rect 69664 39782 69716 39788
rect 69676 39302 69704 39782
rect 69664 39296 69716 39302
rect 69664 39238 69716 39244
rect 69664 37664 69716 37670
rect 69664 37606 69716 37612
rect 69676 37330 69704 37606
rect 69664 37324 69716 37330
rect 69664 37266 69716 37272
rect 69664 36576 69716 36582
rect 69664 36518 69716 36524
rect 69676 36038 69704 36518
rect 69664 36032 69716 36038
rect 69664 35974 69716 35980
rect 68008 35488 68060 35494
rect 68008 35430 68060 35436
rect 68020 34950 68048 35430
rect 68008 34944 68060 34950
rect 68008 34886 68060 34892
rect 69664 32224 69716 32230
rect 69664 32166 69716 32172
rect 69676 31890 69704 32166
rect 69664 31884 69716 31890
rect 69664 31826 69716 31832
rect 68008 31136 68060 31142
rect 68008 31078 68060 31084
rect 68020 30598 68048 31078
rect 68008 30592 68060 30598
rect 68008 30534 68060 30540
rect 69664 30048 69716 30054
rect 69664 29990 69716 29996
rect 69676 29510 69704 29990
rect 69664 29504 69716 29510
rect 69664 29446 69716 29452
rect 69664 26784 69716 26790
rect 69664 26726 69716 26732
rect 69676 26314 69704 26726
rect 69664 26308 69716 26314
rect 69664 26250 69716 26256
rect 69664 25764 69716 25770
rect 69664 25706 69716 25712
rect 69676 25158 69704 25706
rect 69664 25152 69716 25158
rect 69664 25094 69716 25100
rect 69664 24608 69716 24614
rect 69664 24550 69716 24556
rect 69676 24070 69704 24550
rect 69664 24064 69716 24070
rect 69664 24006 69716 24012
rect 68008 20256 68060 20262
rect 68008 20198 68060 20204
rect 68020 19718 68048 20198
rect 68008 19712 68060 19718
rect 68008 19654 68060 19660
rect 68008 14816 68060 14822
rect 68008 14758 68060 14764
rect 68020 14278 68048 14758
rect 68008 14272 68060 14278
rect 68008 14214 68060 14220
rect 69664 9376 69716 9382
rect 69664 9318 69716 9324
rect 69676 8838 69704 9318
rect 69664 8832 69716 8838
rect 69664 8774 69716 8780
rect 69664 5024 69716 5030
rect 69664 4966 69716 4972
rect 69676 4486 69704 4966
rect 69664 4480 69716 4486
rect 69664 4422 69716 4428
rect 69664 3596 69716 3602
rect 69664 3538 69716 3544
rect 69294 3224 69350 3233
rect 69294 3159 69296 3168
rect 69348 3159 69350 3168
rect 69296 3130 69348 3136
rect 68192 3120 68244 3126
rect 68192 3062 68244 3068
rect 68204 2446 68232 3062
rect 68928 3052 68980 3058
rect 68928 2994 68980 3000
rect 68940 2446 68968 2994
rect 69020 2576 69072 2582
rect 69020 2518 69072 2524
rect 68192 2440 68244 2446
rect 68192 2382 68244 2388
rect 68928 2440 68980 2446
rect 68928 2382 68980 2388
rect 67364 2372 67416 2378
rect 67364 2314 67416 2320
rect 65340 2304 65392 2310
rect 65340 2246 65392 2252
rect 66076 2304 66128 2310
rect 66076 2246 66128 2252
rect 66812 2304 66864 2310
rect 66812 2246 66864 2252
rect 67548 2304 67600 2310
rect 67548 2246 67600 2252
rect 68560 2304 68612 2310
rect 68560 2246 68612 2252
rect 65352 800 65380 2246
rect 66088 800 66116 2246
rect 66824 800 66852 2246
rect 67560 800 67588 2246
rect 68296 870 68416 898
rect 68296 800 68324 870
rect 63236 734 63448 762
rect 63866 0 63922 800
rect 64602 0 64658 800
rect 65338 0 65394 800
rect 66074 0 66130 800
rect 66810 0 66866 800
rect 67546 0 67602 800
rect 68282 0 68338 800
rect 68388 762 68416 870
rect 68572 762 68600 2246
rect 69032 800 69060 2518
rect 69676 2446 69704 3538
rect 70584 3460 70636 3466
rect 70584 3402 70636 3408
rect 70596 3194 70624 3402
rect 72054 3360 72110 3369
rect 72054 3295 72110 3304
rect 72068 3194 72096 3295
rect 70584 3188 70636 3194
rect 70584 3130 70636 3136
rect 72056 3188 72108 3194
rect 72056 3130 72108 3136
rect 69756 2848 69808 2854
rect 69756 2790 69808 2796
rect 69664 2440 69716 2446
rect 69664 2382 69716 2388
rect 69768 800 69796 2790
rect 70596 2446 70624 3130
rect 71504 2916 71556 2922
rect 71504 2858 71556 2864
rect 71516 2446 71544 2858
rect 72068 2446 72096 3130
rect 73344 2848 73396 2854
rect 73344 2790 73396 2796
rect 73356 2446 73384 2790
rect 73540 2650 73568 68614
rect 73896 2848 73948 2854
rect 73896 2790 73948 2796
rect 73528 2644 73580 2650
rect 73528 2586 73580 2592
rect 73908 2446 73936 2790
rect 74276 2650 74304 69702
rect 74724 3392 74776 3398
rect 74724 3334 74776 3340
rect 74264 2644 74316 2650
rect 74264 2586 74316 2592
rect 74736 2446 74764 3334
rect 74908 3052 74960 3058
rect 74908 2994 74960 3000
rect 70584 2440 70636 2446
rect 70584 2382 70636 2388
rect 71504 2440 71556 2446
rect 71504 2382 71556 2388
rect 72056 2440 72108 2446
rect 72056 2382 72108 2388
rect 72700 2440 72752 2446
rect 72700 2382 72752 2388
rect 73344 2440 73396 2446
rect 73344 2382 73396 2388
rect 73436 2440 73488 2446
rect 73436 2382 73488 2388
rect 73896 2440 73948 2446
rect 74724 2440 74776 2446
rect 73896 2382 73948 2388
rect 74460 2400 74724 2428
rect 70492 2304 70544 2310
rect 70492 2246 70544 2252
rect 71228 2304 71280 2310
rect 71228 2246 71280 2252
rect 71964 2304 72016 2310
rect 71964 2246 72016 2252
rect 70504 800 70532 2246
rect 71240 800 71268 2246
rect 71976 800 72004 2246
rect 72712 800 72740 2382
rect 73448 800 73476 2382
rect 74184 870 74304 898
rect 74184 800 74212 870
rect 68388 734 68600 762
rect 69018 0 69074 800
rect 69754 0 69810 800
rect 70490 0 70546 800
rect 71226 0 71282 800
rect 71962 0 72018 800
rect 72698 0 72754 800
rect 73434 0 73490 800
rect 74170 0 74226 800
rect 74276 762 74304 870
rect 74460 762 74488 2400
rect 74724 2382 74776 2388
rect 74920 800 74948 2994
rect 75012 2650 75040 70450
rect 75840 70106 75868 70858
rect 75932 70650 75960 72014
rect 76116 71194 76144 72626
rect 76208 71738 76236 73102
rect 76196 71732 76248 71738
rect 76196 71674 76248 71680
rect 76288 71596 76340 71602
rect 76288 71538 76340 71544
rect 76300 71398 76328 71538
rect 76288 71392 76340 71398
rect 76288 71334 76340 71340
rect 76104 71188 76156 71194
rect 76104 71130 76156 71136
rect 76012 70984 76064 70990
rect 76012 70926 76064 70932
rect 75920 70644 75972 70650
rect 75920 70586 75972 70592
rect 76024 70530 76052 70926
rect 75932 70502 76052 70530
rect 75828 70100 75880 70106
rect 75828 70042 75880 70048
rect 75184 68128 75236 68134
rect 75184 68070 75236 68076
rect 75196 61198 75224 68070
rect 75184 61192 75236 61198
rect 75184 61134 75236 61140
rect 75932 3194 75960 70502
rect 76012 65408 76064 65414
rect 76012 65350 76064 65356
rect 76024 60042 76052 65350
rect 76012 60036 76064 60042
rect 76012 59978 76064 59984
rect 76196 56704 76248 56710
rect 76196 56646 76248 56652
rect 76208 56370 76236 56646
rect 76196 56364 76248 56370
rect 76196 56306 76248 56312
rect 76196 54528 76248 54534
rect 76196 54470 76248 54476
rect 76208 53990 76236 54470
rect 76196 53984 76248 53990
rect 76196 53926 76248 53932
rect 76012 7200 76064 7206
rect 76012 7142 76064 7148
rect 76024 6662 76052 7142
rect 76012 6656 76064 6662
rect 76012 6598 76064 6604
rect 75920 3188 75972 3194
rect 75920 3130 75972 3136
rect 75736 2848 75788 2854
rect 75736 2790 75788 2796
rect 75000 2644 75052 2650
rect 75000 2586 75052 2592
rect 75748 2428 75776 2790
rect 76300 2650 76328 71334
rect 76576 60654 76604 75142
rect 78048 75041 78076 75142
rect 78034 75032 78090 75041
rect 78034 74967 78090 74976
rect 78128 74860 78180 74866
rect 78128 74802 78180 74808
rect 77576 74724 77628 74730
rect 77576 74666 77628 74672
rect 77024 73568 77076 73574
rect 77024 73510 77076 73516
rect 76656 69216 76708 69222
rect 76656 69158 76708 69164
rect 76564 60648 76616 60654
rect 76564 60590 76616 60596
rect 76668 60314 76696 69158
rect 77036 61130 77064 73510
rect 77484 64320 77536 64326
rect 77484 64262 77536 64268
rect 77300 62688 77352 62694
rect 77300 62630 77352 62636
rect 77024 61124 77076 61130
rect 77024 61066 77076 61072
rect 76656 60308 76708 60314
rect 76656 60250 76708 60256
rect 77312 57866 77340 62630
rect 77392 62144 77444 62150
rect 77392 62086 77444 62092
rect 77300 57860 77352 57866
rect 77300 57802 77352 57808
rect 77404 57322 77432 62086
rect 77496 57798 77524 64262
rect 77484 57792 77536 57798
rect 77484 57734 77536 57740
rect 77392 57316 77444 57322
rect 77392 57258 77444 57264
rect 77588 55214 77616 74666
rect 78140 74390 78168 74802
rect 78128 74384 78180 74390
rect 78126 74352 78128 74361
rect 78180 74352 78182 74361
rect 78126 74287 78182 74296
rect 78140 74261 78168 74287
rect 77850 73672 77906 73681
rect 77850 73607 77852 73616
rect 77904 73607 77906 73616
rect 77852 73578 77904 73584
rect 78036 73024 78088 73030
rect 78034 72992 78036 73001
rect 78088 72992 78090 73001
rect 78034 72927 78090 72936
rect 77852 72480 77904 72486
rect 77852 72422 77904 72428
rect 77864 72321 77892 72422
rect 77850 72312 77906 72321
rect 77850 72247 77906 72256
rect 78036 71936 78088 71942
rect 78036 71878 78088 71884
rect 78048 71641 78076 71878
rect 78034 71632 78090 71641
rect 78034 71567 78090 71576
rect 78034 70952 78090 70961
rect 78034 70887 78090 70896
rect 78048 70854 78076 70887
rect 78036 70848 78088 70854
rect 78036 70790 78088 70796
rect 77852 70304 77904 70310
rect 77850 70272 77852 70281
rect 77904 70272 77906 70281
rect 77850 70207 77906 70216
rect 78128 69896 78180 69902
rect 78128 69838 78180 69844
rect 77944 69760 77996 69766
rect 77944 69702 77996 69708
rect 77956 69562 77984 69702
rect 78140 69601 78168 69838
rect 78126 69592 78182 69601
rect 77944 69556 77996 69562
rect 78126 69527 78182 69536
rect 77944 69498 77996 69504
rect 77944 69420 77996 69426
rect 77944 69362 77996 69368
rect 77956 68921 77984 69362
rect 77942 68912 77998 68921
rect 77942 68847 77998 68856
rect 77944 68672 77996 68678
rect 77944 68614 77996 68620
rect 77956 68338 77984 68614
rect 77944 68332 77996 68338
rect 77944 68274 77996 68280
rect 77956 68241 77984 68274
rect 77942 68232 77998 68241
rect 77942 68167 77998 68176
rect 78128 67720 78180 67726
rect 78128 67662 78180 67668
rect 78140 67561 78168 67662
rect 78126 67552 78182 67561
rect 78126 67487 78182 67496
rect 77944 67244 77996 67250
rect 77944 67186 77996 67192
rect 77956 66881 77984 67186
rect 77942 66872 77998 66881
rect 77942 66807 77998 66816
rect 78128 66632 78180 66638
rect 78128 66574 78180 66580
rect 77944 66496 77996 66502
rect 77944 66438 77996 66444
rect 77956 66298 77984 66438
rect 77944 66292 77996 66298
rect 77944 66234 77996 66240
rect 78140 66201 78168 66574
rect 78126 66192 78182 66201
rect 78126 66127 78182 66136
rect 78128 65544 78180 65550
rect 78126 65512 78128 65521
rect 78180 65512 78182 65521
rect 78126 65447 78182 65456
rect 77944 65068 77996 65074
rect 77944 65010 77996 65016
rect 77956 64841 77984 65010
rect 77942 64832 77998 64841
rect 77942 64767 77998 64776
rect 78128 64456 78180 64462
rect 78128 64398 78180 64404
rect 78140 64161 78168 64398
rect 78126 64152 78182 64161
rect 78126 64087 78182 64096
rect 77944 63980 77996 63986
rect 77944 63922 77996 63928
rect 77956 63481 77984 63922
rect 77942 63472 77998 63481
rect 77942 63407 77998 63416
rect 77944 63232 77996 63238
rect 77944 63174 77996 63180
rect 77956 62898 77984 63174
rect 77944 62892 77996 62898
rect 77944 62834 77996 62840
rect 77956 62801 77984 62834
rect 77942 62792 77998 62801
rect 77942 62727 77998 62736
rect 78128 62280 78180 62286
rect 78128 62222 78180 62228
rect 78140 62121 78168 62222
rect 78126 62112 78182 62121
rect 78126 62047 78182 62056
rect 77944 61804 77996 61810
rect 77944 61746 77996 61752
rect 77760 61600 77812 61606
rect 77760 61542 77812 61548
rect 77772 61266 77800 61542
rect 77956 61441 77984 61746
rect 77942 61432 77998 61441
rect 77942 61367 77998 61376
rect 77760 61260 77812 61266
rect 77760 61202 77812 61208
rect 78128 61192 78180 61198
rect 78128 61134 78180 61140
rect 77944 61056 77996 61062
rect 77944 60998 77996 61004
rect 77956 60790 77984 60998
rect 77944 60784 77996 60790
rect 78140 60761 78168 61134
rect 77944 60726 77996 60732
rect 78126 60752 78182 60761
rect 78126 60687 78182 60696
rect 78128 60104 78180 60110
rect 78126 60072 78128 60081
rect 78180 60072 78182 60081
rect 78126 60007 78182 60016
rect 77944 59968 77996 59974
rect 77944 59910 77996 59916
rect 77956 59770 77984 59910
rect 77944 59764 77996 59770
rect 77944 59706 77996 59712
rect 77944 59628 77996 59634
rect 77944 59570 77996 59576
rect 77760 59424 77812 59430
rect 77956 59401 77984 59570
rect 77760 59366 77812 59372
rect 77942 59392 77998 59401
rect 77772 58954 77800 59366
rect 77942 59327 77998 59336
rect 78128 59016 78180 59022
rect 78128 58958 78180 58964
rect 77760 58948 77812 58954
rect 77760 58890 77812 58896
rect 77944 58880 77996 58886
rect 77944 58822 77996 58828
rect 77956 58682 77984 58822
rect 78140 58721 78168 58958
rect 78126 58712 78182 58721
rect 77944 58676 77996 58682
rect 78126 58647 78182 58656
rect 77944 58618 77996 58624
rect 77944 58540 77996 58546
rect 77944 58482 77996 58488
rect 77760 58336 77812 58342
rect 77760 58278 77812 58284
rect 77772 57526 77800 58278
rect 77956 58041 77984 58482
rect 77942 58032 77998 58041
rect 77942 57967 77998 57976
rect 77944 57792 77996 57798
rect 77944 57734 77996 57740
rect 77760 57520 77812 57526
rect 77760 57462 77812 57468
rect 77956 57458 77984 57734
rect 77944 57452 77996 57458
rect 77944 57394 77996 57400
rect 77956 57361 77984 57394
rect 77942 57352 77998 57361
rect 77942 57287 77998 57296
rect 77760 57248 77812 57254
rect 77760 57190 77812 57196
rect 77772 57050 77800 57190
rect 77760 57044 77812 57050
rect 77760 56986 77812 56992
rect 78128 56840 78180 56846
rect 78128 56782 78180 56788
rect 78140 56681 78168 56782
rect 78126 56672 78182 56681
rect 78126 56607 78182 56616
rect 77944 56364 77996 56370
rect 77944 56306 77996 56312
rect 77956 56001 77984 56306
rect 77942 55992 77998 56001
rect 77942 55927 77998 55936
rect 78128 55752 78180 55758
rect 78128 55694 78180 55700
rect 78140 55321 78168 55694
rect 78126 55312 78182 55321
rect 78126 55247 78182 55256
rect 77588 55186 77800 55214
rect 77484 54120 77536 54126
rect 77484 54062 77536 54068
rect 77300 53576 77352 53582
rect 77300 53518 77352 53524
rect 77392 53576 77444 53582
rect 77392 53518 77444 53524
rect 77312 53281 77340 53518
rect 77298 53272 77354 53281
rect 77298 53207 77354 53216
rect 77404 52562 77432 53518
rect 77496 52902 77524 54062
rect 77668 53508 77720 53514
rect 77668 53450 77720 53456
rect 77680 53106 77708 53450
rect 77668 53100 77720 53106
rect 77668 53042 77720 53048
rect 77576 53032 77628 53038
rect 77576 52974 77628 52980
rect 77484 52896 77536 52902
rect 77484 52838 77536 52844
rect 77588 52630 77616 52974
rect 77576 52624 77628 52630
rect 77574 52592 77576 52601
rect 77628 52592 77630 52601
rect 77392 52556 77444 52562
rect 77574 52527 77630 52536
rect 77392 52498 77444 52504
rect 77300 51400 77352 51406
rect 77300 51342 77352 51348
rect 77312 51241 77340 51342
rect 77298 51232 77354 51241
rect 77298 51167 77354 51176
rect 77116 50856 77168 50862
rect 77116 50798 77168 50804
rect 77208 50856 77260 50862
rect 77208 50798 77260 50804
rect 77128 50561 77156 50798
rect 77114 50552 77170 50561
rect 77114 50487 77170 50496
rect 77220 50250 77248 50798
rect 77392 50312 77444 50318
rect 77392 50254 77444 50260
rect 77576 50312 77628 50318
rect 77576 50254 77628 50260
rect 77208 50244 77260 50250
rect 77208 50186 77260 50192
rect 77404 49910 77432 50254
rect 77392 49904 77444 49910
rect 77390 49872 77392 49881
rect 77444 49872 77446 49881
rect 77390 49807 77446 49816
rect 77588 49774 77616 50254
rect 77772 50182 77800 55186
rect 78128 55072 78180 55078
rect 78128 55014 78180 55020
rect 78140 54670 78168 55014
rect 77944 54664 77996 54670
rect 78128 54664 78180 54670
rect 77944 54606 77996 54612
rect 78126 54632 78128 54641
rect 78180 54632 78182 54641
rect 77956 54126 77984 54606
rect 78126 54567 78182 54576
rect 77944 54120 77996 54126
rect 77944 54062 77996 54068
rect 77956 53961 77984 54062
rect 77942 53952 77998 53961
rect 77942 53887 77998 53896
rect 77944 52352 77996 52358
rect 77944 52294 77996 52300
rect 77956 51950 77984 52294
rect 77944 51944 77996 51950
rect 77942 51912 77944 51921
rect 77996 51912 77998 51921
rect 77942 51847 77998 51856
rect 77760 50176 77812 50182
rect 77760 50118 77812 50124
rect 77576 49768 77628 49774
rect 77576 49710 77628 49716
rect 78128 49632 78180 49638
rect 78128 49574 78180 49580
rect 78140 49230 78168 49574
rect 78128 49224 78180 49230
rect 78126 49192 78128 49201
rect 78180 49192 78182 49201
rect 78126 49127 78182 49136
rect 77116 48680 77168 48686
rect 77116 48622 77168 48628
rect 77128 48521 77156 48622
rect 77114 48512 77170 48521
rect 77114 48447 77170 48456
rect 77024 48000 77076 48006
rect 77024 47942 77076 47948
rect 78036 48000 78088 48006
rect 78036 47942 78088 47948
rect 77036 47530 77064 47942
rect 78048 47841 78076 47942
rect 78034 47832 78090 47841
rect 78034 47767 78090 47776
rect 77024 47524 77076 47530
rect 77024 47466 77076 47472
rect 77852 47456 77904 47462
rect 77852 47398 77904 47404
rect 77864 47161 77892 47398
rect 77850 47152 77906 47161
rect 77850 47087 77906 47096
rect 77850 46472 77906 46481
rect 77850 46407 77852 46416
rect 77904 46407 77906 46416
rect 77852 46378 77904 46384
rect 78036 45824 78088 45830
rect 78034 45792 78036 45801
rect 78088 45792 78090 45801
rect 78034 45727 78090 45736
rect 77852 45280 77904 45286
rect 77852 45222 77904 45228
rect 77864 45121 77892 45222
rect 77850 45112 77906 45121
rect 77850 45047 77906 45056
rect 77300 44736 77352 44742
rect 77300 44678 77352 44684
rect 78036 44736 78088 44742
rect 78036 44678 78088 44684
rect 77312 44198 77340 44678
rect 78048 44441 78076 44678
rect 78034 44432 78090 44441
rect 78034 44367 78090 44376
rect 77300 44192 77352 44198
rect 77300 44134 77352 44140
rect 78034 43752 78090 43761
rect 78034 43687 78090 43696
rect 78048 43654 78076 43687
rect 77300 43648 77352 43654
rect 77300 43590 77352 43596
rect 78036 43648 78088 43654
rect 78036 43590 78088 43596
rect 77312 43178 77340 43590
rect 77300 43172 77352 43178
rect 77300 43114 77352 43120
rect 76932 43104 76984 43110
rect 77852 43104 77904 43110
rect 76932 43046 76984 43052
rect 77850 43072 77852 43081
rect 77904 43072 77906 43081
rect 76944 42566 76972 43046
rect 77850 43007 77906 43016
rect 76932 42560 76984 42566
rect 76932 42502 76984 42508
rect 77024 42560 77076 42566
rect 77024 42502 77076 42508
rect 78036 42560 78088 42566
rect 78036 42502 78088 42508
rect 77036 42090 77064 42502
rect 78048 42401 78076 42502
rect 78034 42392 78090 42401
rect 78034 42327 78090 42336
rect 77024 42084 77076 42090
rect 77024 42026 77076 42032
rect 77852 42016 77904 42022
rect 77852 41958 77904 41964
rect 77864 41721 77892 41958
rect 77850 41712 77906 41721
rect 77850 41647 77906 41656
rect 77850 41032 77906 41041
rect 77850 40967 77852 40976
rect 77904 40967 77906 40976
rect 77852 40938 77904 40944
rect 77116 40928 77168 40934
rect 77116 40870 77168 40876
rect 77128 40458 77156 40870
rect 77116 40452 77168 40458
rect 77116 40394 77168 40400
rect 78036 40384 78088 40390
rect 78034 40352 78036 40361
rect 78088 40352 78090 40361
rect 78034 40287 78090 40296
rect 77852 39840 77904 39846
rect 77852 39782 77904 39788
rect 77864 39681 77892 39782
rect 77850 39672 77906 39681
rect 77850 39607 77906 39616
rect 77300 39296 77352 39302
rect 77300 39238 77352 39244
rect 78036 39296 78088 39302
rect 78036 39238 78088 39244
rect 77312 38758 77340 39238
rect 78048 39001 78076 39238
rect 78034 38992 78090 39001
rect 78034 38927 78090 38936
rect 77300 38752 77352 38758
rect 77300 38694 77352 38700
rect 78034 38312 78090 38321
rect 78034 38247 78090 38256
rect 78048 38214 78076 38247
rect 77024 38208 77076 38214
rect 77024 38150 77076 38156
rect 78036 38208 78088 38214
rect 78036 38150 78088 38156
rect 77036 37738 77064 38150
rect 77024 37732 77076 37738
rect 77024 37674 77076 37680
rect 77852 37664 77904 37670
rect 77850 37632 77852 37641
rect 77904 37632 77906 37641
rect 77850 37567 77906 37576
rect 77300 37120 77352 37126
rect 77300 37062 77352 37068
rect 78036 37120 78088 37126
rect 78036 37062 78088 37068
rect 77312 36854 77340 37062
rect 78048 36961 78076 37062
rect 78034 36952 78090 36961
rect 78034 36887 78090 36896
rect 77300 36848 77352 36854
rect 77300 36790 77352 36796
rect 77852 36576 77904 36582
rect 77852 36518 77904 36524
rect 77864 36281 77892 36518
rect 77850 36272 77906 36281
rect 77850 36207 77906 36216
rect 77850 35592 77906 35601
rect 77850 35527 77852 35536
rect 77904 35527 77906 35536
rect 77852 35498 77904 35504
rect 77300 34944 77352 34950
rect 78036 34944 78088 34950
rect 77300 34886 77352 34892
rect 78034 34912 78036 34921
rect 78088 34912 78090 34921
rect 77312 34678 77340 34886
rect 78034 34847 78090 34856
rect 77300 34672 77352 34678
rect 77300 34614 77352 34620
rect 77116 34536 77168 34542
rect 77116 34478 77168 34484
rect 77128 33862 77156 34478
rect 77852 34400 77904 34406
rect 77852 34342 77904 34348
rect 77864 34241 77892 34342
rect 77850 34232 77906 34241
rect 77850 34167 77906 34176
rect 77116 33856 77168 33862
rect 77116 33798 77168 33804
rect 77300 33856 77352 33862
rect 77300 33798 77352 33804
rect 78036 33856 78088 33862
rect 78036 33798 78088 33804
rect 77312 33318 77340 33798
rect 78048 33561 78076 33798
rect 78034 33552 78090 33561
rect 78034 33487 78090 33496
rect 77300 33312 77352 33318
rect 77300 33254 77352 33260
rect 78034 32872 78090 32881
rect 78034 32807 78090 32816
rect 78048 32774 78076 32807
rect 77024 32768 77076 32774
rect 77024 32710 77076 32716
rect 78036 32768 78088 32774
rect 78036 32710 78088 32716
rect 77036 32298 77064 32710
rect 77024 32292 77076 32298
rect 77024 32234 77076 32240
rect 77852 32224 77904 32230
rect 77850 32192 77852 32201
rect 77904 32192 77906 32201
rect 77850 32127 77906 32136
rect 78036 31952 78088 31958
rect 78036 31894 78088 31900
rect 78048 31521 78076 31894
rect 78034 31512 78090 31521
rect 78034 31447 78090 31456
rect 77852 31136 77904 31142
rect 77852 31078 77904 31084
rect 77864 30841 77892 31078
rect 77850 30832 77906 30841
rect 77850 30767 77906 30776
rect 77850 30152 77906 30161
rect 77850 30087 77852 30096
rect 77904 30087 77906 30096
rect 77852 30058 77904 30064
rect 77300 29504 77352 29510
rect 78036 29504 78088 29510
rect 77300 29446 77352 29452
rect 78034 29472 78036 29481
rect 78088 29472 78090 29481
rect 77312 29170 77340 29446
rect 78034 29407 78090 29416
rect 77300 29164 77352 29170
rect 77300 29106 77352 29112
rect 77116 29028 77168 29034
rect 77116 28970 77168 28976
rect 77852 29028 77904 29034
rect 77852 28970 77904 28976
rect 77128 28422 77156 28970
rect 77864 28801 77892 28970
rect 77850 28792 77906 28801
rect 77850 28727 77906 28736
rect 77116 28416 77168 28422
rect 77116 28358 77168 28364
rect 77300 28416 77352 28422
rect 77300 28358 77352 28364
rect 78036 28416 78088 28422
rect 78036 28358 78088 28364
rect 77312 27878 77340 28358
rect 78048 28121 78076 28358
rect 78034 28112 78090 28121
rect 78034 28047 78090 28056
rect 77300 27872 77352 27878
rect 77300 27814 77352 27820
rect 78034 27432 78090 27441
rect 78034 27367 78090 27376
rect 78048 27334 78076 27367
rect 77024 27328 77076 27334
rect 77024 27270 77076 27276
rect 78036 27328 78088 27334
rect 78036 27270 78088 27276
rect 77036 26858 77064 27270
rect 77024 26852 77076 26858
rect 77024 26794 77076 26800
rect 77852 26784 77904 26790
rect 77850 26752 77852 26761
rect 77904 26752 77906 26761
rect 77850 26687 77906 26696
rect 78036 26512 78088 26518
rect 78036 26454 78088 26460
rect 77392 26376 77444 26382
rect 77392 26318 77444 26324
rect 77404 25702 77432 26318
rect 78048 26081 78076 26454
rect 78034 26072 78090 26081
rect 78034 26007 78090 26016
rect 77392 25696 77444 25702
rect 77392 25638 77444 25644
rect 77852 25696 77904 25702
rect 77852 25638 77904 25644
rect 77864 25401 77892 25638
rect 77850 25392 77906 25401
rect 77850 25327 77906 25336
rect 77850 24712 77906 24721
rect 77850 24647 77852 24656
rect 77904 24647 77906 24656
rect 77852 24618 77904 24624
rect 77300 24064 77352 24070
rect 78036 24064 78088 24070
rect 77300 24006 77352 24012
rect 78034 24032 78036 24041
rect 78088 24032 78090 24041
rect 77116 23724 77168 23730
rect 77116 23666 77168 23672
rect 77128 23526 77156 23666
rect 77312 23662 77340 24006
rect 78034 23967 78090 23976
rect 77300 23656 77352 23662
rect 77300 23598 77352 23604
rect 77116 23520 77168 23526
rect 77116 23462 77168 23468
rect 77852 23520 77904 23526
rect 77852 23462 77904 23468
rect 77128 23186 77156 23462
rect 77864 23361 77892 23462
rect 77850 23352 77906 23361
rect 77850 23287 77906 23296
rect 77116 23180 77168 23186
rect 77116 23122 77168 23128
rect 77300 22976 77352 22982
rect 77300 22918 77352 22924
rect 78036 22976 78088 22982
rect 78036 22918 78088 22924
rect 77312 22506 77340 22918
rect 78048 22681 78076 22918
rect 78034 22672 78090 22681
rect 78034 22607 78090 22616
rect 77300 22500 77352 22506
rect 77300 22442 77352 22448
rect 78034 21992 78090 22001
rect 78034 21927 78090 21936
rect 78048 21894 78076 21927
rect 78036 21888 78088 21894
rect 78036 21830 78088 21836
rect 77116 21344 77168 21350
rect 77852 21344 77904 21350
rect 77116 21286 77168 21292
rect 77850 21312 77852 21321
rect 77904 21312 77906 21321
rect 77128 20806 77156 21286
rect 77850 21247 77906 21256
rect 77116 20800 77168 20806
rect 77116 20742 77168 20748
rect 78036 20800 78088 20806
rect 78036 20742 78088 20748
rect 78048 20641 78076 20742
rect 78034 20632 78090 20641
rect 78034 20567 78090 20576
rect 77852 20256 77904 20262
rect 77852 20198 77904 20204
rect 77864 19961 77892 20198
rect 77850 19952 77906 19961
rect 77850 19887 77906 19896
rect 77852 19508 77904 19514
rect 77852 19450 77904 19456
rect 77864 19281 77892 19450
rect 77850 19272 77906 19281
rect 77850 19207 77906 19216
rect 78036 18624 78088 18630
rect 78034 18592 78036 18601
rect 78088 18592 78090 18601
rect 78034 18527 78090 18536
rect 77116 18284 77168 18290
rect 77116 18226 77168 18232
rect 77128 18086 77156 18226
rect 77116 18080 77168 18086
rect 77116 18022 77168 18028
rect 77852 18080 77904 18086
rect 77852 18022 77904 18028
rect 77024 17536 77076 17542
rect 77024 17478 77076 17484
rect 77036 16658 77064 17478
rect 77128 16998 77156 18022
rect 77864 17921 77892 18022
rect 77850 17912 77906 17921
rect 77850 17847 77906 17856
rect 78036 17536 78088 17542
rect 78036 17478 78088 17484
rect 78048 17241 78076 17478
rect 78034 17232 78090 17241
rect 78034 17167 78090 17176
rect 77116 16992 77168 16998
rect 77116 16934 77168 16940
rect 77024 16652 77076 16658
rect 77024 16594 77076 16600
rect 78034 16552 78090 16561
rect 78034 16487 78090 16496
rect 78048 16454 78076 16487
rect 78036 16448 78088 16454
rect 78036 16390 78088 16396
rect 77852 15904 77904 15910
rect 77850 15872 77852 15881
rect 77904 15872 77906 15881
rect 77850 15807 77906 15816
rect 78036 15360 78088 15366
rect 78036 15302 78088 15308
rect 78048 15201 78076 15302
rect 78034 15192 78090 15201
rect 78034 15127 78090 15136
rect 77852 14816 77904 14822
rect 77852 14758 77904 14764
rect 77864 14521 77892 14758
rect 77850 14512 77906 14521
rect 77850 14447 77906 14456
rect 77852 14068 77904 14074
rect 77852 14010 77904 14016
rect 77864 13841 77892 14010
rect 77850 13832 77906 13841
rect 77850 13767 77906 13776
rect 78036 13184 78088 13190
rect 78034 13152 78036 13161
rect 78088 13152 78090 13161
rect 78034 13087 78090 13096
rect 77116 12844 77168 12850
rect 77116 12786 77168 12792
rect 77128 12646 77156 12786
rect 77116 12640 77168 12646
rect 77116 12582 77168 12588
rect 77852 12640 77904 12646
rect 77852 12582 77904 12588
rect 77128 12102 77156 12582
rect 77864 12481 77892 12582
rect 77850 12472 77906 12481
rect 77850 12407 77906 12416
rect 77116 12096 77168 12102
rect 77116 12038 77168 12044
rect 77300 12096 77352 12102
rect 77300 12038 77352 12044
rect 78036 12096 78088 12102
rect 78036 12038 78088 12044
rect 77312 11558 77340 12038
rect 78048 11801 78076 12038
rect 78034 11792 78090 11801
rect 78034 11727 78090 11736
rect 77300 11552 77352 11558
rect 77300 11494 77352 11500
rect 78036 11280 78088 11286
rect 78036 11222 78088 11228
rect 78048 11121 78076 11222
rect 78034 11112 78090 11121
rect 78034 11047 78090 11056
rect 77116 10464 77168 10470
rect 77852 10464 77904 10470
rect 77116 10406 77168 10412
rect 77850 10432 77852 10441
rect 77904 10432 77906 10441
rect 77128 9994 77156 10406
rect 77850 10367 77906 10376
rect 77116 9988 77168 9994
rect 77116 9930 77168 9936
rect 78036 9920 78088 9926
rect 78036 9862 78088 9868
rect 78048 9761 78076 9862
rect 78034 9752 78090 9761
rect 78034 9687 78090 9696
rect 77852 9376 77904 9382
rect 77852 9318 77904 9324
rect 77864 9081 77892 9318
rect 77850 9072 77906 9081
rect 77850 9007 77906 9016
rect 77850 8392 77906 8401
rect 77116 8356 77168 8362
rect 77850 8327 77852 8336
rect 77116 8298 77168 8304
rect 77904 8327 77906 8336
rect 77852 8298 77904 8304
rect 77024 7812 77076 7818
rect 77024 7754 77076 7760
rect 77036 7274 77064 7754
rect 77128 7750 77156 8298
rect 77116 7744 77168 7750
rect 78036 7744 78088 7750
rect 77116 7686 77168 7692
rect 78034 7712 78036 7721
rect 78088 7712 78090 7721
rect 78034 7647 78090 7656
rect 77024 7268 77076 7274
rect 77024 7210 77076 7216
rect 77852 7200 77904 7206
rect 77852 7142 77904 7148
rect 77864 7041 77892 7142
rect 77850 7032 77906 7041
rect 77850 6967 77906 6976
rect 77300 6656 77352 6662
rect 77300 6598 77352 6604
rect 78036 6656 78088 6662
rect 78036 6598 78088 6604
rect 77312 6118 77340 6598
rect 78048 6361 78076 6598
rect 78034 6352 78090 6361
rect 78034 6287 78090 6296
rect 77300 6112 77352 6118
rect 77300 6054 77352 6060
rect 78034 5672 78090 5681
rect 78034 5607 78090 5616
rect 78048 5574 78076 5607
rect 78036 5568 78088 5574
rect 78036 5510 78088 5516
rect 77852 5024 77904 5030
rect 77850 4992 77852 5001
rect 77904 4992 77906 5001
rect 77850 4927 77906 4936
rect 77852 3392 77904 3398
rect 77852 3334 77904 3340
rect 77864 3058 77892 3334
rect 77852 3052 77904 3058
rect 77852 2994 77904 3000
rect 77114 2952 77170 2961
rect 77114 2887 77116 2896
rect 77168 2887 77170 2896
rect 77392 2916 77444 2922
rect 77116 2858 77168 2864
rect 77392 2858 77444 2864
rect 76380 2848 76432 2854
rect 76380 2790 76432 2796
rect 76288 2644 76340 2650
rect 76288 2586 76340 2592
rect 76392 2446 76420 2790
rect 77404 2446 77432 2858
rect 75920 2440 75972 2446
rect 75656 2400 75920 2428
rect 75656 800 75684 2400
rect 75920 2382 75972 2388
rect 76380 2440 76432 2446
rect 76380 2382 76432 2388
rect 77392 2440 77444 2446
rect 77392 2382 77444 2388
rect 76392 800 76420 2382
rect 77116 2304 77168 2310
rect 77116 2246 77168 2252
rect 77128 800 77156 2246
rect 77864 800 77892 2994
rect 74276 734 74488 762
rect 74906 0 74962 800
rect 75642 0 75698 800
rect 76378 0 76434 800
rect 77114 0 77170 800
rect 77850 0 77906 800
<< via2 >>
rect 4220 77818 4276 77820
rect 4300 77818 4356 77820
rect 4380 77818 4436 77820
rect 4460 77818 4516 77820
rect 4220 77766 4266 77818
rect 4266 77766 4276 77818
rect 4300 77766 4330 77818
rect 4330 77766 4342 77818
rect 4342 77766 4356 77818
rect 4380 77766 4394 77818
rect 4394 77766 4406 77818
rect 4406 77766 4436 77818
rect 4460 77766 4470 77818
rect 4470 77766 4516 77818
rect 4220 77764 4276 77766
rect 4300 77764 4356 77766
rect 4380 77764 4436 77766
rect 4460 77764 4516 77766
rect 34940 77818 34996 77820
rect 35020 77818 35076 77820
rect 35100 77818 35156 77820
rect 35180 77818 35236 77820
rect 34940 77766 34986 77818
rect 34986 77766 34996 77818
rect 35020 77766 35050 77818
rect 35050 77766 35062 77818
rect 35062 77766 35076 77818
rect 35100 77766 35114 77818
rect 35114 77766 35126 77818
rect 35126 77766 35156 77818
rect 35180 77766 35190 77818
rect 35190 77766 35236 77818
rect 34940 77764 34996 77766
rect 35020 77764 35076 77766
rect 35100 77764 35156 77766
rect 35180 77764 35236 77766
rect 65660 77818 65716 77820
rect 65740 77818 65796 77820
rect 65820 77818 65876 77820
rect 65900 77818 65956 77820
rect 65660 77766 65706 77818
rect 65706 77766 65716 77818
rect 65740 77766 65770 77818
rect 65770 77766 65782 77818
rect 65782 77766 65796 77818
rect 65820 77766 65834 77818
rect 65834 77766 65846 77818
rect 65846 77766 65876 77818
rect 65900 77766 65910 77818
rect 65910 77766 65956 77818
rect 65660 77764 65716 77766
rect 65740 77764 65796 77766
rect 65820 77764 65876 77766
rect 65900 77764 65956 77766
rect 19580 77274 19636 77276
rect 19660 77274 19716 77276
rect 19740 77274 19796 77276
rect 19820 77274 19876 77276
rect 19580 77222 19626 77274
rect 19626 77222 19636 77274
rect 19660 77222 19690 77274
rect 19690 77222 19702 77274
rect 19702 77222 19716 77274
rect 19740 77222 19754 77274
rect 19754 77222 19766 77274
rect 19766 77222 19796 77274
rect 19820 77222 19830 77274
rect 19830 77222 19876 77274
rect 19580 77220 19636 77222
rect 19660 77220 19716 77222
rect 19740 77220 19796 77222
rect 19820 77220 19876 77222
rect 50300 77274 50356 77276
rect 50380 77274 50436 77276
rect 50460 77274 50516 77276
rect 50540 77274 50596 77276
rect 50300 77222 50346 77274
rect 50346 77222 50356 77274
rect 50380 77222 50410 77274
rect 50410 77222 50422 77274
rect 50422 77222 50436 77274
rect 50460 77222 50474 77274
rect 50474 77222 50486 77274
rect 50486 77222 50516 77274
rect 50540 77222 50550 77274
rect 50550 77222 50596 77274
rect 50300 77220 50356 77222
rect 50380 77220 50436 77222
rect 50460 77220 50516 77222
rect 50540 77220 50596 77222
rect 4220 76730 4276 76732
rect 4300 76730 4356 76732
rect 4380 76730 4436 76732
rect 4460 76730 4516 76732
rect 4220 76678 4266 76730
rect 4266 76678 4276 76730
rect 4300 76678 4330 76730
rect 4330 76678 4342 76730
rect 4342 76678 4356 76730
rect 4380 76678 4394 76730
rect 4394 76678 4406 76730
rect 4406 76678 4436 76730
rect 4460 76678 4470 76730
rect 4470 76678 4516 76730
rect 4220 76676 4276 76678
rect 4300 76676 4356 76678
rect 4380 76676 4436 76678
rect 4460 76676 4516 76678
rect 34940 76730 34996 76732
rect 35020 76730 35076 76732
rect 35100 76730 35156 76732
rect 35180 76730 35236 76732
rect 34940 76678 34986 76730
rect 34986 76678 34996 76730
rect 35020 76678 35050 76730
rect 35050 76678 35062 76730
rect 35062 76678 35076 76730
rect 35100 76678 35114 76730
rect 35114 76678 35126 76730
rect 35126 76678 35156 76730
rect 35180 76678 35190 76730
rect 35190 76678 35236 76730
rect 34940 76676 34996 76678
rect 35020 76676 35076 76678
rect 35100 76676 35156 76678
rect 35180 76676 35236 76678
rect 65660 76730 65716 76732
rect 65740 76730 65796 76732
rect 65820 76730 65876 76732
rect 65900 76730 65956 76732
rect 65660 76678 65706 76730
rect 65706 76678 65716 76730
rect 65740 76678 65770 76730
rect 65770 76678 65782 76730
rect 65782 76678 65796 76730
rect 65820 76678 65834 76730
rect 65834 76678 65846 76730
rect 65846 76678 65876 76730
rect 65900 76678 65910 76730
rect 65910 76678 65956 76730
rect 65660 76676 65716 76678
rect 65740 76676 65796 76678
rect 65820 76676 65876 76678
rect 65900 76676 65956 76678
rect 19580 76186 19636 76188
rect 19660 76186 19716 76188
rect 19740 76186 19796 76188
rect 19820 76186 19876 76188
rect 19580 76134 19626 76186
rect 19626 76134 19636 76186
rect 19660 76134 19690 76186
rect 19690 76134 19702 76186
rect 19702 76134 19716 76186
rect 19740 76134 19754 76186
rect 19754 76134 19766 76186
rect 19766 76134 19796 76186
rect 19820 76134 19830 76186
rect 19830 76134 19876 76186
rect 19580 76132 19636 76134
rect 19660 76132 19716 76134
rect 19740 76132 19796 76134
rect 19820 76132 19876 76134
rect 50300 76186 50356 76188
rect 50380 76186 50436 76188
rect 50460 76186 50516 76188
rect 50540 76186 50596 76188
rect 50300 76134 50346 76186
rect 50346 76134 50356 76186
rect 50380 76134 50410 76186
rect 50410 76134 50422 76186
rect 50422 76134 50436 76186
rect 50460 76134 50474 76186
rect 50474 76134 50486 76186
rect 50486 76134 50516 76186
rect 50540 76134 50550 76186
rect 50550 76134 50596 76186
rect 50300 76132 50356 76134
rect 50380 76132 50436 76134
rect 50460 76132 50516 76134
rect 50540 76132 50596 76134
rect 4220 75642 4276 75644
rect 4300 75642 4356 75644
rect 4380 75642 4436 75644
rect 4460 75642 4516 75644
rect 4220 75590 4266 75642
rect 4266 75590 4276 75642
rect 4300 75590 4330 75642
rect 4330 75590 4342 75642
rect 4342 75590 4356 75642
rect 4380 75590 4394 75642
rect 4394 75590 4406 75642
rect 4406 75590 4436 75642
rect 4460 75590 4470 75642
rect 4470 75590 4516 75642
rect 4220 75588 4276 75590
rect 4300 75588 4356 75590
rect 4380 75588 4436 75590
rect 4460 75588 4516 75590
rect 34940 75642 34996 75644
rect 35020 75642 35076 75644
rect 35100 75642 35156 75644
rect 35180 75642 35236 75644
rect 34940 75590 34986 75642
rect 34986 75590 34996 75642
rect 35020 75590 35050 75642
rect 35050 75590 35062 75642
rect 35062 75590 35076 75642
rect 35100 75590 35114 75642
rect 35114 75590 35126 75642
rect 35126 75590 35156 75642
rect 35180 75590 35190 75642
rect 35190 75590 35236 75642
rect 34940 75588 34996 75590
rect 35020 75588 35076 75590
rect 35100 75588 35156 75590
rect 35180 75588 35236 75590
rect 65660 75642 65716 75644
rect 65740 75642 65796 75644
rect 65820 75642 65876 75644
rect 65900 75642 65956 75644
rect 65660 75590 65706 75642
rect 65706 75590 65716 75642
rect 65740 75590 65770 75642
rect 65770 75590 65782 75642
rect 65782 75590 65796 75642
rect 65820 75590 65834 75642
rect 65834 75590 65846 75642
rect 65846 75590 65876 75642
rect 65900 75590 65910 75642
rect 65910 75590 65956 75642
rect 65660 75588 65716 75590
rect 65740 75588 65796 75590
rect 65820 75588 65876 75590
rect 65900 75588 65956 75590
rect 1674 75284 1676 75304
rect 1676 75284 1728 75304
rect 1728 75284 1730 75304
rect 1674 75248 1730 75284
rect 19580 75098 19636 75100
rect 19660 75098 19716 75100
rect 19740 75098 19796 75100
rect 19820 75098 19876 75100
rect 19580 75046 19626 75098
rect 19626 75046 19636 75098
rect 19660 75046 19690 75098
rect 19690 75046 19702 75098
rect 19702 75046 19716 75098
rect 19740 75046 19754 75098
rect 19754 75046 19766 75098
rect 19766 75046 19796 75098
rect 19820 75046 19830 75098
rect 19830 75046 19876 75098
rect 19580 75044 19636 75046
rect 19660 75044 19716 75046
rect 19740 75044 19796 75046
rect 19820 75044 19876 75046
rect 50300 75098 50356 75100
rect 50380 75098 50436 75100
rect 50460 75098 50516 75100
rect 50540 75098 50596 75100
rect 50300 75046 50346 75098
rect 50346 75046 50356 75098
rect 50380 75046 50410 75098
rect 50410 75046 50422 75098
rect 50422 75046 50436 75098
rect 50460 75046 50474 75098
rect 50474 75046 50486 75098
rect 50486 75046 50516 75098
rect 50540 75046 50550 75098
rect 50550 75046 50596 75098
rect 50300 75044 50356 75046
rect 50380 75044 50436 75046
rect 50460 75044 50516 75046
rect 50540 75044 50596 75046
rect 1490 74976 1546 75032
rect 4220 74554 4276 74556
rect 4300 74554 4356 74556
rect 4380 74554 4436 74556
rect 4460 74554 4516 74556
rect 1398 74332 1400 74352
rect 1400 74332 1452 74352
rect 1452 74332 1454 74352
rect 1398 74296 1454 74332
rect 1490 73636 1546 73672
rect 1490 73616 1492 73636
rect 1492 73616 1544 73636
rect 1544 73616 1546 73636
rect 1490 72972 1492 72992
rect 1492 72972 1544 72992
rect 1544 72972 1546 72992
rect 1490 72936 1546 72972
rect 1490 72256 1546 72312
rect 1490 71576 1546 71632
rect 1490 70896 1546 70952
rect 1490 70252 1492 70272
rect 1492 70252 1544 70272
rect 1544 70252 1546 70272
rect 1490 70216 1546 70252
rect 1398 69536 1454 69592
rect 1398 68856 1454 68912
rect 1398 68176 1454 68232
rect 1398 67496 1454 67552
rect 1398 66816 1454 66872
rect 1398 66136 1454 66192
rect 1398 65492 1400 65512
rect 1400 65492 1452 65512
rect 1452 65492 1454 65512
rect 1398 65456 1454 65492
rect 1398 64776 1454 64832
rect 1398 64096 1454 64152
rect 1398 63416 1454 63472
rect 1398 62736 1454 62792
rect 1398 62056 1454 62112
rect 1398 61376 1454 61432
rect 1398 60696 1454 60752
rect 1398 60052 1400 60072
rect 1400 60052 1452 60072
rect 1452 60052 1454 60072
rect 1398 60016 1454 60052
rect 1398 59336 1454 59392
rect 1398 58656 1454 58712
rect 1398 57976 1454 58032
rect 1674 60152 1730 60208
rect 1858 59608 1914 59664
rect 1398 57296 1454 57352
rect 1398 56616 1454 56672
rect 1398 55936 1454 55992
rect 1490 55256 1546 55312
rect 1490 54612 1492 54632
rect 1492 54612 1544 54632
rect 1544 54612 1546 54632
rect 1490 54576 1546 54612
rect 1490 53896 1546 53952
rect 1490 53216 1546 53272
rect 1490 52536 1546 52592
rect 1490 51856 1546 51912
rect 1490 51176 1546 51232
rect 1490 50496 1546 50552
rect 4220 74502 4266 74554
rect 4266 74502 4276 74554
rect 4300 74502 4330 74554
rect 4330 74502 4342 74554
rect 4342 74502 4356 74554
rect 4380 74502 4394 74554
rect 4394 74502 4406 74554
rect 4406 74502 4436 74554
rect 4460 74502 4470 74554
rect 4470 74502 4516 74554
rect 4220 74500 4276 74502
rect 4300 74500 4356 74502
rect 4380 74500 4436 74502
rect 4460 74500 4516 74502
rect 34940 74554 34996 74556
rect 35020 74554 35076 74556
rect 35100 74554 35156 74556
rect 35180 74554 35236 74556
rect 34940 74502 34986 74554
rect 34986 74502 34996 74554
rect 35020 74502 35050 74554
rect 35050 74502 35062 74554
rect 35062 74502 35076 74554
rect 35100 74502 35114 74554
rect 35114 74502 35126 74554
rect 35126 74502 35156 74554
rect 35180 74502 35190 74554
rect 35190 74502 35236 74554
rect 34940 74500 34996 74502
rect 35020 74500 35076 74502
rect 35100 74500 35156 74502
rect 35180 74500 35236 74502
rect 65660 74554 65716 74556
rect 65740 74554 65796 74556
rect 65820 74554 65876 74556
rect 65900 74554 65956 74556
rect 65660 74502 65706 74554
rect 65706 74502 65716 74554
rect 65740 74502 65770 74554
rect 65770 74502 65782 74554
rect 65782 74502 65796 74554
rect 65820 74502 65834 74554
rect 65834 74502 65846 74554
rect 65846 74502 65876 74554
rect 65900 74502 65910 74554
rect 65910 74502 65956 74554
rect 65660 74500 65716 74502
rect 65740 74500 65796 74502
rect 65820 74500 65876 74502
rect 65900 74500 65956 74502
rect 19580 74010 19636 74012
rect 19660 74010 19716 74012
rect 19740 74010 19796 74012
rect 19820 74010 19876 74012
rect 19580 73958 19626 74010
rect 19626 73958 19636 74010
rect 19660 73958 19690 74010
rect 19690 73958 19702 74010
rect 19702 73958 19716 74010
rect 19740 73958 19754 74010
rect 19754 73958 19766 74010
rect 19766 73958 19796 74010
rect 19820 73958 19830 74010
rect 19830 73958 19876 74010
rect 19580 73956 19636 73958
rect 19660 73956 19716 73958
rect 19740 73956 19796 73958
rect 19820 73956 19876 73958
rect 50300 74010 50356 74012
rect 50380 74010 50436 74012
rect 50460 74010 50516 74012
rect 50540 74010 50596 74012
rect 50300 73958 50346 74010
rect 50346 73958 50356 74010
rect 50380 73958 50410 74010
rect 50410 73958 50422 74010
rect 50422 73958 50436 74010
rect 50460 73958 50474 74010
rect 50474 73958 50486 74010
rect 50486 73958 50516 74010
rect 50540 73958 50550 74010
rect 50550 73958 50596 74010
rect 50300 73956 50356 73958
rect 50380 73956 50436 73958
rect 50460 73956 50516 73958
rect 50540 73956 50596 73958
rect 4220 73466 4276 73468
rect 4300 73466 4356 73468
rect 4380 73466 4436 73468
rect 4460 73466 4516 73468
rect 4220 73414 4266 73466
rect 4266 73414 4276 73466
rect 4300 73414 4330 73466
rect 4330 73414 4342 73466
rect 4342 73414 4356 73466
rect 4380 73414 4394 73466
rect 4394 73414 4406 73466
rect 4406 73414 4436 73466
rect 4460 73414 4470 73466
rect 4470 73414 4516 73466
rect 4220 73412 4276 73414
rect 4300 73412 4356 73414
rect 4380 73412 4436 73414
rect 4460 73412 4516 73414
rect 34940 73466 34996 73468
rect 35020 73466 35076 73468
rect 35100 73466 35156 73468
rect 35180 73466 35236 73468
rect 34940 73414 34986 73466
rect 34986 73414 34996 73466
rect 35020 73414 35050 73466
rect 35050 73414 35062 73466
rect 35062 73414 35076 73466
rect 35100 73414 35114 73466
rect 35114 73414 35126 73466
rect 35126 73414 35156 73466
rect 35180 73414 35190 73466
rect 35190 73414 35236 73466
rect 34940 73412 34996 73414
rect 35020 73412 35076 73414
rect 35100 73412 35156 73414
rect 35180 73412 35236 73414
rect 65660 73466 65716 73468
rect 65740 73466 65796 73468
rect 65820 73466 65876 73468
rect 65900 73466 65956 73468
rect 65660 73414 65706 73466
rect 65706 73414 65716 73466
rect 65740 73414 65770 73466
rect 65770 73414 65782 73466
rect 65782 73414 65796 73466
rect 65820 73414 65834 73466
rect 65834 73414 65846 73466
rect 65846 73414 65876 73466
rect 65900 73414 65910 73466
rect 65910 73414 65956 73466
rect 65660 73412 65716 73414
rect 65740 73412 65796 73414
rect 65820 73412 65876 73414
rect 65900 73412 65956 73414
rect 19580 72922 19636 72924
rect 19660 72922 19716 72924
rect 19740 72922 19796 72924
rect 19820 72922 19876 72924
rect 19580 72870 19626 72922
rect 19626 72870 19636 72922
rect 19660 72870 19690 72922
rect 19690 72870 19702 72922
rect 19702 72870 19716 72922
rect 19740 72870 19754 72922
rect 19754 72870 19766 72922
rect 19766 72870 19796 72922
rect 19820 72870 19830 72922
rect 19830 72870 19876 72922
rect 19580 72868 19636 72870
rect 19660 72868 19716 72870
rect 19740 72868 19796 72870
rect 19820 72868 19876 72870
rect 50300 72922 50356 72924
rect 50380 72922 50436 72924
rect 50460 72922 50516 72924
rect 50540 72922 50596 72924
rect 50300 72870 50346 72922
rect 50346 72870 50356 72922
rect 50380 72870 50410 72922
rect 50410 72870 50422 72922
rect 50422 72870 50436 72922
rect 50460 72870 50474 72922
rect 50474 72870 50486 72922
rect 50486 72870 50516 72922
rect 50540 72870 50550 72922
rect 50550 72870 50596 72922
rect 50300 72868 50356 72870
rect 50380 72868 50436 72870
rect 50460 72868 50516 72870
rect 50540 72868 50596 72870
rect 4220 72378 4276 72380
rect 4300 72378 4356 72380
rect 4380 72378 4436 72380
rect 4460 72378 4516 72380
rect 4220 72326 4266 72378
rect 4266 72326 4276 72378
rect 4300 72326 4330 72378
rect 4330 72326 4342 72378
rect 4342 72326 4356 72378
rect 4380 72326 4394 72378
rect 4394 72326 4406 72378
rect 4406 72326 4436 72378
rect 4460 72326 4470 72378
rect 4470 72326 4516 72378
rect 4220 72324 4276 72326
rect 4300 72324 4356 72326
rect 4380 72324 4436 72326
rect 4460 72324 4516 72326
rect 34940 72378 34996 72380
rect 35020 72378 35076 72380
rect 35100 72378 35156 72380
rect 35180 72378 35236 72380
rect 34940 72326 34986 72378
rect 34986 72326 34996 72378
rect 35020 72326 35050 72378
rect 35050 72326 35062 72378
rect 35062 72326 35076 72378
rect 35100 72326 35114 72378
rect 35114 72326 35126 72378
rect 35126 72326 35156 72378
rect 35180 72326 35190 72378
rect 35190 72326 35236 72378
rect 34940 72324 34996 72326
rect 35020 72324 35076 72326
rect 35100 72324 35156 72326
rect 35180 72324 35236 72326
rect 65660 72378 65716 72380
rect 65740 72378 65796 72380
rect 65820 72378 65876 72380
rect 65900 72378 65956 72380
rect 65660 72326 65706 72378
rect 65706 72326 65716 72378
rect 65740 72326 65770 72378
rect 65770 72326 65782 72378
rect 65782 72326 65796 72378
rect 65820 72326 65834 72378
rect 65834 72326 65846 72378
rect 65846 72326 65876 72378
rect 65900 72326 65910 72378
rect 65910 72326 65956 72378
rect 65660 72324 65716 72326
rect 65740 72324 65796 72326
rect 65820 72324 65876 72326
rect 65900 72324 65956 72326
rect 19580 71834 19636 71836
rect 19660 71834 19716 71836
rect 19740 71834 19796 71836
rect 19820 71834 19876 71836
rect 19580 71782 19626 71834
rect 19626 71782 19636 71834
rect 19660 71782 19690 71834
rect 19690 71782 19702 71834
rect 19702 71782 19716 71834
rect 19740 71782 19754 71834
rect 19754 71782 19766 71834
rect 19766 71782 19796 71834
rect 19820 71782 19830 71834
rect 19830 71782 19876 71834
rect 19580 71780 19636 71782
rect 19660 71780 19716 71782
rect 19740 71780 19796 71782
rect 19820 71780 19876 71782
rect 50300 71834 50356 71836
rect 50380 71834 50436 71836
rect 50460 71834 50516 71836
rect 50540 71834 50596 71836
rect 50300 71782 50346 71834
rect 50346 71782 50356 71834
rect 50380 71782 50410 71834
rect 50410 71782 50422 71834
rect 50422 71782 50436 71834
rect 50460 71782 50474 71834
rect 50474 71782 50486 71834
rect 50486 71782 50516 71834
rect 50540 71782 50550 71834
rect 50550 71782 50596 71834
rect 50300 71780 50356 71782
rect 50380 71780 50436 71782
rect 50460 71780 50516 71782
rect 50540 71780 50596 71782
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 34940 71290 34996 71292
rect 35020 71290 35076 71292
rect 35100 71290 35156 71292
rect 35180 71290 35236 71292
rect 34940 71238 34986 71290
rect 34986 71238 34996 71290
rect 35020 71238 35050 71290
rect 35050 71238 35062 71290
rect 35062 71238 35076 71290
rect 35100 71238 35114 71290
rect 35114 71238 35126 71290
rect 35126 71238 35156 71290
rect 35180 71238 35190 71290
rect 35190 71238 35236 71290
rect 34940 71236 34996 71238
rect 35020 71236 35076 71238
rect 35100 71236 35156 71238
rect 35180 71236 35236 71238
rect 65660 71290 65716 71292
rect 65740 71290 65796 71292
rect 65820 71290 65876 71292
rect 65900 71290 65956 71292
rect 65660 71238 65706 71290
rect 65706 71238 65716 71290
rect 65740 71238 65770 71290
rect 65770 71238 65782 71290
rect 65782 71238 65796 71290
rect 65820 71238 65834 71290
rect 65834 71238 65846 71290
rect 65846 71238 65876 71290
rect 65900 71238 65910 71290
rect 65910 71238 65956 71290
rect 65660 71236 65716 71238
rect 65740 71236 65796 71238
rect 65820 71236 65876 71238
rect 65900 71236 65956 71238
rect 19580 70746 19636 70748
rect 19660 70746 19716 70748
rect 19740 70746 19796 70748
rect 19820 70746 19876 70748
rect 19580 70694 19626 70746
rect 19626 70694 19636 70746
rect 19660 70694 19690 70746
rect 19690 70694 19702 70746
rect 19702 70694 19716 70746
rect 19740 70694 19754 70746
rect 19754 70694 19766 70746
rect 19766 70694 19796 70746
rect 19820 70694 19830 70746
rect 19830 70694 19876 70746
rect 19580 70692 19636 70694
rect 19660 70692 19716 70694
rect 19740 70692 19796 70694
rect 19820 70692 19876 70694
rect 50300 70746 50356 70748
rect 50380 70746 50436 70748
rect 50460 70746 50516 70748
rect 50540 70746 50596 70748
rect 50300 70694 50346 70746
rect 50346 70694 50356 70746
rect 50380 70694 50410 70746
rect 50410 70694 50422 70746
rect 50422 70694 50436 70746
rect 50460 70694 50474 70746
rect 50474 70694 50486 70746
rect 50486 70694 50516 70746
rect 50540 70694 50550 70746
rect 50550 70694 50596 70746
rect 50300 70692 50356 70694
rect 50380 70692 50436 70694
rect 50460 70692 50516 70694
rect 50540 70692 50596 70694
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 34940 70202 34996 70204
rect 35020 70202 35076 70204
rect 35100 70202 35156 70204
rect 35180 70202 35236 70204
rect 34940 70150 34986 70202
rect 34986 70150 34996 70202
rect 35020 70150 35050 70202
rect 35050 70150 35062 70202
rect 35062 70150 35076 70202
rect 35100 70150 35114 70202
rect 35114 70150 35126 70202
rect 35126 70150 35156 70202
rect 35180 70150 35190 70202
rect 35190 70150 35236 70202
rect 34940 70148 34996 70150
rect 35020 70148 35076 70150
rect 35100 70148 35156 70150
rect 35180 70148 35236 70150
rect 65660 70202 65716 70204
rect 65740 70202 65796 70204
rect 65820 70202 65876 70204
rect 65900 70202 65956 70204
rect 65660 70150 65706 70202
rect 65706 70150 65716 70202
rect 65740 70150 65770 70202
rect 65770 70150 65782 70202
rect 65782 70150 65796 70202
rect 65820 70150 65834 70202
rect 65834 70150 65846 70202
rect 65846 70150 65876 70202
rect 65900 70150 65910 70202
rect 65910 70150 65956 70202
rect 65660 70148 65716 70150
rect 65740 70148 65796 70150
rect 65820 70148 65876 70150
rect 65900 70148 65956 70150
rect 19580 69658 19636 69660
rect 19660 69658 19716 69660
rect 19740 69658 19796 69660
rect 19820 69658 19876 69660
rect 19580 69606 19626 69658
rect 19626 69606 19636 69658
rect 19660 69606 19690 69658
rect 19690 69606 19702 69658
rect 19702 69606 19716 69658
rect 19740 69606 19754 69658
rect 19754 69606 19766 69658
rect 19766 69606 19796 69658
rect 19820 69606 19830 69658
rect 19830 69606 19876 69658
rect 19580 69604 19636 69606
rect 19660 69604 19716 69606
rect 19740 69604 19796 69606
rect 19820 69604 19876 69606
rect 50300 69658 50356 69660
rect 50380 69658 50436 69660
rect 50460 69658 50516 69660
rect 50540 69658 50596 69660
rect 50300 69606 50346 69658
rect 50346 69606 50356 69658
rect 50380 69606 50410 69658
rect 50410 69606 50422 69658
rect 50422 69606 50436 69658
rect 50460 69606 50474 69658
rect 50474 69606 50486 69658
rect 50486 69606 50516 69658
rect 50540 69606 50550 69658
rect 50550 69606 50596 69658
rect 50300 69604 50356 69606
rect 50380 69604 50436 69606
rect 50460 69604 50516 69606
rect 50540 69604 50596 69606
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 34940 69114 34996 69116
rect 35020 69114 35076 69116
rect 35100 69114 35156 69116
rect 35180 69114 35236 69116
rect 34940 69062 34986 69114
rect 34986 69062 34996 69114
rect 35020 69062 35050 69114
rect 35050 69062 35062 69114
rect 35062 69062 35076 69114
rect 35100 69062 35114 69114
rect 35114 69062 35126 69114
rect 35126 69062 35156 69114
rect 35180 69062 35190 69114
rect 35190 69062 35236 69114
rect 34940 69060 34996 69062
rect 35020 69060 35076 69062
rect 35100 69060 35156 69062
rect 35180 69060 35236 69062
rect 65660 69114 65716 69116
rect 65740 69114 65796 69116
rect 65820 69114 65876 69116
rect 65900 69114 65956 69116
rect 65660 69062 65706 69114
rect 65706 69062 65716 69114
rect 65740 69062 65770 69114
rect 65770 69062 65782 69114
rect 65782 69062 65796 69114
rect 65820 69062 65834 69114
rect 65834 69062 65846 69114
rect 65846 69062 65876 69114
rect 65900 69062 65910 69114
rect 65910 69062 65956 69114
rect 65660 69060 65716 69062
rect 65740 69060 65796 69062
rect 65820 69060 65876 69062
rect 65900 69060 65956 69062
rect 19580 68570 19636 68572
rect 19660 68570 19716 68572
rect 19740 68570 19796 68572
rect 19820 68570 19876 68572
rect 19580 68518 19626 68570
rect 19626 68518 19636 68570
rect 19660 68518 19690 68570
rect 19690 68518 19702 68570
rect 19702 68518 19716 68570
rect 19740 68518 19754 68570
rect 19754 68518 19766 68570
rect 19766 68518 19796 68570
rect 19820 68518 19830 68570
rect 19830 68518 19876 68570
rect 19580 68516 19636 68518
rect 19660 68516 19716 68518
rect 19740 68516 19796 68518
rect 19820 68516 19876 68518
rect 50300 68570 50356 68572
rect 50380 68570 50436 68572
rect 50460 68570 50516 68572
rect 50540 68570 50596 68572
rect 50300 68518 50346 68570
rect 50346 68518 50356 68570
rect 50380 68518 50410 68570
rect 50410 68518 50422 68570
rect 50422 68518 50436 68570
rect 50460 68518 50474 68570
rect 50474 68518 50486 68570
rect 50486 68518 50516 68570
rect 50540 68518 50550 68570
rect 50550 68518 50596 68570
rect 50300 68516 50356 68518
rect 50380 68516 50436 68518
rect 50460 68516 50516 68518
rect 50540 68516 50596 68518
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 34940 68026 34996 68028
rect 35020 68026 35076 68028
rect 35100 68026 35156 68028
rect 35180 68026 35236 68028
rect 34940 67974 34986 68026
rect 34986 67974 34996 68026
rect 35020 67974 35050 68026
rect 35050 67974 35062 68026
rect 35062 67974 35076 68026
rect 35100 67974 35114 68026
rect 35114 67974 35126 68026
rect 35126 67974 35156 68026
rect 35180 67974 35190 68026
rect 35190 67974 35236 68026
rect 34940 67972 34996 67974
rect 35020 67972 35076 67974
rect 35100 67972 35156 67974
rect 35180 67972 35236 67974
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 19580 67482 19636 67484
rect 19660 67482 19716 67484
rect 19740 67482 19796 67484
rect 19820 67482 19876 67484
rect 19580 67430 19626 67482
rect 19626 67430 19636 67482
rect 19660 67430 19690 67482
rect 19690 67430 19702 67482
rect 19702 67430 19716 67482
rect 19740 67430 19754 67482
rect 19754 67430 19766 67482
rect 19766 67430 19796 67482
rect 19820 67430 19830 67482
rect 19830 67430 19876 67482
rect 19580 67428 19636 67430
rect 19660 67428 19716 67430
rect 19740 67428 19796 67430
rect 19820 67428 19876 67430
rect 50300 67482 50356 67484
rect 50380 67482 50436 67484
rect 50460 67482 50516 67484
rect 50540 67482 50596 67484
rect 50300 67430 50346 67482
rect 50346 67430 50356 67482
rect 50380 67430 50410 67482
rect 50410 67430 50422 67482
rect 50422 67430 50436 67482
rect 50460 67430 50474 67482
rect 50474 67430 50486 67482
rect 50486 67430 50516 67482
rect 50540 67430 50550 67482
rect 50550 67430 50596 67482
rect 50300 67428 50356 67430
rect 50380 67428 50436 67430
rect 50460 67428 50516 67430
rect 50540 67428 50596 67430
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 19580 66394 19636 66396
rect 19660 66394 19716 66396
rect 19740 66394 19796 66396
rect 19820 66394 19876 66396
rect 19580 66342 19626 66394
rect 19626 66342 19636 66394
rect 19660 66342 19690 66394
rect 19690 66342 19702 66394
rect 19702 66342 19716 66394
rect 19740 66342 19754 66394
rect 19754 66342 19766 66394
rect 19766 66342 19796 66394
rect 19820 66342 19830 66394
rect 19830 66342 19876 66394
rect 19580 66340 19636 66342
rect 19660 66340 19716 66342
rect 19740 66340 19796 66342
rect 19820 66340 19876 66342
rect 50300 66394 50356 66396
rect 50380 66394 50436 66396
rect 50460 66394 50516 66396
rect 50540 66394 50596 66396
rect 50300 66342 50346 66394
rect 50346 66342 50356 66394
rect 50380 66342 50410 66394
rect 50410 66342 50422 66394
rect 50422 66342 50436 66394
rect 50460 66342 50474 66394
rect 50474 66342 50486 66394
rect 50486 66342 50516 66394
rect 50540 66342 50550 66394
rect 50550 66342 50596 66394
rect 50300 66340 50356 66342
rect 50380 66340 50436 66342
rect 50460 66340 50516 66342
rect 50540 66340 50596 66342
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 19580 65306 19636 65308
rect 19660 65306 19716 65308
rect 19740 65306 19796 65308
rect 19820 65306 19876 65308
rect 19580 65254 19626 65306
rect 19626 65254 19636 65306
rect 19660 65254 19690 65306
rect 19690 65254 19702 65306
rect 19702 65254 19716 65306
rect 19740 65254 19754 65306
rect 19754 65254 19766 65306
rect 19766 65254 19796 65306
rect 19820 65254 19830 65306
rect 19830 65254 19876 65306
rect 19580 65252 19636 65254
rect 19660 65252 19716 65254
rect 19740 65252 19796 65254
rect 19820 65252 19876 65254
rect 50300 65306 50356 65308
rect 50380 65306 50436 65308
rect 50460 65306 50516 65308
rect 50540 65306 50596 65308
rect 50300 65254 50346 65306
rect 50346 65254 50356 65306
rect 50380 65254 50410 65306
rect 50410 65254 50422 65306
rect 50422 65254 50436 65306
rect 50460 65254 50474 65306
rect 50474 65254 50486 65306
rect 50486 65254 50516 65306
rect 50540 65254 50550 65306
rect 50550 65254 50596 65306
rect 50300 65252 50356 65254
rect 50380 65252 50436 65254
rect 50460 65252 50516 65254
rect 50540 65252 50596 65254
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 34940 64762 34996 64764
rect 35020 64762 35076 64764
rect 35100 64762 35156 64764
rect 35180 64762 35236 64764
rect 34940 64710 34986 64762
rect 34986 64710 34996 64762
rect 35020 64710 35050 64762
rect 35050 64710 35062 64762
rect 35062 64710 35076 64762
rect 35100 64710 35114 64762
rect 35114 64710 35126 64762
rect 35126 64710 35156 64762
rect 35180 64710 35190 64762
rect 35190 64710 35236 64762
rect 34940 64708 34996 64710
rect 35020 64708 35076 64710
rect 35100 64708 35156 64710
rect 35180 64708 35236 64710
rect 19580 64218 19636 64220
rect 19660 64218 19716 64220
rect 19740 64218 19796 64220
rect 19820 64218 19876 64220
rect 19580 64166 19626 64218
rect 19626 64166 19636 64218
rect 19660 64166 19690 64218
rect 19690 64166 19702 64218
rect 19702 64166 19716 64218
rect 19740 64166 19754 64218
rect 19754 64166 19766 64218
rect 19766 64166 19796 64218
rect 19820 64166 19830 64218
rect 19830 64166 19876 64218
rect 19580 64164 19636 64166
rect 19660 64164 19716 64166
rect 19740 64164 19796 64166
rect 19820 64164 19876 64166
rect 50300 64218 50356 64220
rect 50380 64218 50436 64220
rect 50460 64218 50516 64220
rect 50540 64218 50596 64220
rect 50300 64166 50346 64218
rect 50346 64166 50356 64218
rect 50380 64166 50410 64218
rect 50410 64166 50422 64218
rect 50422 64166 50436 64218
rect 50460 64166 50474 64218
rect 50474 64166 50486 64218
rect 50486 64166 50516 64218
rect 50540 64166 50550 64218
rect 50550 64166 50596 64218
rect 50300 64164 50356 64166
rect 50380 64164 50436 64166
rect 50460 64164 50516 64166
rect 50540 64164 50596 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 34940 63674 34996 63676
rect 35020 63674 35076 63676
rect 35100 63674 35156 63676
rect 35180 63674 35236 63676
rect 34940 63622 34986 63674
rect 34986 63622 34996 63674
rect 35020 63622 35050 63674
rect 35050 63622 35062 63674
rect 35062 63622 35076 63674
rect 35100 63622 35114 63674
rect 35114 63622 35126 63674
rect 35126 63622 35156 63674
rect 35180 63622 35190 63674
rect 35190 63622 35236 63674
rect 34940 63620 34996 63622
rect 35020 63620 35076 63622
rect 35100 63620 35156 63622
rect 35180 63620 35236 63622
rect 19580 63130 19636 63132
rect 19660 63130 19716 63132
rect 19740 63130 19796 63132
rect 19820 63130 19876 63132
rect 19580 63078 19626 63130
rect 19626 63078 19636 63130
rect 19660 63078 19690 63130
rect 19690 63078 19702 63130
rect 19702 63078 19716 63130
rect 19740 63078 19754 63130
rect 19754 63078 19766 63130
rect 19766 63078 19796 63130
rect 19820 63078 19830 63130
rect 19830 63078 19876 63130
rect 19580 63076 19636 63078
rect 19660 63076 19716 63078
rect 19740 63076 19796 63078
rect 19820 63076 19876 63078
rect 50300 63130 50356 63132
rect 50380 63130 50436 63132
rect 50460 63130 50516 63132
rect 50540 63130 50596 63132
rect 50300 63078 50346 63130
rect 50346 63078 50356 63130
rect 50380 63078 50410 63130
rect 50410 63078 50422 63130
rect 50422 63078 50436 63130
rect 50460 63078 50474 63130
rect 50474 63078 50486 63130
rect 50486 63078 50516 63130
rect 50540 63078 50550 63130
rect 50550 63078 50596 63130
rect 50300 63076 50356 63078
rect 50380 63076 50436 63078
rect 50460 63076 50516 63078
rect 50540 63076 50596 63078
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 34940 62586 34996 62588
rect 35020 62586 35076 62588
rect 35100 62586 35156 62588
rect 35180 62586 35236 62588
rect 34940 62534 34986 62586
rect 34986 62534 34996 62586
rect 35020 62534 35050 62586
rect 35050 62534 35062 62586
rect 35062 62534 35076 62586
rect 35100 62534 35114 62586
rect 35114 62534 35126 62586
rect 35126 62534 35156 62586
rect 35180 62534 35190 62586
rect 35190 62534 35236 62586
rect 34940 62532 34996 62534
rect 35020 62532 35076 62534
rect 35100 62532 35156 62534
rect 35180 62532 35236 62534
rect 19580 62042 19636 62044
rect 19660 62042 19716 62044
rect 19740 62042 19796 62044
rect 19820 62042 19876 62044
rect 19580 61990 19626 62042
rect 19626 61990 19636 62042
rect 19660 61990 19690 62042
rect 19690 61990 19702 62042
rect 19702 61990 19716 62042
rect 19740 61990 19754 62042
rect 19754 61990 19766 62042
rect 19766 61990 19796 62042
rect 19820 61990 19830 62042
rect 19830 61990 19876 62042
rect 19580 61988 19636 61990
rect 19660 61988 19716 61990
rect 19740 61988 19796 61990
rect 19820 61988 19876 61990
rect 50300 62042 50356 62044
rect 50380 62042 50436 62044
rect 50460 62042 50516 62044
rect 50540 62042 50596 62044
rect 50300 61990 50346 62042
rect 50346 61990 50356 62042
rect 50380 61990 50410 62042
rect 50410 61990 50422 62042
rect 50422 61990 50436 62042
rect 50460 61990 50474 62042
rect 50474 61990 50486 62042
rect 50486 61990 50516 62042
rect 50540 61990 50550 62042
rect 50550 61990 50596 62042
rect 50300 61988 50356 61990
rect 50380 61988 50436 61990
rect 50460 61988 50516 61990
rect 50540 61988 50596 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 19580 60954 19636 60956
rect 19660 60954 19716 60956
rect 19740 60954 19796 60956
rect 19820 60954 19876 60956
rect 19580 60902 19626 60954
rect 19626 60902 19636 60954
rect 19660 60902 19690 60954
rect 19690 60902 19702 60954
rect 19702 60902 19716 60954
rect 19740 60902 19754 60954
rect 19754 60902 19766 60954
rect 19766 60902 19796 60954
rect 19820 60902 19830 60954
rect 19830 60902 19876 60954
rect 19580 60900 19636 60902
rect 19660 60900 19716 60902
rect 19740 60900 19796 60902
rect 19820 60900 19876 60902
rect 50300 60954 50356 60956
rect 50380 60954 50436 60956
rect 50460 60954 50516 60956
rect 50540 60954 50596 60956
rect 50300 60902 50346 60954
rect 50346 60902 50356 60954
rect 50380 60902 50410 60954
rect 50410 60902 50422 60954
rect 50422 60902 50436 60954
rect 50460 60902 50474 60954
rect 50474 60902 50486 60954
rect 50486 60902 50516 60954
rect 50540 60902 50550 60954
rect 50550 60902 50596 60954
rect 50300 60900 50356 60902
rect 50380 60900 50436 60902
rect 50460 60900 50516 60902
rect 50540 60900 50596 60902
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 19580 59866 19636 59868
rect 19660 59866 19716 59868
rect 19740 59866 19796 59868
rect 19820 59866 19876 59868
rect 19580 59814 19626 59866
rect 19626 59814 19636 59866
rect 19660 59814 19690 59866
rect 19690 59814 19702 59866
rect 19702 59814 19716 59866
rect 19740 59814 19754 59866
rect 19754 59814 19766 59866
rect 19766 59814 19796 59866
rect 19820 59814 19830 59866
rect 19830 59814 19876 59866
rect 19580 59812 19636 59814
rect 19660 59812 19716 59814
rect 19740 59812 19796 59814
rect 19820 59812 19876 59814
rect 50300 59866 50356 59868
rect 50380 59866 50436 59868
rect 50460 59866 50516 59868
rect 50540 59866 50596 59868
rect 50300 59814 50346 59866
rect 50346 59814 50356 59866
rect 50380 59814 50410 59866
rect 50410 59814 50422 59866
rect 50422 59814 50436 59866
rect 50460 59814 50474 59866
rect 50474 59814 50486 59866
rect 50486 59814 50516 59866
rect 50540 59814 50550 59866
rect 50550 59814 50596 59866
rect 50300 59812 50356 59814
rect 50380 59812 50436 59814
rect 50460 59812 50516 59814
rect 50540 59812 50596 59814
rect 4220 59322 4276 59324
rect 4300 59322 4356 59324
rect 4380 59322 4436 59324
rect 4460 59322 4516 59324
rect 4220 59270 4266 59322
rect 4266 59270 4276 59322
rect 4300 59270 4330 59322
rect 4330 59270 4342 59322
rect 4342 59270 4356 59322
rect 4380 59270 4394 59322
rect 4394 59270 4406 59322
rect 4406 59270 4436 59322
rect 4460 59270 4470 59322
rect 4470 59270 4516 59322
rect 4220 59268 4276 59270
rect 4300 59268 4356 59270
rect 4380 59268 4436 59270
rect 4460 59268 4516 59270
rect 34940 59322 34996 59324
rect 35020 59322 35076 59324
rect 35100 59322 35156 59324
rect 35180 59322 35236 59324
rect 34940 59270 34986 59322
rect 34986 59270 34996 59322
rect 35020 59270 35050 59322
rect 35050 59270 35062 59322
rect 35062 59270 35076 59322
rect 35100 59270 35114 59322
rect 35114 59270 35126 59322
rect 35126 59270 35156 59322
rect 35180 59270 35190 59322
rect 35190 59270 35236 59322
rect 34940 59268 34996 59270
rect 35020 59268 35076 59270
rect 35100 59268 35156 59270
rect 35180 59268 35236 59270
rect 19580 58778 19636 58780
rect 19660 58778 19716 58780
rect 19740 58778 19796 58780
rect 19820 58778 19876 58780
rect 19580 58726 19626 58778
rect 19626 58726 19636 58778
rect 19660 58726 19690 58778
rect 19690 58726 19702 58778
rect 19702 58726 19716 58778
rect 19740 58726 19754 58778
rect 19754 58726 19766 58778
rect 19766 58726 19796 58778
rect 19820 58726 19830 58778
rect 19830 58726 19876 58778
rect 19580 58724 19636 58726
rect 19660 58724 19716 58726
rect 19740 58724 19796 58726
rect 19820 58724 19876 58726
rect 50300 58778 50356 58780
rect 50380 58778 50436 58780
rect 50460 58778 50516 58780
rect 50540 58778 50596 58780
rect 50300 58726 50346 58778
rect 50346 58726 50356 58778
rect 50380 58726 50410 58778
rect 50410 58726 50422 58778
rect 50422 58726 50436 58778
rect 50460 58726 50474 58778
rect 50474 58726 50486 58778
rect 50486 58726 50516 58778
rect 50540 58726 50550 58778
rect 50550 58726 50596 58778
rect 50300 58724 50356 58726
rect 50380 58724 50436 58726
rect 50460 58724 50516 58726
rect 50540 58724 50596 58726
rect 4220 58234 4276 58236
rect 4300 58234 4356 58236
rect 4380 58234 4436 58236
rect 4460 58234 4516 58236
rect 4220 58182 4266 58234
rect 4266 58182 4276 58234
rect 4300 58182 4330 58234
rect 4330 58182 4342 58234
rect 4342 58182 4356 58234
rect 4380 58182 4394 58234
rect 4394 58182 4406 58234
rect 4406 58182 4436 58234
rect 4460 58182 4470 58234
rect 4470 58182 4516 58234
rect 4220 58180 4276 58182
rect 4300 58180 4356 58182
rect 4380 58180 4436 58182
rect 4460 58180 4516 58182
rect 34940 58234 34996 58236
rect 35020 58234 35076 58236
rect 35100 58234 35156 58236
rect 35180 58234 35236 58236
rect 34940 58182 34986 58234
rect 34986 58182 34996 58234
rect 35020 58182 35050 58234
rect 35050 58182 35062 58234
rect 35062 58182 35076 58234
rect 35100 58182 35114 58234
rect 35114 58182 35126 58234
rect 35126 58182 35156 58234
rect 35180 58182 35190 58234
rect 35190 58182 35236 58234
rect 34940 58180 34996 58182
rect 35020 58180 35076 58182
rect 35100 58180 35156 58182
rect 35180 58180 35236 58182
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 1490 49816 1546 49872
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 1490 49172 1492 49192
rect 1492 49172 1544 49192
rect 1544 49172 1546 49192
rect 1490 49136 1546 49172
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 1490 48456 1546 48512
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 1490 47776 1546 47832
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 1490 47096 1546 47152
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 1490 46436 1546 46472
rect 1490 46416 1492 46436
rect 1492 46416 1544 46436
rect 1544 46416 1546 46436
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 1490 45772 1492 45792
rect 1492 45772 1544 45792
rect 1544 45772 1546 45792
rect 1490 45736 1546 45772
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 1490 45056 1546 45112
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 1490 44376 1546 44432
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 1490 43696 1546 43752
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 1490 43052 1492 43072
rect 1492 43052 1544 43072
rect 1544 43052 1546 43072
rect 1490 43016 1546 43052
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 1490 42336 1546 42392
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 1490 41656 1546 41712
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 1490 40996 1546 41032
rect 1490 40976 1492 40996
rect 1492 40976 1544 40996
rect 1544 40976 1546 40996
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 1490 40332 1492 40352
rect 1492 40332 1544 40352
rect 1544 40332 1546 40352
rect 1490 40296 1546 40332
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 1490 39616 1546 39672
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 1490 38936 1546 38992
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 1490 38256 1546 38312
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 1490 37612 1492 37632
rect 1492 37612 1544 37632
rect 1544 37612 1546 37632
rect 1490 37576 1546 37612
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 1490 36896 1546 36952
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 1490 36216 1546 36272
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 1490 35556 1546 35592
rect 1490 35536 1492 35556
rect 1492 35536 1544 35556
rect 1544 35536 1546 35556
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 1490 34892 1492 34912
rect 1492 34892 1544 34912
rect 1544 34892 1546 34912
rect 1490 34856 1546 34892
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 1490 34176 1546 34232
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 1490 33496 1546 33552
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 1490 32816 1546 32872
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 1490 32172 1492 32192
rect 1492 32172 1544 32192
rect 1544 32172 1546 32192
rect 1490 32136 1546 32172
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 1490 31456 1546 31512
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 1490 30776 1546 30832
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 1490 30116 1546 30152
rect 1490 30096 1492 30116
rect 1492 30096 1544 30116
rect 1544 30096 1546 30116
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 1490 29452 1492 29472
rect 1492 29452 1544 29472
rect 1544 29452 1546 29472
rect 1490 29416 1546 29452
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 1490 28736 1546 28792
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 1490 28056 1546 28112
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 1490 27376 1546 27432
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 1490 26732 1492 26752
rect 1492 26732 1544 26752
rect 1544 26732 1546 26752
rect 1490 26696 1546 26732
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 1490 26016 1546 26072
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 1490 25336 1546 25392
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 1490 24676 1546 24712
rect 1490 24656 1492 24676
rect 1492 24656 1544 24676
rect 1544 24656 1546 24676
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 1490 24012 1492 24032
rect 1492 24012 1544 24032
rect 1544 24012 1546 24032
rect 1490 23976 1546 24012
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 1490 23296 1546 23352
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 1490 22616 1546 22672
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 1490 21936 1546 21992
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 1490 21292 1492 21312
rect 1492 21292 1544 21312
rect 1544 21292 1546 21312
rect 1490 21256 1546 21292
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 1490 20576 1546 20632
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 1490 19896 1546 19952
rect 1490 19236 1546 19272
rect 1490 19216 1492 19236
rect 1492 19216 1544 19236
rect 1544 19216 1546 19236
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 1490 18572 1492 18592
rect 1492 18572 1544 18592
rect 1544 18572 1546 18592
rect 1490 18536 1546 18572
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1490 17856 1546 17912
rect 1490 17176 1546 17232
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 1490 16496 1546 16552
rect 1490 15852 1492 15872
rect 1492 15852 1544 15872
rect 1544 15852 1546 15872
rect 1490 15816 1546 15852
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1490 15136 1546 15192
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1490 14456 1546 14512
rect 1490 13796 1546 13832
rect 1490 13776 1492 13796
rect 1492 13776 1544 13796
rect 1544 13776 1546 13796
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 1490 13132 1492 13152
rect 1492 13132 1544 13152
rect 1544 13132 1546 13152
rect 1490 13096 1546 13132
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 1490 12416 1546 12472
rect 1490 11736 1546 11792
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1490 11056 1546 11112
rect 1490 10412 1492 10432
rect 1492 10412 1544 10432
rect 1544 10412 1546 10432
rect 1490 10376 1546 10412
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1490 9696 1546 9752
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 1490 9016 1546 9072
rect 1490 8356 1546 8392
rect 1490 8336 1492 8356
rect 1492 8336 1544 8356
rect 1544 8336 1546 8356
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 1490 7692 1492 7712
rect 1492 7692 1544 7712
rect 1544 7692 1546 7712
rect 1490 7656 1546 7692
rect 1490 6976 1546 7032
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1490 6296 1546 6352
rect 1490 5616 1546 5672
rect 1490 4972 1492 4992
rect 1492 4972 1544 4992
rect 1544 4972 1546 4992
rect 1490 4936 1546 4972
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 53378 2896 53434 2952
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 63774 61104 63830 61160
rect 65660 64762 65716 64764
rect 65740 64762 65796 64764
rect 65820 64762 65876 64764
rect 65900 64762 65956 64764
rect 65660 64710 65706 64762
rect 65706 64710 65716 64762
rect 65740 64710 65770 64762
rect 65770 64710 65782 64762
rect 65782 64710 65796 64762
rect 65820 64710 65834 64762
rect 65834 64710 65846 64762
rect 65846 64710 65876 64762
rect 65900 64710 65910 64762
rect 65910 64710 65956 64762
rect 65660 64708 65716 64710
rect 65740 64708 65796 64710
rect 65820 64708 65876 64710
rect 65900 64708 65956 64710
rect 65660 63674 65716 63676
rect 65740 63674 65796 63676
rect 65820 63674 65876 63676
rect 65900 63674 65956 63676
rect 65660 63622 65706 63674
rect 65706 63622 65716 63674
rect 65740 63622 65770 63674
rect 65770 63622 65782 63674
rect 65782 63622 65796 63674
rect 65820 63622 65834 63674
rect 65834 63622 65846 63674
rect 65846 63622 65876 63674
rect 65900 63622 65910 63674
rect 65910 63622 65956 63674
rect 65660 63620 65716 63622
rect 65740 63620 65796 63622
rect 65820 63620 65876 63622
rect 65900 63620 65956 63622
rect 65660 62586 65716 62588
rect 65740 62586 65796 62588
rect 65820 62586 65876 62588
rect 65900 62586 65956 62588
rect 65660 62534 65706 62586
rect 65706 62534 65716 62586
rect 65740 62534 65770 62586
rect 65770 62534 65782 62586
rect 65782 62534 65796 62586
rect 65820 62534 65834 62586
rect 65834 62534 65846 62586
rect 65846 62534 65876 62586
rect 65900 62534 65910 62586
rect 65910 62534 65956 62586
rect 65660 62532 65716 62534
rect 65740 62532 65796 62534
rect 65820 62532 65876 62534
rect 65900 62532 65956 62534
rect 63590 60052 63592 60072
rect 63592 60052 63644 60072
rect 63644 60052 63646 60072
rect 63590 60016 63646 60052
rect 63774 59880 63830 59936
rect 64786 59880 64842 59936
rect 64602 59472 64658 59528
rect 65660 61498 65716 61500
rect 65740 61498 65796 61500
rect 65820 61498 65876 61500
rect 65900 61498 65956 61500
rect 65660 61446 65706 61498
rect 65706 61446 65716 61498
rect 65740 61446 65770 61498
rect 65770 61446 65782 61498
rect 65782 61446 65796 61498
rect 65820 61446 65834 61498
rect 65834 61446 65846 61498
rect 65846 61446 65876 61498
rect 65900 61446 65910 61498
rect 65910 61446 65956 61498
rect 65660 61444 65716 61446
rect 65740 61444 65796 61446
rect 65820 61444 65876 61446
rect 65900 61444 65956 61446
rect 64970 3304 65026 3360
rect 65338 59608 65394 59664
rect 65660 60410 65716 60412
rect 65740 60410 65796 60412
rect 65820 60410 65876 60412
rect 65900 60410 65956 60412
rect 65660 60358 65706 60410
rect 65706 60358 65716 60410
rect 65740 60358 65770 60410
rect 65770 60358 65782 60410
rect 65782 60358 65796 60410
rect 65820 60358 65834 60410
rect 65834 60358 65846 60410
rect 65846 60358 65876 60410
rect 65900 60358 65910 60410
rect 65910 60358 65956 60410
rect 65660 60356 65716 60358
rect 65740 60356 65796 60358
rect 65820 60356 65876 60358
rect 65900 60356 65956 60358
rect 65614 60152 65670 60208
rect 65522 60016 65578 60072
rect 65706 59492 65762 59528
rect 65706 59472 65708 59492
rect 65708 59472 65760 59492
rect 65760 59472 65762 59492
rect 65660 59322 65716 59324
rect 65740 59322 65796 59324
rect 65820 59322 65876 59324
rect 65900 59322 65956 59324
rect 65660 59270 65706 59322
rect 65706 59270 65716 59322
rect 65740 59270 65770 59322
rect 65770 59270 65782 59322
rect 65782 59270 65796 59322
rect 65820 59270 65834 59322
rect 65834 59270 65846 59322
rect 65846 59270 65876 59322
rect 65900 59270 65910 59322
rect 65910 59270 65956 59322
rect 65660 59268 65716 59270
rect 65740 59268 65796 59270
rect 65820 59268 65876 59270
rect 65900 59268 65956 59270
rect 65660 58234 65716 58236
rect 65740 58234 65796 58236
rect 65820 58234 65876 58236
rect 65900 58234 65956 58236
rect 65660 58182 65706 58234
rect 65706 58182 65716 58234
rect 65740 58182 65770 58234
rect 65770 58182 65782 58234
rect 65782 58182 65796 58234
rect 65820 58182 65834 58234
rect 65834 58182 65846 58234
rect 65846 58182 65876 58234
rect 65900 58182 65910 58234
rect 65910 58182 65956 58234
rect 65660 58180 65716 58182
rect 65740 58180 65796 58182
rect 65820 58180 65876 58182
rect 65900 58180 65956 58182
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 65982 3168 66038 3224
rect 68098 60188 68100 60208
rect 68100 60188 68152 60208
rect 68152 60188 68154 60208
rect 68098 60152 68154 60188
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
rect 69294 3188 69350 3224
rect 69294 3168 69296 3188
rect 69296 3168 69348 3188
rect 69348 3168 69350 3188
rect 72054 3304 72110 3360
rect 78034 74976 78090 75032
rect 78126 74332 78128 74352
rect 78128 74332 78180 74352
rect 78180 74332 78182 74352
rect 78126 74296 78182 74332
rect 77850 73636 77906 73672
rect 77850 73616 77852 73636
rect 77852 73616 77904 73636
rect 77904 73616 77906 73636
rect 78034 72972 78036 72992
rect 78036 72972 78088 72992
rect 78088 72972 78090 72992
rect 78034 72936 78090 72972
rect 77850 72256 77906 72312
rect 78034 71576 78090 71632
rect 78034 70896 78090 70952
rect 77850 70252 77852 70272
rect 77852 70252 77904 70272
rect 77904 70252 77906 70272
rect 77850 70216 77906 70252
rect 78126 69536 78182 69592
rect 77942 68856 77998 68912
rect 77942 68176 77998 68232
rect 78126 67496 78182 67552
rect 77942 66816 77998 66872
rect 78126 66136 78182 66192
rect 78126 65492 78128 65512
rect 78128 65492 78180 65512
rect 78180 65492 78182 65512
rect 78126 65456 78182 65492
rect 77942 64776 77998 64832
rect 78126 64096 78182 64152
rect 77942 63416 77998 63472
rect 77942 62736 77998 62792
rect 78126 62056 78182 62112
rect 77942 61376 77998 61432
rect 78126 60696 78182 60752
rect 78126 60052 78128 60072
rect 78128 60052 78180 60072
rect 78180 60052 78182 60072
rect 78126 60016 78182 60052
rect 77942 59336 77998 59392
rect 78126 58656 78182 58712
rect 77942 57976 77998 58032
rect 77942 57296 77998 57352
rect 78126 56616 78182 56672
rect 77942 55936 77998 55992
rect 78126 55256 78182 55312
rect 77298 53216 77354 53272
rect 77574 52572 77576 52592
rect 77576 52572 77628 52592
rect 77628 52572 77630 52592
rect 77574 52536 77630 52572
rect 77298 51176 77354 51232
rect 77114 50496 77170 50552
rect 77390 49852 77392 49872
rect 77392 49852 77444 49872
rect 77444 49852 77446 49872
rect 77390 49816 77446 49852
rect 78126 54612 78128 54632
rect 78128 54612 78180 54632
rect 78180 54612 78182 54632
rect 78126 54576 78182 54612
rect 77942 53896 77998 53952
rect 77942 51892 77944 51912
rect 77944 51892 77996 51912
rect 77996 51892 77998 51912
rect 77942 51856 77998 51892
rect 78126 49172 78128 49192
rect 78128 49172 78180 49192
rect 78180 49172 78182 49192
rect 78126 49136 78182 49172
rect 77114 48456 77170 48512
rect 78034 47776 78090 47832
rect 77850 47096 77906 47152
rect 77850 46436 77906 46472
rect 77850 46416 77852 46436
rect 77852 46416 77904 46436
rect 77904 46416 77906 46436
rect 78034 45772 78036 45792
rect 78036 45772 78088 45792
rect 78088 45772 78090 45792
rect 78034 45736 78090 45772
rect 77850 45056 77906 45112
rect 78034 44376 78090 44432
rect 78034 43696 78090 43752
rect 77850 43052 77852 43072
rect 77852 43052 77904 43072
rect 77904 43052 77906 43072
rect 77850 43016 77906 43052
rect 78034 42336 78090 42392
rect 77850 41656 77906 41712
rect 77850 40996 77906 41032
rect 77850 40976 77852 40996
rect 77852 40976 77904 40996
rect 77904 40976 77906 40996
rect 78034 40332 78036 40352
rect 78036 40332 78088 40352
rect 78088 40332 78090 40352
rect 78034 40296 78090 40332
rect 77850 39616 77906 39672
rect 78034 38936 78090 38992
rect 78034 38256 78090 38312
rect 77850 37612 77852 37632
rect 77852 37612 77904 37632
rect 77904 37612 77906 37632
rect 77850 37576 77906 37612
rect 78034 36896 78090 36952
rect 77850 36216 77906 36272
rect 77850 35556 77906 35592
rect 77850 35536 77852 35556
rect 77852 35536 77904 35556
rect 77904 35536 77906 35556
rect 78034 34892 78036 34912
rect 78036 34892 78088 34912
rect 78088 34892 78090 34912
rect 78034 34856 78090 34892
rect 77850 34176 77906 34232
rect 78034 33496 78090 33552
rect 78034 32816 78090 32872
rect 77850 32172 77852 32192
rect 77852 32172 77904 32192
rect 77904 32172 77906 32192
rect 77850 32136 77906 32172
rect 78034 31456 78090 31512
rect 77850 30776 77906 30832
rect 77850 30116 77906 30152
rect 77850 30096 77852 30116
rect 77852 30096 77904 30116
rect 77904 30096 77906 30116
rect 78034 29452 78036 29472
rect 78036 29452 78088 29472
rect 78088 29452 78090 29472
rect 78034 29416 78090 29452
rect 77850 28736 77906 28792
rect 78034 28056 78090 28112
rect 78034 27376 78090 27432
rect 77850 26732 77852 26752
rect 77852 26732 77904 26752
rect 77904 26732 77906 26752
rect 77850 26696 77906 26732
rect 78034 26016 78090 26072
rect 77850 25336 77906 25392
rect 77850 24676 77906 24712
rect 77850 24656 77852 24676
rect 77852 24656 77904 24676
rect 77904 24656 77906 24676
rect 78034 24012 78036 24032
rect 78036 24012 78088 24032
rect 78088 24012 78090 24032
rect 78034 23976 78090 24012
rect 77850 23296 77906 23352
rect 78034 22616 78090 22672
rect 78034 21936 78090 21992
rect 77850 21292 77852 21312
rect 77852 21292 77904 21312
rect 77904 21292 77906 21312
rect 77850 21256 77906 21292
rect 78034 20576 78090 20632
rect 77850 19896 77906 19952
rect 77850 19216 77906 19272
rect 78034 18572 78036 18592
rect 78036 18572 78088 18592
rect 78088 18572 78090 18592
rect 78034 18536 78090 18572
rect 77850 17856 77906 17912
rect 78034 17176 78090 17232
rect 78034 16496 78090 16552
rect 77850 15852 77852 15872
rect 77852 15852 77904 15872
rect 77904 15852 77906 15872
rect 77850 15816 77906 15852
rect 78034 15136 78090 15192
rect 77850 14456 77906 14512
rect 77850 13776 77906 13832
rect 78034 13132 78036 13152
rect 78036 13132 78088 13152
rect 78088 13132 78090 13152
rect 78034 13096 78090 13132
rect 77850 12416 77906 12472
rect 78034 11736 78090 11792
rect 78034 11056 78090 11112
rect 77850 10412 77852 10432
rect 77852 10412 77904 10432
rect 77904 10412 77906 10432
rect 77850 10376 77906 10412
rect 78034 9696 78090 9752
rect 77850 9016 77906 9072
rect 77850 8356 77906 8392
rect 77850 8336 77852 8356
rect 77852 8336 77904 8356
rect 77904 8336 77906 8356
rect 78034 7692 78036 7712
rect 78036 7692 78088 7712
rect 78088 7692 78090 7712
rect 78034 7656 78090 7692
rect 77850 6976 77906 7032
rect 78034 6296 78090 6352
rect 78034 5616 78090 5672
rect 77850 4972 77852 4992
rect 77852 4972 77904 4992
rect 77904 4972 77906 4992
rect 77850 4936 77906 4972
rect 77114 2916 77170 2952
rect 77114 2896 77116 2916
rect 77116 2896 77168 2916
rect 77168 2896 77170 2916
<< metal3 >>
rect 4210 77824 4526 77825
rect 4210 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4526 77824
rect 4210 77759 4526 77760
rect 34930 77824 35246 77825
rect 34930 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35246 77824
rect 34930 77759 35246 77760
rect 65650 77824 65966 77825
rect 65650 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65966 77824
rect 65650 77759 65966 77760
rect 19570 77280 19886 77281
rect 19570 77216 19576 77280
rect 19640 77216 19656 77280
rect 19720 77216 19736 77280
rect 19800 77216 19816 77280
rect 19880 77216 19886 77280
rect 19570 77215 19886 77216
rect 50290 77280 50606 77281
rect 50290 77216 50296 77280
rect 50360 77216 50376 77280
rect 50440 77216 50456 77280
rect 50520 77216 50536 77280
rect 50600 77216 50606 77280
rect 50290 77215 50606 77216
rect 4210 76736 4526 76737
rect 4210 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4526 76736
rect 4210 76671 4526 76672
rect 34930 76736 35246 76737
rect 34930 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35246 76736
rect 34930 76671 35246 76672
rect 65650 76736 65966 76737
rect 65650 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65966 76736
rect 65650 76671 65966 76672
rect 19570 76192 19886 76193
rect 19570 76128 19576 76192
rect 19640 76128 19656 76192
rect 19720 76128 19736 76192
rect 19800 76128 19816 76192
rect 19880 76128 19886 76192
rect 19570 76127 19886 76128
rect 50290 76192 50606 76193
rect 50290 76128 50296 76192
rect 50360 76128 50376 76192
rect 50440 76128 50456 76192
rect 50520 76128 50536 76192
rect 50600 76128 50606 76192
rect 50290 76127 50606 76128
rect 4210 75648 4526 75649
rect 4210 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4526 75648
rect 4210 75583 4526 75584
rect 34930 75648 35246 75649
rect 34930 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35246 75648
rect 34930 75583 35246 75584
rect 65650 75648 65966 75649
rect 65650 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65966 75648
rect 65650 75583 65966 75584
rect 1669 75308 1735 75309
rect 1669 75306 1716 75308
rect 1624 75304 1716 75306
rect 1624 75248 1674 75304
rect 1624 75246 1716 75248
rect 1669 75244 1716 75246
rect 1780 75244 1786 75308
rect 1669 75243 1735 75244
rect 19570 75104 19886 75105
rect 0 75034 800 75064
rect 19570 75040 19576 75104
rect 19640 75040 19656 75104
rect 19720 75040 19736 75104
rect 19800 75040 19816 75104
rect 19880 75040 19886 75104
rect 19570 75039 19886 75040
rect 50290 75104 50606 75105
rect 50290 75040 50296 75104
rect 50360 75040 50376 75104
rect 50440 75040 50456 75104
rect 50520 75040 50536 75104
rect 50600 75040 50606 75104
rect 50290 75039 50606 75040
rect 1485 75034 1551 75037
rect 0 75032 1551 75034
rect 0 74976 1490 75032
rect 1546 74976 1551 75032
rect 0 74974 1551 74976
rect 0 74944 800 74974
rect 1485 74971 1551 74974
rect 78029 75034 78095 75037
rect 79200 75034 80000 75064
rect 78029 75032 80000 75034
rect 78029 74976 78034 75032
rect 78090 74976 80000 75032
rect 78029 74974 80000 74976
rect 78029 74971 78095 74974
rect 79200 74944 80000 74974
rect 4210 74560 4526 74561
rect 4210 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4526 74560
rect 4210 74495 4526 74496
rect 34930 74560 35246 74561
rect 34930 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35246 74560
rect 34930 74495 35246 74496
rect 65650 74560 65966 74561
rect 65650 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65966 74560
rect 65650 74495 65966 74496
rect 0 74354 800 74384
rect 1393 74354 1459 74357
rect 0 74352 1459 74354
rect 0 74296 1398 74352
rect 1454 74296 1459 74352
rect 0 74294 1459 74296
rect 0 74264 800 74294
rect 1393 74291 1459 74294
rect 78121 74354 78187 74357
rect 79200 74354 80000 74384
rect 78121 74352 80000 74354
rect 78121 74296 78126 74352
rect 78182 74296 80000 74352
rect 78121 74294 80000 74296
rect 78121 74291 78187 74294
rect 79200 74264 80000 74294
rect 19570 74016 19886 74017
rect 19570 73952 19576 74016
rect 19640 73952 19656 74016
rect 19720 73952 19736 74016
rect 19800 73952 19816 74016
rect 19880 73952 19886 74016
rect 19570 73951 19886 73952
rect 50290 74016 50606 74017
rect 50290 73952 50296 74016
rect 50360 73952 50376 74016
rect 50440 73952 50456 74016
rect 50520 73952 50536 74016
rect 50600 73952 50606 74016
rect 50290 73951 50606 73952
rect 0 73674 800 73704
rect 1485 73674 1551 73677
rect 0 73672 1551 73674
rect 0 73616 1490 73672
rect 1546 73616 1551 73672
rect 0 73614 1551 73616
rect 0 73584 800 73614
rect 1485 73611 1551 73614
rect 77845 73674 77911 73677
rect 79200 73674 80000 73704
rect 77845 73672 80000 73674
rect 77845 73616 77850 73672
rect 77906 73616 80000 73672
rect 77845 73614 80000 73616
rect 77845 73611 77911 73614
rect 79200 73584 80000 73614
rect 4210 73472 4526 73473
rect 4210 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4526 73472
rect 4210 73407 4526 73408
rect 34930 73472 35246 73473
rect 34930 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35246 73472
rect 34930 73407 35246 73408
rect 65650 73472 65966 73473
rect 65650 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65966 73472
rect 65650 73407 65966 73408
rect 0 72994 800 73024
rect 1485 72994 1551 72997
rect 0 72992 1551 72994
rect 0 72936 1490 72992
rect 1546 72936 1551 72992
rect 0 72934 1551 72936
rect 0 72904 800 72934
rect 1485 72931 1551 72934
rect 78029 72994 78095 72997
rect 79200 72994 80000 73024
rect 78029 72992 80000 72994
rect 78029 72936 78034 72992
rect 78090 72936 80000 72992
rect 78029 72934 80000 72936
rect 78029 72931 78095 72934
rect 19570 72928 19886 72929
rect 19570 72864 19576 72928
rect 19640 72864 19656 72928
rect 19720 72864 19736 72928
rect 19800 72864 19816 72928
rect 19880 72864 19886 72928
rect 19570 72863 19886 72864
rect 50290 72928 50606 72929
rect 50290 72864 50296 72928
rect 50360 72864 50376 72928
rect 50440 72864 50456 72928
rect 50520 72864 50536 72928
rect 50600 72864 50606 72928
rect 79200 72904 80000 72934
rect 50290 72863 50606 72864
rect 4210 72384 4526 72385
rect 0 72314 800 72344
rect 4210 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4526 72384
rect 4210 72319 4526 72320
rect 34930 72384 35246 72385
rect 34930 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35246 72384
rect 34930 72319 35246 72320
rect 65650 72384 65966 72385
rect 65650 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65966 72384
rect 65650 72319 65966 72320
rect 1485 72314 1551 72317
rect 0 72312 1551 72314
rect 0 72256 1490 72312
rect 1546 72256 1551 72312
rect 0 72254 1551 72256
rect 0 72224 800 72254
rect 1485 72251 1551 72254
rect 77845 72314 77911 72317
rect 79200 72314 80000 72344
rect 77845 72312 80000 72314
rect 77845 72256 77850 72312
rect 77906 72256 80000 72312
rect 77845 72254 80000 72256
rect 77845 72251 77911 72254
rect 79200 72224 80000 72254
rect 19570 71840 19886 71841
rect 19570 71776 19576 71840
rect 19640 71776 19656 71840
rect 19720 71776 19736 71840
rect 19800 71776 19816 71840
rect 19880 71776 19886 71840
rect 19570 71775 19886 71776
rect 50290 71840 50606 71841
rect 50290 71776 50296 71840
rect 50360 71776 50376 71840
rect 50440 71776 50456 71840
rect 50520 71776 50536 71840
rect 50600 71776 50606 71840
rect 50290 71775 50606 71776
rect 0 71634 800 71664
rect 1485 71634 1551 71637
rect 0 71632 1551 71634
rect 0 71576 1490 71632
rect 1546 71576 1551 71632
rect 0 71574 1551 71576
rect 0 71544 800 71574
rect 1485 71571 1551 71574
rect 78029 71634 78095 71637
rect 79200 71634 80000 71664
rect 78029 71632 80000 71634
rect 78029 71576 78034 71632
rect 78090 71576 80000 71632
rect 78029 71574 80000 71576
rect 78029 71571 78095 71574
rect 79200 71544 80000 71574
rect 4210 71296 4526 71297
rect 4210 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4526 71296
rect 4210 71231 4526 71232
rect 34930 71296 35246 71297
rect 34930 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35246 71296
rect 34930 71231 35246 71232
rect 65650 71296 65966 71297
rect 65650 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65966 71296
rect 65650 71231 65966 71232
rect 0 70954 800 70984
rect 1485 70954 1551 70957
rect 0 70952 1551 70954
rect 0 70896 1490 70952
rect 1546 70896 1551 70952
rect 0 70894 1551 70896
rect 0 70864 800 70894
rect 1485 70891 1551 70894
rect 78029 70954 78095 70957
rect 79200 70954 80000 70984
rect 78029 70952 80000 70954
rect 78029 70896 78034 70952
rect 78090 70896 80000 70952
rect 78029 70894 80000 70896
rect 78029 70891 78095 70894
rect 79200 70864 80000 70894
rect 19570 70752 19886 70753
rect 19570 70688 19576 70752
rect 19640 70688 19656 70752
rect 19720 70688 19736 70752
rect 19800 70688 19816 70752
rect 19880 70688 19886 70752
rect 19570 70687 19886 70688
rect 50290 70752 50606 70753
rect 50290 70688 50296 70752
rect 50360 70688 50376 70752
rect 50440 70688 50456 70752
rect 50520 70688 50536 70752
rect 50600 70688 50606 70752
rect 50290 70687 50606 70688
rect 0 70274 800 70304
rect 1485 70274 1551 70277
rect 0 70272 1551 70274
rect 0 70216 1490 70272
rect 1546 70216 1551 70272
rect 0 70214 1551 70216
rect 0 70184 800 70214
rect 1485 70211 1551 70214
rect 77845 70274 77911 70277
rect 79200 70274 80000 70304
rect 77845 70272 80000 70274
rect 77845 70216 77850 70272
rect 77906 70216 80000 70272
rect 77845 70214 80000 70216
rect 77845 70211 77911 70214
rect 4210 70208 4526 70209
rect 4210 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4526 70208
rect 4210 70143 4526 70144
rect 34930 70208 35246 70209
rect 34930 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35246 70208
rect 34930 70143 35246 70144
rect 65650 70208 65966 70209
rect 65650 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65966 70208
rect 79200 70184 80000 70214
rect 65650 70143 65966 70144
rect 19570 69664 19886 69665
rect 0 69594 800 69624
rect 19570 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19886 69664
rect 19570 69599 19886 69600
rect 50290 69664 50606 69665
rect 50290 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50606 69664
rect 50290 69599 50606 69600
rect 1393 69594 1459 69597
rect 0 69592 1459 69594
rect 0 69536 1398 69592
rect 1454 69536 1459 69592
rect 0 69534 1459 69536
rect 0 69504 800 69534
rect 1393 69531 1459 69534
rect 78121 69594 78187 69597
rect 79200 69594 80000 69624
rect 78121 69592 80000 69594
rect 78121 69536 78126 69592
rect 78182 69536 80000 69592
rect 78121 69534 80000 69536
rect 78121 69531 78187 69534
rect 79200 69504 80000 69534
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 34930 69120 35246 69121
rect 34930 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35246 69120
rect 34930 69055 35246 69056
rect 65650 69120 65966 69121
rect 65650 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65966 69120
rect 65650 69055 65966 69056
rect 0 68914 800 68944
rect 1393 68914 1459 68917
rect 0 68912 1459 68914
rect 0 68856 1398 68912
rect 1454 68856 1459 68912
rect 0 68854 1459 68856
rect 0 68824 800 68854
rect 1393 68851 1459 68854
rect 77937 68914 78003 68917
rect 79200 68914 80000 68944
rect 77937 68912 80000 68914
rect 77937 68856 77942 68912
rect 77998 68856 80000 68912
rect 77937 68854 80000 68856
rect 77937 68851 78003 68854
rect 79200 68824 80000 68854
rect 19570 68576 19886 68577
rect 19570 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19886 68576
rect 19570 68511 19886 68512
rect 50290 68576 50606 68577
rect 50290 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50606 68576
rect 50290 68511 50606 68512
rect 0 68234 800 68264
rect 1393 68234 1459 68237
rect 0 68232 1459 68234
rect 0 68176 1398 68232
rect 1454 68176 1459 68232
rect 0 68174 1459 68176
rect 0 68144 800 68174
rect 1393 68171 1459 68174
rect 77937 68234 78003 68237
rect 79200 68234 80000 68264
rect 77937 68232 80000 68234
rect 77937 68176 77942 68232
rect 77998 68176 80000 68232
rect 77937 68174 80000 68176
rect 77937 68171 78003 68174
rect 79200 68144 80000 68174
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 4210 67967 4526 67968
rect 34930 68032 35246 68033
rect 34930 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35246 68032
rect 34930 67967 35246 67968
rect 65650 68032 65966 68033
rect 65650 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65966 68032
rect 65650 67967 65966 67968
rect 0 67554 800 67584
rect 1393 67554 1459 67557
rect 0 67552 1459 67554
rect 0 67496 1398 67552
rect 1454 67496 1459 67552
rect 0 67494 1459 67496
rect 0 67464 800 67494
rect 1393 67491 1459 67494
rect 78121 67554 78187 67557
rect 79200 67554 80000 67584
rect 78121 67552 80000 67554
rect 78121 67496 78126 67552
rect 78182 67496 80000 67552
rect 78121 67494 80000 67496
rect 78121 67491 78187 67494
rect 19570 67488 19886 67489
rect 19570 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19886 67488
rect 19570 67423 19886 67424
rect 50290 67488 50606 67489
rect 50290 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50606 67488
rect 79200 67464 80000 67494
rect 50290 67423 50606 67424
rect 4210 66944 4526 66945
rect 0 66874 800 66904
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 34930 66944 35246 66945
rect 34930 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35246 66944
rect 34930 66879 35246 66880
rect 65650 66944 65966 66945
rect 65650 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65966 66944
rect 65650 66879 65966 66880
rect 1393 66874 1459 66877
rect 0 66872 1459 66874
rect 0 66816 1398 66872
rect 1454 66816 1459 66872
rect 0 66814 1459 66816
rect 0 66784 800 66814
rect 1393 66811 1459 66814
rect 77937 66874 78003 66877
rect 79200 66874 80000 66904
rect 77937 66872 80000 66874
rect 77937 66816 77942 66872
rect 77998 66816 80000 66872
rect 77937 66814 80000 66816
rect 77937 66811 78003 66814
rect 79200 66784 80000 66814
rect 19570 66400 19886 66401
rect 19570 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19886 66400
rect 19570 66335 19886 66336
rect 50290 66400 50606 66401
rect 50290 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50606 66400
rect 50290 66335 50606 66336
rect 0 66194 800 66224
rect 1393 66194 1459 66197
rect 0 66192 1459 66194
rect 0 66136 1398 66192
rect 1454 66136 1459 66192
rect 0 66134 1459 66136
rect 0 66104 800 66134
rect 1393 66131 1459 66134
rect 78121 66194 78187 66197
rect 79200 66194 80000 66224
rect 78121 66192 80000 66194
rect 78121 66136 78126 66192
rect 78182 66136 80000 66192
rect 78121 66134 80000 66136
rect 78121 66131 78187 66134
rect 79200 66104 80000 66134
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 34930 65856 35246 65857
rect 34930 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35246 65856
rect 34930 65791 35246 65792
rect 65650 65856 65966 65857
rect 65650 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65966 65856
rect 65650 65791 65966 65792
rect 0 65514 800 65544
rect 1393 65514 1459 65517
rect 0 65512 1459 65514
rect 0 65456 1398 65512
rect 1454 65456 1459 65512
rect 0 65454 1459 65456
rect 0 65424 800 65454
rect 1393 65451 1459 65454
rect 78121 65514 78187 65517
rect 79200 65514 80000 65544
rect 78121 65512 80000 65514
rect 78121 65456 78126 65512
rect 78182 65456 80000 65512
rect 78121 65454 80000 65456
rect 78121 65451 78187 65454
rect 79200 65424 80000 65454
rect 19570 65312 19886 65313
rect 19570 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19886 65312
rect 19570 65247 19886 65248
rect 50290 65312 50606 65313
rect 50290 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50606 65312
rect 50290 65247 50606 65248
rect 0 64834 800 64864
rect 1393 64834 1459 64837
rect 0 64832 1459 64834
rect 0 64776 1398 64832
rect 1454 64776 1459 64832
rect 0 64774 1459 64776
rect 0 64744 800 64774
rect 1393 64771 1459 64774
rect 77937 64834 78003 64837
rect 79200 64834 80000 64864
rect 77937 64832 80000 64834
rect 77937 64776 77942 64832
rect 77998 64776 80000 64832
rect 77937 64774 80000 64776
rect 77937 64771 78003 64774
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 34930 64768 35246 64769
rect 34930 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35246 64768
rect 34930 64703 35246 64704
rect 65650 64768 65966 64769
rect 65650 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65966 64768
rect 79200 64744 80000 64774
rect 65650 64703 65966 64704
rect 19570 64224 19886 64225
rect 0 64154 800 64184
rect 19570 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19886 64224
rect 19570 64159 19886 64160
rect 50290 64224 50606 64225
rect 50290 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50606 64224
rect 50290 64159 50606 64160
rect 1393 64154 1459 64157
rect 0 64152 1459 64154
rect 0 64096 1398 64152
rect 1454 64096 1459 64152
rect 0 64094 1459 64096
rect 0 64064 800 64094
rect 1393 64091 1459 64094
rect 78121 64154 78187 64157
rect 79200 64154 80000 64184
rect 78121 64152 80000 64154
rect 78121 64096 78126 64152
rect 78182 64096 80000 64152
rect 78121 64094 80000 64096
rect 78121 64091 78187 64094
rect 79200 64064 80000 64094
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 34930 63680 35246 63681
rect 34930 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35246 63680
rect 34930 63615 35246 63616
rect 65650 63680 65966 63681
rect 65650 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65966 63680
rect 65650 63615 65966 63616
rect 0 63474 800 63504
rect 1393 63474 1459 63477
rect 0 63472 1459 63474
rect 0 63416 1398 63472
rect 1454 63416 1459 63472
rect 0 63414 1459 63416
rect 0 63384 800 63414
rect 1393 63411 1459 63414
rect 77937 63474 78003 63477
rect 79200 63474 80000 63504
rect 77937 63472 80000 63474
rect 77937 63416 77942 63472
rect 77998 63416 80000 63472
rect 77937 63414 80000 63416
rect 77937 63411 78003 63414
rect 79200 63384 80000 63414
rect 19570 63136 19886 63137
rect 19570 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19886 63136
rect 19570 63071 19886 63072
rect 50290 63136 50606 63137
rect 50290 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50606 63136
rect 50290 63071 50606 63072
rect 0 62794 800 62824
rect 1393 62794 1459 62797
rect 0 62792 1459 62794
rect 0 62736 1398 62792
rect 1454 62736 1459 62792
rect 0 62734 1459 62736
rect 0 62704 800 62734
rect 1393 62731 1459 62734
rect 77937 62794 78003 62797
rect 79200 62794 80000 62824
rect 77937 62792 80000 62794
rect 77937 62736 77942 62792
rect 77998 62736 80000 62792
rect 77937 62734 80000 62736
rect 77937 62731 78003 62734
rect 79200 62704 80000 62734
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 34930 62592 35246 62593
rect 34930 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35246 62592
rect 34930 62527 35246 62528
rect 65650 62592 65966 62593
rect 65650 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65966 62592
rect 65650 62527 65966 62528
rect 0 62114 800 62144
rect 1393 62114 1459 62117
rect 0 62112 1459 62114
rect 0 62056 1398 62112
rect 1454 62056 1459 62112
rect 0 62054 1459 62056
rect 0 62024 800 62054
rect 1393 62051 1459 62054
rect 78121 62114 78187 62117
rect 79200 62114 80000 62144
rect 78121 62112 80000 62114
rect 78121 62056 78126 62112
rect 78182 62056 80000 62112
rect 78121 62054 80000 62056
rect 78121 62051 78187 62054
rect 19570 62048 19886 62049
rect 19570 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19886 62048
rect 19570 61983 19886 61984
rect 50290 62048 50606 62049
rect 50290 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50606 62048
rect 79200 62024 80000 62054
rect 50290 61983 50606 61984
rect 4210 61504 4526 61505
rect 0 61434 800 61464
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 34930 61504 35246 61505
rect 34930 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35246 61504
rect 34930 61439 35246 61440
rect 65650 61504 65966 61505
rect 65650 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65966 61504
rect 65650 61439 65966 61440
rect 1393 61434 1459 61437
rect 0 61432 1459 61434
rect 0 61376 1398 61432
rect 1454 61376 1459 61432
rect 0 61374 1459 61376
rect 0 61344 800 61374
rect 1393 61371 1459 61374
rect 77937 61434 78003 61437
rect 79200 61434 80000 61464
rect 77937 61432 80000 61434
rect 77937 61376 77942 61432
rect 77998 61376 80000 61432
rect 77937 61374 80000 61376
rect 77937 61371 78003 61374
rect 79200 61344 80000 61374
rect 1710 61100 1716 61164
rect 1780 61162 1786 61164
rect 63769 61162 63835 61165
rect 1780 61160 63835 61162
rect 1780 61104 63774 61160
rect 63830 61104 63835 61160
rect 1780 61102 63835 61104
rect 1780 61100 1786 61102
rect 63769 61099 63835 61102
rect 19570 60960 19886 60961
rect 19570 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19886 60960
rect 19570 60895 19886 60896
rect 50290 60960 50606 60961
rect 50290 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50606 60960
rect 50290 60895 50606 60896
rect 0 60754 800 60784
rect 1393 60754 1459 60757
rect 0 60752 1459 60754
rect 0 60696 1398 60752
rect 1454 60696 1459 60752
rect 0 60694 1459 60696
rect 0 60664 800 60694
rect 1393 60691 1459 60694
rect 78121 60754 78187 60757
rect 79200 60754 80000 60784
rect 78121 60752 80000 60754
rect 78121 60696 78126 60752
rect 78182 60696 80000 60752
rect 78121 60694 80000 60696
rect 78121 60691 78187 60694
rect 79200 60664 80000 60694
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 34930 60416 35246 60417
rect 34930 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35246 60416
rect 34930 60351 35246 60352
rect 65650 60416 65966 60417
rect 65650 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65966 60416
rect 65650 60351 65966 60352
rect 1669 60210 1735 60213
rect 65609 60210 65675 60213
rect 68093 60210 68159 60213
rect 1669 60208 68159 60210
rect 1669 60152 1674 60208
rect 1730 60152 65614 60208
rect 65670 60152 68098 60208
rect 68154 60152 68159 60208
rect 1669 60150 68159 60152
rect 1669 60147 1735 60150
rect 65609 60147 65675 60150
rect 68093 60147 68159 60150
rect 0 60074 800 60104
rect 1393 60074 1459 60077
rect 0 60072 1459 60074
rect 0 60016 1398 60072
rect 1454 60016 1459 60072
rect 0 60014 1459 60016
rect 0 59984 800 60014
rect 1393 60011 1459 60014
rect 63585 60074 63651 60077
rect 65517 60074 65583 60077
rect 63585 60072 65583 60074
rect 63585 60016 63590 60072
rect 63646 60016 65522 60072
rect 65578 60016 65583 60072
rect 63585 60014 65583 60016
rect 63585 60011 63651 60014
rect 65517 60011 65583 60014
rect 78121 60074 78187 60077
rect 79200 60074 80000 60104
rect 78121 60072 80000 60074
rect 78121 60016 78126 60072
rect 78182 60016 80000 60072
rect 78121 60014 80000 60016
rect 78121 60011 78187 60014
rect 79200 59984 80000 60014
rect 63769 59938 63835 59941
rect 64781 59938 64847 59941
rect 63769 59936 64847 59938
rect 63769 59880 63774 59936
rect 63830 59880 64786 59936
rect 64842 59880 64847 59936
rect 63769 59878 64847 59880
rect 63769 59875 63835 59878
rect 64781 59875 64847 59878
rect 19570 59872 19886 59873
rect 19570 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19886 59872
rect 19570 59807 19886 59808
rect 50290 59872 50606 59873
rect 50290 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50606 59872
rect 50290 59807 50606 59808
rect 1853 59666 1919 59669
rect 65333 59666 65399 59669
rect 1853 59664 65399 59666
rect 1853 59608 1858 59664
rect 1914 59608 65338 59664
rect 65394 59608 65399 59664
rect 1853 59606 65399 59608
rect 1853 59603 1919 59606
rect 65333 59603 65399 59606
rect 64597 59530 64663 59533
rect 65701 59530 65767 59533
rect 64597 59528 65767 59530
rect 64597 59472 64602 59528
rect 64658 59472 65706 59528
rect 65762 59472 65767 59528
rect 64597 59470 65767 59472
rect 64597 59467 64663 59470
rect 65701 59467 65767 59470
rect 0 59394 800 59424
rect 1393 59394 1459 59397
rect 0 59392 1459 59394
rect 0 59336 1398 59392
rect 1454 59336 1459 59392
rect 0 59334 1459 59336
rect 0 59304 800 59334
rect 1393 59331 1459 59334
rect 77937 59394 78003 59397
rect 79200 59394 80000 59424
rect 77937 59392 80000 59394
rect 77937 59336 77942 59392
rect 77998 59336 80000 59392
rect 77937 59334 80000 59336
rect 77937 59331 78003 59334
rect 4210 59328 4526 59329
rect 4210 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4526 59328
rect 4210 59263 4526 59264
rect 34930 59328 35246 59329
rect 34930 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35246 59328
rect 34930 59263 35246 59264
rect 65650 59328 65966 59329
rect 65650 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65966 59328
rect 79200 59304 80000 59334
rect 65650 59263 65966 59264
rect 19570 58784 19886 58785
rect 0 58714 800 58744
rect 19570 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19886 58784
rect 19570 58719 19886 58720
rect 50290 58784 50606 58785
rect 50290 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50606 58784
rect 50290 58719 50606 58720
rect 1393 58714 1459 58717
rect 0 58712 1459 58714
rect 0 58656 1398 58712
rect 1454 58656 1459 58712
rect 0 58654 1459 58656
rect 0 58624 800 58654
rect 1393 58651 1459 58654
rect 78121 58714 78187 58717
rect 79200 58714 80000 58744
rect 78121 58712 80000 58714
rect 78121 58656 78126 58712
rect 78182 58656 80000 58712
rect 78121 58654 80000 58656
rect 78121 58651 78187 58654
rect 79200 58624 80000 58654
rect 4210 58240 4526 58241
rect 4210 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4526 58240
rect 4210 58175 4526 58176
rect 34930 58240 35246 58241
rect 34930 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35246 58240
rect 34930 58175 35246 58176
rect 65650 58240 65966 58241
rect 65650 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65966 58240
rect 65650 58175 65966 58176
rect 0 58034 800 58064
rect 1393 58034 1459 58037
rect 0 58032 1459 58034
rect 0 57976 1398 58032
rect 1454 57976 1459 58032
rect 0 57974 1459 57976
rect 0 57944 800 57974
rect 1393 57971 1459 57974
rect 77937 58034 78003 58037
rect 79200 58034 80000 58064
rect 77937 58032 80000 58034
rect 77937 57976 77942 58032
rect 77998 57976 80000 58032
rect 77937 57974 80000 57976
rect 77937 57971 78003 57974
rect 79200 57944 80000 57974
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 0 57354 800 57384
rect 1393 57354 1459 57357
rect 0 57352 1459 57354
rect 0 57296 1398 57352
rect 1454 57296 1459 57352
rect 0 57294 1459 57296
rect 0 57264 800 57294
rect 1393 57291 1459 57294
rect 77937 57354 78003 57357
rect 79200 57354 80000 57384
rect 77937 57352 80000 57354
rect 77937 57296 77942 57352
rect 77998 57296 80000 57352
rect 77937 57294 80000 57296
rect 77937 57291 78003 57294
rect 79200 57264 80000 57294
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 65650 57152 65966 57153
rect 65650 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65966 57152
rect 65650 57087 65966 57088
rect 0 56674 800 56704
rect 1393 56674 1459 56677
rect 0 56672 1459 56674
rect 0 56616 1398 56672
rect 1454 56616 1459 56672
rect 0 56614 1459 56616
rect 0 56584 800 56614
rect 1393 56611 1459 56614
rect 78121 56674 78187 56677
rect 79200 56674 80000 56704
rect 78121 56672 80000 56674
rect 78121 56616 78126 56672
rect 78182 56616 80000 56672
rect 78121 56614 80000 56616
rect 78121 56611 78187 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 79200 56584 80000 56614
rect 50290 56543 50606 56544
rect 4210 56064 4526 56065
rect 0 55994 800 56024
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 65650 56064 65966 56065
rect 65650 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65966 56064
rect 65650 55999 65966 56000
rect 1393 55994 1459 55997
rect 0 55992 1459 55994
rect 0 55936 1398 55992
rect 1454 55936 1459 55992
rect 0 55934 1459 55936
rect 0 55904 800 55934
rect 1393 55931 1459 55934
rect 77937 55994 78003 55997
rect 79200 55994 80000 56024
rect 77937 55992 80000 55994
rect 77937 55936 77942 55992
rect 77998 55936 80000 55992
rect 77937 55934 80000 55936
rect 77937 55931 78003 55934
rect 79200 55904 80000 55934
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 0 55314 800 55344
rect 1485 55314 1551 55317
rect 0 55312 1551 55314
rect 0 55256 1490 55312
rect 1546 55256 1551 55312
rect 0 55254 1551 55256
rect 0 55224 800 55254
rect 1485 55251 1551 55254
rect 78121 55314 78187 55317
rect 79200 55314 80000 55344
rect 78121 55312 80000 55314
rect 78121 55256 78126 55312
rect 78182 55256 80000 55312
rect 78121 55254 80000 55256
rect 78121 55251 78187 55254
rect 79200 55224 80000 55254
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 65650 54976 65966 54977
rect 65650 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65966 54976
rect 65650 54911 65966 54912
rect 0 54634 800 54664
rect 1485 54634 1551 54637
rect 0 54632 1551 54634
rect 0 54576 1490 54632
rect 1546 54576 1551 54632
rect 0 54574 1551 54576
rect 0 54544 800 54574
rect 1485 54571 1551 54574
rect 78121 54634 78187 54637
rect 79200 54634 80000 54664
rect 78121 54632 80000 54634
rect 78121 54576 78126 54632
rect 78182 54576 80000 54632
rect 78121 54574 80000 54576
rect 78121 54571 78187 54574
rect 79200 54544 80000 54574
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 0 53954 800 53984
rect 1485 53954 1551 53957
rect 0 53952 1551 53954
rect 0 53896 1490 53952
rect 1546 53896 1551 53952
rect 0 53894 1551 53896
rect 0 53864 800 53894
rect 1485 53891 1551 53894
rect 77937 53954 78003 53957
rect 79200 53954 80000 53984
rect 77937 53952 80000 53954
rect 77937 53896 77942 53952
rect 77998 53896 80000 53952
rect 77937 53894 80000 53896
rect 77937 53891 78003 53894
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 65650 53888 65966 53889
rect 65650 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65966 53888
rect 79200 53864 80000 53894
rect 65650 53823 65966 53824
rect 19570 53344 19886 53345
rect 0 53274 800 53304
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 1485 53274 1551 53277
rect 0 53272 1551 53274
rect 0 53216 1490 53272
rect 1546 53216 1551 53272
rect 0 53214 1551 53216
rect 0 53184 800 53214
rect 1485 53211 1551 53214
rect 77293 53274 77359 53277
rect 79200 53274 80000 53304
rect 77293 53272 80000 53274
rect 77293 53216 77298 53272
rect 77354 53216 80000 53272
rect 77293 53214 80000 53216
rect 77293 53211 77359 53214
rect 79200 53184 80000 53214
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 65650 52800 65966 52801
rect 65650 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65966 52800
rect 65650 52735 65966 52736
rect 0 52594 800 52624
rect 1485 52594 1551 52597
rect 0 52592 1551 52594
rect 0 52536 1490 52592
rect 1546 52536 1551 52592
rect 0 52534 1551 52536
rect 0 52504 800 52534
rect 1485 52531 1551 52534
rect 77569 52594 77635 52597
rect 79200 52594 80000 52624
rect 77569 52592 80000 52594
rect 77569 52536 77574 52592
rect 77630 52536 80000 52592
rect 77569 52534 80000 52536
rect 77569 52531 77635 52534
rect 79200 52504 80000 52534
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 0 51914 800 51944
rect 1485 51914 1551 51917
rect 0 51912 1551 51914
rect 0 51856 1490 51912
rect 1546 51856 1551 51912
rect 0 51854 1551 51856
rect 0 51824 800 51854
rect 1485 51851 1551 51854
rect 77937 51914 78003 51917
rect 79200 51914 80000 51944
rect 77937 51912 80000 51914
rect 77937 51856 77942 51912
rect 77998 51856 80000 51912
rect 77937 51854 80000 51856
rect 77937 51851 78003 51854
rect 79200 51824 80000 51854
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 65650 51712 65966 51713
rect 65650 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65966 51712
rect 65650 51647 65966 51648
rect 0 51234 800 51264
rect 1485 51234 1551 51237
rect 0 51232 1551 51234
rect 0 51176 1490 51232
rect 1546 51176 1551 51232
rect 0 51174 1551 51176
rect 0 51144 800 51174
rect 1485 51171 1551 51174
rect 77293 51234 77359 51237
rect 79200 51234 80000 51264
rect 77293 51232 80000 51234
rect 77293 51176 77298 51232
rect 77354 51176 80000 51232
rect 77293 51174 80000 51176
rect 77293 51171 77359 51174
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 79200 51144 80000 51174
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 0 50554 800 50584
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 65650 50624 65966 50625
rect 65650 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65966 50624
rect 65650 50559 65966 50560
rect 1485 50554 1551 50557
rect 0 50552 1551 50554
rect 0 50496 1490 50552
rect 1546 50496 1551 50552
rect 0 50494 1551 50496
rect 0 50464 800 50494
rect 1485 50491 1551 50494
rect 77109 50554 77175 50557
rect 79200 50554 80000 50584
rect 77109 50552 80000 50554
rect 77109 50496 77114 50552
rect 77170 50496 80000 50552
rect 77109 50494 80000 50496
rect 77109 50491 77175 50494
rect 79200 50464 80000 50494
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 0 49874 800 49904
rect 1485 49874 1551 49877
rect 0 49872 1551 49874
rect 0 49816 1490 49872
rect 1546 49816 1551 49872
rect 0 49814 1551 49816
rect 0 49784 800 49814
rect 1485 49811 1551 49814
rect 77385 49874 77451 49877
rect 79200 49874 80000 49904
rect 77385 49872 80000 49874
rect 77385 49816 77390 49872
rect 77446 49816 80000 49872
rect 77385 49814 80000 49816
rect 77385 49811 77451 49814
rect 79200 49784 80000 49814
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 65650 49536 65966 49537
rect 65650 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65966 49536
rect 65650 49471 65966 49472
rect 0 49194 800 49224
rect 1485 49194 1551 49197
rect 0 49192 1551 49194
rect 0 49136 1490 49192
rect 1546 49136 1551 49192
rect 0 49134 1551 49136
rect 0 49104 800 49134
rect 1485 49131 1551 49134
rect 78121 49194 78187 49197
rect 79200 49194 80000 49224
rect 78121 49192 80000 49194
rect 78121 49136 78126 49192
rect 78182 49136 80000 49192
rect 78121 49134 80000 49136
rect 78121 49131 78187 49134
rect 79200 49104 80000 49134
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 0 48514 800 48544
rect 1485 48514 1551 48517
rect 0 48512 1551 48514
rect 0 48456 1490 48512
rect 1546 48456 1551 48512
rect 0 48454 1551 48456
rect 0 48424 800 48454
rect 1485 48451 1551 48454
rect 77109 48514 77175 48517
rect 79200 48514 80000 48544
rect 77109 48512 80000 48514
rect 77109 48456 77114 48512
rect 77170 48456 80000 48512
rect 77109 48454 80000 48456
rect 77109 48451 77175 48454
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 65650 48448 65966 48449
rect 65650 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65966 48448
rect 79200 48424 80000 48454
rect 65650 48383 65966 48384
rect 19570 47904 19886 47905
rect 0 47834 800 47864
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 1485 47834 1551 47837
rect 0 47832 1551 47834
rect 0 47776 1490 47832
rect 1546 47776 1551 47832
rect 0 47774 1551 47776
rect 0 47744 800 47774
rect 1485 47771 1551 47774
rect 78029 47834 78095 47837
rect 79200 47834 80000 47864
rect 78029 47832 80000 47834
rect 78029 47776 78034 47832
rect 78090 47776 80000 47832
rect 78029 47774 80000 47776
rect 78029 47771 78095 47774
rect 79200 47744 80000 47774
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 65650 47360 65966 47361
rect 65650 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65966 47360
rect 65650 47295 65966 47296
rect 0 47154 800 47184
rect 1485 47154 1551 47157
rect 0 47152 1551 47154
rect 0 47096 1490 47152
rect 1546 47096 1551 47152
rect 0 47094 1551 47096
rect 0 47064 800 47094
rect 1485 47091 1551 47094
rect 77845 47154 77911 47157
rect 79200 47154 80000 47184
rect 77845 47152 80000 47154
rect 77845 47096 77850 47152
rect 77906 47096 80000 47152
rect 77845 47094 80000 47096
rect 77845 47091 77911 47094
rect 79200 47064 80000 47094
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 0 46474 800 46504
rect 1485 46474 1551 46477
rect 0 46472 1551 46474
rect 0 46416 1490 46472
rect 1546 46416 1551 46472
rect 0 46414 1551 46416
rect 0 46384 800 46414
rect 1485 46411 1551 46414
rect 77845 46474 77911 46477
rect 79200 46474 80000 46504
rect 77845 46472 80000 46474
rect 77845 46416 77850 46472
rect 77906 46416 80000 46472
rect 77845 46414 80000 46416
rect 77845 46411 77911 46414
rect 79200 46384 80000 46414
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 65650 46272 65966 46273
rect 65650 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65966 46272
rect 65650 46207 65966 46208
rect 0 45794 800 45824
rect 1485 45794 1551 45797
rect 0 45792 1551 45794
rect 0 45736 1490 45792
rect 1546 45736 1551 45792
rect 0 45734 1551 45736
rect 0 45704 800 45734
rect 1485 45731 1551 45734
rect 78029 45794 78095 45797
rect 79200 45794 80000 45824
rect 78029 45792 80000 45794
rect 78029 45736 78034 45792
rect 78090 45736 80000 45792
rect 78029 45734 80000 45736
rect 78029 45731 78095 45734
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 79200 45704 80000 45734
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 0 45114 800 45144
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 65650 45184 65966 45185
rect 65650 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65966 45184
rect 65650 45119 65966 45120
rect 1485 45114 1551 45117
rect 0 45112 1551 45114
rect 0 45056 1490 45112
rect 1546 45056 1551 45112
rect 0 45054 1551 45056
rect 0 45024 800 45054
rect 1485 45051 1551 45054
rect 77845 45114 77911 45117
rect 79200 45114 80000 45144
rect 77845 45112 80000 45114
rect 77845 45056 77850 45112
rect 77906 45056 80000 45112
rect 77845 45054 80000 45056
rect 77845 45051 77911 45054
rect 79200 45024 80000 45054
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 0 44434 800 44464
rect 1485 44434 1551 44437
rect 0 44432 1551 44434
rect 0 44376 1490 44432
rect 1546 44376 1551 44432
rect 0 44374 1551 44376
rect 0 44344 800 44374
rect 1485 44371 1551 44374
rect 78029 44434 78095 44437
rect 79200 44434 80000 44464
rect 78029 44432 80000 44434
rect 78029 44376 78034 44432
rect 78090 44376 80000 44432
rect 78029 44374 80000 44376
rect 78029 44371 78095 44374
rect 79200 44344 80000 44374
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 65650 44096 65966 44097
rect 65650 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65966 44096
rect 65650 44031 65966 44032
rect 0 43754 800 43784
rect 1485 43754 1551 43757
rect 0 43752 1551 43754
rect 0 43696 1490 43752
rect 1546 43696 1551 43752
rect 0 43694 1551 43696
rect 0 43664 800 43694
rect 1485 43691 1551 43694
rect 78029 43754 78095 43757
rect 79200 43754 80000 43784
rect 78029 43752 80000 43754
rect 78029 43696 78034 43752
rect 78090 43696 80000 43752
rect 78029 43694 80000 43696
rect 78029 43691 78095 43694
rect 79200 43664 80000 43694
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 0 43074 800 43104
rect 1485 43074 1551 43077
rect 0 43072 1551 43074
rect 0 43016 1490 43072
rect 1546 43016 1551 43072
rect 0 43014 1551 43016
rect 0 42984 800 43014
rect 1485 43011 1551 43014
rect 77845 43074 77911 43077
rect 79200 43074 80000 43104
rect 77845 43072 80000 43074
rect 77845 43016 77850 43072
rect 77906 43016 80000 43072
rect 77845 43014 80000 43016
rect 77845 43011 77911 43014
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 65650 43008 65966 43009
rect 65650 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65966 43008
rect 79200 42984 80000 43014
rect 65650 42943 65966 42944
rect 19570 42464 19886 42465
rect 0 42394 800 42424
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 1485 42394 1551 42397
rect 0 42392 1551 42394
rect 0 42336 1490 42392
rect 1546 42336 1551 42392
rect 0 42334 1551 42336
rect 0 42304 800 42334
rect 1485 42331 1551 42334
rect 78029 42394 78095 42397
rect 79200 42394 80000 42424
rect 78029 42392 80000 42394
rect 78029 42336 78034 42392
rect 78090 42336 80000 42392
rect 78029 42334 80000 42336
rect 78029 42331 78095 42334
rect 79200 42304 80000 42334
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 65650 41920 65966 41921
rect 65650 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65966 41920
rect 65650 41855 65966 41856
rect 0 41714 800 41744
rect 1485 41714 1551 41717
rect 0 41712 1551 41714
rect 0 41656 1490 41712
rect 1546 41656 1551 41712
rect 0 41654 1551 41656
rect 0 41624 800 41654
rect 1485 41651 1551 41654
rect 77845 41714 77911 41717
rect 79200 41714 80000 41744
rect 77845 41712 80000 41714
rect 77845 41656 77850 41712
rect 77906 41656 80000 41712
rect 77845 41654 80000 41656
rect 77845 41651 77911 41654
rect 79200 41624 80000 41654
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 41034 800 41064
rect 1485 41034 1551 41037
rect 0 41032 1551 41034
rect 0 40976 1490 41032
rect 1546 40976 1551 41032
rect 0 40974 1551 40976
rect 0 40944 800 40974
rect 1485 40971 1551 40974
rect 77845 41034 77911 41037
rect 79200 41034 80000 41064
rect 77845 41032 80000 41034
rect 77845 40976 77850 41032
rect 77906 40976 80000 41032
rect 77845 40974 80000 40976
rect 77845 40971 77911 40974
rect 79200 40944 80000 40974
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 65650 40832 65966 40833
rect 65650 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65966 40832
rect 65650 40767 65966 40768
rect 0 40354 800 40384
rect 1485 40354 1551 40357
rect 0 40352 1551 40354
rect 0 40296 1490 40352
rect 1546 40296 1551 40352
rect 0 40294 1551 40296
rect 0 40264 800 40294
rect 1485 40291 1551 40294
rect 78029 40354 78095 40357
rect 79200 40354 80000 40384
rect 78029 40352 80000 40354
rect 78029 40296 78034 40352
rect 78090 40296 80000 40352
rect 78029 40294 80000 40296
rect 78029 40291 78095 40294
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 79200 40264 80000 40294
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 0 39674 800 39704
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 65650 39744 65966 39745
rect 65650 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65966 39744
rect 65650 39679 65966 39680
rect 1485 39674 1551 39677
rect 0 39672 1551 39674
rect 0 39616 1490 39672
rect 1546 39616 1551 39672
rect 0 39614 1551 39616
rect 0 39584 800 39614
rect 1485 39611 1551 39614
rect 77845 39674 77911 39677
rect 79200 39674 80000 39704
rect 77845 39672 80000 39674
rect 77845 39616 77850 39672
rect 77906 39616 80000 39672
rect 77845 39614 80000 39616
rect 77845 39611 77911 39614
rect 79200 39584 80000 39614
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 0 38994 800 39024
rect 1485 38994 1551 38997
rect 0 38992 1551 38994
rect 0 38936 1490 38992
rect 1546 38936 1551 38992
rect 0 38934 1551 38936
rect 0 38904 800 38934
rect 1485 38931 1551 38934
rect 78029 38994 78095 38997
rect 79200 38994 80000 39024
rect 78029 38992 80000 38994
rect 78029 38936 78034 38992
rect 78090 38936 80000 38992
rect 78029 38934 80000 38936
rect 78029 38931 78095 38934
rect 79200 38904 80000 38934
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 65650 38656 65966 38657
rect 65650 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65966 38656
rect 65650 38591 65966 38592
rect 0 38314 800 38344
rect 1485 38314 1551 38317
rect 0 38312 1551 38314
rect 0 38256 1490 38312
rect 1546 38256 1551 38312
rect 0 38254 1551 38256
rect 0 38224 800 38254
rect 1485 38251 1551 38254
rect 78029 38314 78095 38317
rect 79200 38314 80000 38344
rect 78029 38312 80000 38314
rect 78029 38256 78034 38312
rect 78090 38256 80000 38312
rect 78029 38254 80000 38256
rect 78029 38251 78095 38254
rect 79200 38224 80000 38254
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 0 37634 800 37664
rect 1485 37634 1551 37637
rect 0 37632 1551 37634
rect 0 37576 1490 37632
rect 1546 37576 1551 37632
rect 0 37574 1551 37576
rect 0 37544 800 37574
rect 1485 37571 1551 37574
rect 77845 37634 77911 37637
rect 79200 37634 80000 37664
rect 77845 37632 80000 37634
rect 77845 37576 77850 37632
rect 77906 37576 80000 37632
rect 77845 37574 80000 37576
rect 77845 37571 77911 37574
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 79200 37544 80000 37574
rect 65650 37503 65966 37504
rect 19570 37024 19886 37025
rect 0 36954 800 36984
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 1485 36954 1551 36957
rect 0 36952 1551 36954
rect 0 36896 1490 36952
rect 1546 36896 1551 36952
rect 0 36894 1551 36896
rect 0 36864 800 36894
rect 1485 36891 1551 36894
rect 78029 36954 78095 36957
rect 79200 36954 80000 36984
rect 78029 36952 80000 36954
rect 78029 36896 78034 36952
rect 78090 36896 80000 36952
rect 78029 36894 80000 36896
rect 78029 36891 78095 36894
rect 79200 36864 80000 36894
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 0 36274 800 36304
rect 1485 36274 1551 36277
rect 0 36272 1551 36274
rect 0 36216 1490 36272
rect 1546 36216 1551 36272
rect 0 36214 1551 36216
rect 0 36184 800 36214
rect 1485 36211 1551 36214
rect 77845 36274 77911 36277
rect 79200 36274 80000 36304
rect 77845 36272 80000 36274
rect 77845 36216 77850 36272
rect 77906 36216 80000 36272
rect 77845 36214 80000 36216
rect 77845 36211 77911 36214
rect 79200 36184 80000 36214
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 0 35594 800 35624
rect 1485 35594 1551 35597
rect 0 35592 1551 35594
rect 0 35536 1490 35592
rect 1546 35536 1551 35592
rect 0 35534 1551 35536
rect 0 35504 800 35534
rect 1485 35531 1551 35534
rect 77845 35594 77911 35597
rect 79200 35594 80000 35624
rect 77845 35592 80000 35594
rect 77845 35536 77850 35592
rect 77906 35536 80000 35592
rect 77845 35534 80000 35536
rect 77845 35531 77911 35534
rect 79200 35504 80000 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 0 34914 800 34944
rect 1485 34914 1551 34917
rect 0 34912 1551 34914
rect 0 34856 1490 34912
rect 1546 34856 1551 34912
rect 0 34854 1551 34856
rect 0 34824 800 34854
rect 1485 34851 1551 34854
rect 78029 34914 78095 34917
rect 79200 34914 80000 34944
rect 78029 34912 80000 34914
rect 78029 34856 78034 34912
rect 78090 34856 80000 34912
rect 78029 34854 80000 34856
rect 78029 34851 78095 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 79200 34824 80000 34854
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 0 34234 800 34264
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 1485 34234 1551 34237
rect 0 34232 1551 34234
rect 0 34176 1490 34232
rect 1546 34176 1551 34232
rect 0 34174 1551 34176
rect 0 34144 800 34174
rect 1485 34171 1551 34174
rect 77845 34234 77911 34237
rect 79200 34234 80000 34264
rect 77845 34232 80000 34234
rect 77845 34176 77850 34232
rect 77906 34176 80000 34232
rect 77845 34174 80000 34176
rect 77845 34171 77911 34174
rect 79200 34144 80000 34174
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 0 33554 800 33584
rect 1485 33554 1551 33557
rect 0 33552 1551 33554
rect 0 33496 1490 33552
rect 1546 33496 1551 33552
rect 0 33494 1551 33496
rect 0 33464 800 33494
rect 1485 33491 1551 33494
rect 78029 33554 78095 33557
rect 79200 33554 80000 33584
rect 78029 33552 80000 33554
rect 78029 33496 78034 33552
rect 78090 33496 80000 33552
rect 78029 33494 80000 33496
rect 78029 33491 78095 33494
rect 79200 33464 80000 33494
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 0 32874 800 32904
rect 1485 32874 1551 32877
rect 0 32872 1551 32874
rect 0 32816 1490 32872
rect 1546 32816 1551 32872
rect 0 32814 1551 32816
rect 0 32784 800 32814
rect 1485 32811 1551 32814
rect 78029 32874 78095 32877
rect 79200 32874 80000 32904
rect 78029 32872 80000 32874
rect 78029 32816 78034 32872
rect 78090 32816 80000 32872
rect 78029 32814 80000 32816
rect 78029 32811 78095 32814
rect 79200 32784 80000 32814
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 0 32194 800 32224
rect 1485 32194 1551 32197
rect 0 32192 1551 32194
rect 0 32136 1490 32192
rect 1546 32136 1551 32192
rect 0 32134 1551 32136
rect 0 32104 800 32134
rect 1485 32131 1551 32134
rect 77845 32194 77911 32197
rect 79200 32194 80000 32224
rect 77845 32192 80000 32194
rect 77845 32136 77850 32192
rect 77906 32136 80000 32192
rect 77845 32134 80000 32136
rect 77845 32131 77911 32134
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 79200 32104 80000 32134
rect 65650 32063 65966 32064
rect 19570 31584 19886 31585
rect 0 31514 800 31544
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 1485 31514 1551 31517
rect 0 31512 1551 31514
rect 0 31456 1490 31512
rect 1546 31456 1551 31512
rect 0 31454 1551 31456
rect 0 31424 800 31454
rect 1485 31451 1551 31454
rect 78029 31514 78095 31517
rect 79200 31514 80000 31544
rect 78029 31512 80000 31514
rect 78029 31456 78034 31512
rect 78090 31456 80000 31512
rect 78029 31454 80000 31456
rect 78029 31451 78095 31454
rect 79200 31424 80000 31454
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 0 30834 800 30864
rect 1485 30834 1551 30837
rect 0 30832 1551 30834
rect 0 30776 1490 30832
rect 1546 30776 1551 30832
rect 0 30774 1551 30776
rect 0 30744 800 30774
rect 1485 30771 1551 30774
rect 77845 30834 77911 30837
rect 79200 30834 80000 30864
rect 77845 30832 80000 30834
rect 77845 30776 77850 30832
rect 77906 30776 80000 30832
rect 77845 30774 80000 30776
rect 77845 30771 77911 30774
rect 79200 30744 80000 30774
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 0 30154 800 30184
rect 1485 30154 1551 30157
rect 0 30152 1551 30154
rect 0 30096 1490 30152
rect 1546 30096 1551 30152
rect 0 30094 1551 30096
rect 0 30064 800 30094
rect 1485 30091 1551 30094
rect 77845 30154 77911 30157
rect 79200 30154 80000 30184
rect 77845 30152 80000 30154
rect 77845 30096 77850 30152
rect 77906 30096 80000 30152
rect 77845 30094 80000 30096
rect 77845 30091 77911 30094
rect 79200 30064 80000 30094
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 0 29474 800 29504
rect 1485 29474 1551 29477
rect 0 29472 1551 29474
rect 0 29416 1490 29472
rect 1546 29416 1551 29472
rect 0 29414 1551 29416
rect 0 29384 800 29414
rect 1485 29411 1551 29414
rect 78029 29474 78095 29477
rect 79200 29474 80000 29504
rect 78029 29472 80000 29474
rect 78029 29416 78034 29472
rect 78090 29416 80000 29472
rect 78029 29414 80000 29416
rect 78029 29411 78095 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 79200 29384 80000 29414
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 0 28794 800 28824
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 1485 28794 1551 28797
rect 0 28792 1551 28794
rect 0 28736 1490 28792
rect 1546 28736 1551 28792
rect 0 28734 1551 28736
rect 0 28704 800 28734
rect 1485 28731 1551 28734
rect 77845 28794 77911 28797
rect 79200 28794 80000 28824
rect 77845 28792 80000 28794
rect 77845 28736 77850 28792
rect 77906 28736 80000 28792
rect 77845 28734 80000 28736
rect 77845 28731 77911 28734
rect 79200 28704 80000 28734
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 0 28114 800 28144
rect 1485 28114 1551 28117
rect 0 28112 1551 28114
rect 0 28056 1490 28112
rect 1546 28056 1551 28112
rect 0 28054 1551 28056
rect 0 28024 800 28054
rect 1485 28051 1551 28054
rect 78029 28114 78095 28117
rect 79200 28114 80000 28144
rect 78029 28112 80000 28114
rect 78029 28056 78034 28112
rect 78090 28056 80000 28112
rect 78029 28054 80000 28056
rect 78029 28051 78095 28054
rect 79200 28024 80000 28054
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 0 27434 800 27464
rect 1485 27434 1551 27437
rect 0 27432 1551 27434
rect 0 27376 1490 27432
rect 1546 27376 1551 27432
rect 0 27374 1551 27376
rect 0 27344 800 27374
rect 1485 27371 1551 27374
rect 78029 27434 78095 27437
rect 79200 27434 80000 27464
rect 78029 27432 80000 27434
rect 78029 27376 78034 27432
rect 78090 27376 80000 27432
rect 78029 27374 80000 27376
rect 78029 27371 78095 27374
rect 79200 27344 80000 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 0 26754 800 26784
rect 1485 26754 1551 26757
rect 0 26752 1551 26754
rect 0 26696 1490 26752
rect 1546 26696 1551 26752
rect 0 26694 1551 26696
rect 0 26664 800 26694
rect 1485 26691 1551 26694
rect 77845 26754 77911 26757
rect 79200 26754 80000 26784
rect 77845 26752 80000 26754
rect 77845 26696 77850 26752
rect 77906 26696 80000 26752
rect 77845 26694 80000 26696
rect 77845 26691 77911 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 79200 26664 80000 26694
rect 65650 26623 65966 26624
rect 19570 26144 19886 26145
rect 0 26074 800 26104
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 1485 26074 1551 26077
rect 0 26072 1551 26074
rect 0 26016 1490 26072
rect 1546 26016 1551 26072
rect 0 26014 1551 26016
rect 0 25984 800 26014
rect 1485 26011 1551 26014
rect 78029 26074 78095 26077
rect 79200 26074 80000 26104
rect 78029 26072 80000 26074
rect 78029 26016 78034 26072
rect 78090 26016 80000 26072
rect 78029 26014 80000 26016
rect 78029 26011 78095 26014
rect 79200 25984 80000 26014
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 0 25394 800 25424
rect 1485 25394 1551 25397
rect 0 25392 1551 25394
rect 0 25336 1490 25392
rect 1546 25336 1551 25392
rect 0 25334 1551 25336
rect 0 25304 800 25334
rect 1485 25331 1551 25334
rect 77845 25394 77911 25397
rect 79200 25394 80000 25424
rect 77845 25392 80000 25394
rect 77845 25336 77850 25392
rect 77906 25336 80000 25392
rect 77845 25334 80000 25336
rect 77845 25331 77911 25334
rect 79200 25304 80000 25334
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 0 24714 800 24744
rect 1485 24714 1551 24717
rect 0 24712 1551 24714
rect 0 24656 1490 24712
rect 1546 24656 1551 24712
rect 0 24654 1551 24656
rect 0 24624 800 24654
rect 1485 24651 1551 24654
rect 77845 24714 77911 24717
rect 79200 24714 80000 24744
rect 77845 24712 80000 24714
rect 77845 24656 77850 24712
rect 77906 24656 80000 24712
rect 77845 24654 80000 24656
rect 77845 24651 77911 24654
rect 79200 24624 80000 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 0 24034 800 24064
rect 1485 24034 1551 24037
rect 0 24032 1551 24034
rect 0 23976 1490 24032
rect 1546 23976 1551 24032
rect 0 23974 1551 23976
rect 0 23944 800 23974
rect 1485 23971 1551 23974
rect 78029 24034 78095 24037
rect 79200 24034 80000 24064
rect 78029 24032 80000 24034
rect 78029 23976 78034 24032
rect 78090 23976 80000 24032
rect 78029 23974 80000 23976
rect 78029 23971 78095 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 79200 23944 80000 23974
rect 50290 23903 50606 23904
rect 4210 23424 4526 23425
rect 0 23354 800 23384
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 1485 23354 1551 23357
rect 0 23352 1551 23354
rect 0 23296 1490 23352
rect 1546 23296 1551 23352
rect 0 23294 1551 23296
rect 0 23264 800 23294
rect 1485 23291 1551 23294
rect 77845 23354 77911 23357
rect 79200 23354 80000 23384
rect 77845 23352 80000 23354
rect 77845 23296 77850 23352
rect 77906 23296 80000 23352
rect 77845 23294 80000 23296
rect 77845 23291 77911 23294
rect 79200 23264 80000 23294
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 0 22674 800 22704
rect 1485 22674 1551 22677
rect 0 22672 1551 22674
rect 0 22616 1490 22672
rect 1546 22616 1551 22672
rect 0 22614 1551 22616
rect 0 22584 800 22614
rect 1485 22611 1551 22614
rect 78029 22674 78095 22677
rect 79200 22674 80000 22704
rect 78029 22672 80000 22674
rect 78029 22616 78034 22672
rect 78090 22616 80000 22672
rect 78029 22614 80000 22616
rect 78029 22611 78095 22614
rect 79200 22584 80000 22614
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 0 21994 800 22024
rect 1485 21994 1551 21997
rect 0 21992 1551 21994
rect 0 21936 1490 21992
rect 1546 21936 1551 21992
rect 0 21934 1551 21936
rect 0 21904 800 21934
rect 1485 21931 1551 21934
rect 78029 21994 78095 21997
rect 79200 21994 80000 22024
rect 78029 21992 80000 21994
rect 78029 21936 78034 21992
rect 78090 21936 80000 21992
rect 78029 21934 80000 21936
rect 78029 21931 78095 21934
rect 79200 21904 80000 21934
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 0 21314 800 21344
rect 1485 21314 1551 21317
rect 0 21312 1551 21314
rect 0 21256 1490 21312
rect 1546 21256 1551 21312
rect 0 21254 1551 21256
rect 0 21224 800 21254
rect 1485 21251 1551 21254
rect 77845 21314 77911 21317
rect 79200 21314 80000 21344
rect 77845 21312 80000 21314
rect 77845 21256 77850 21312
rect 77906 21256 80000 21312
rect 77845 21254 80000 21256
rect 77845 21251 77911 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 79200 21224 80000 21254
rect 65650 21183 65966 21184
rect 19570 20704 19886 20705
rect 0 20634 800 20664
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 1485 20634 1551 20637
rect 0 20632 1551 20634
rect 0 20576 1490 20632
rect 1546 20576 1551 20632
rect 0 20574 1551 20576
rect 0 20544 800 20574
rect 1485 20571 1551 20574
rect 78029 20634 78095 20637
rect 79200 20634 80000 20664
rect 78029 20632 80000 20634
rect 78029 20576 78034 20632
rect 78090 20576 80000 20632
rect 78029 20574 80000 20576
rect 78029 20571 78095 20574
rect 79200 20544 80000 20574
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 0 19954 800 19984
rect 1485 19954 1551 19957
rect 0 19952 1551 19954
rect 0 19896 1490 19952
rect 1546 19896 1551 19952
rect 0 19894 1551 19896
rect 0 19864 800 19894
rect 1485 19891 1551 19894
rect 77845 19954 77911 19957
rect 79200 19954 80000 19984
rect 77845 19952 80000 19954
rect 77845 19896 77850 19952
rect 77906 19896 80000 19952
rect 77845 19894 80000 19896
rect 77845 19891 77911 19894
rect 79200 19864 80000 19894
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 0 19274 800 19304
rect 1485 19274 1551 19277
rect 0 19272 1551 19274
rect 0 19216 1490 19272
rect 1546 19216 1551 19272
rect 0 19214 1551 19216
rect 0 19184 800 19214
rect 1485 19211 1551 19214
rect 77845 19274 77911 19277
rect 79200 19274 80000 19304
rect 77845 19272 80000 19274
rect 77845 19216 77850 19272
rect 77906 19216 80000 19272
rect 77845 19214 80000 19216
rect 77845 19211 77911 19214
rect 79200 19184 80000 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 0 18594 800 18624
rect 1485 18594 1551 18597
rect 0 18592 1551 18594
rect 0 18536 1490 18592
rect 1546 18536 1551 18592
rect 0 18534 1551 18536
rect 0 18504 800 18534
rect 1485 18531 1551 18534
rect 78029 18594 78095 18597
rect 79200 18594 80000 18624
rect 78029 18592 80000 18594
rect 78029 18536 78034 18592
rect 78090 18536 80000 18592
rect 78029 18534 80000 18536
rect 78029 18531 78095 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 79200 18504 80000 18534
rect 50290 18463 50606 18464
rect 4210 17984 4526 17985
rect 0 17914 800 17944
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 1485 17914 1551 17917
rect 0 17912 1551 17914
rect 0 17856 1490 17912
rect 1546 17856 1551 17912
rect 0 17854 1551 17856
rect 0 17824 800 17854
rect 1485 17851 1551 17854
rect 77845 17914 77911 17917
rect 79200 17914 80000 17944
rect 77845 17912 80000 17914
rect 77845 17856 77850 17912
rect 77906 17856 80000 17912
rect 77845 17854 80000 17856
rect 77845 17851 77911 17854
rect 79200 17824 80000 17854
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 78029 17234 78095 17237
rect 79200 17234 80000 17264
rect 78029 17232 80000 17234
rect 78029 17176 78034 17232
rect 78090 17176 80000 17232
rect 78029 17174 80000 17176
rect 78029 17171 78095 17174
rect 79200 17144 80000 17174
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 0 16554 800 16584
rect 1485 16554 1551 16557
rect 0 16552 1551 16554
rect 0 16496 1490 16552
rect 1546 16496 1551 16552
rect 0 16494 1551 16496
rect 0 16464 800 16494
rect 1485 16491 1551 16494
rect 78029 16554 78095 16557
rect 79200 16554 80000 16584
rect 78029 16552 80000 16554
rect 78029 16496 78034 16552
rect 78090 16496 80000 16552
rect 78029 16494 80000 16496
rect 78029 16491 78095 16494
rect 79200 16464 80000 16494
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 0 15874 800 15904
rect 1485 15874 1551 15877
rect 0 15872 1551 15874
rect 0 15816 1490 15872
rect 1546 15816 1551 15872
rect 0 15814 1551 15816
rect 0 15784 800 15814
rect 1485 15811 1551 15814
rect 77845 15874 77911 15877
rect 79200 15874 80000 15904
rect 77845 15872 80000 15874
rect 77845 15816 77850 15872
rect 77906 15816 80000 15872
rect 77845 15814 80000 15816
rect 77845 15811 77911 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 79200 15784 80000 15814
rect 65650 15743 65966 15744
rect 19570 15264 19886 15265
rect 0 15194 800 15224
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 78029 15194 78095 15197
rect 79200 15194 80000 15224
rect 78029 15192 80000 15194
rect 78029 15136 78034 15192
rect 78090 15136 80000 15192
rect 78029 15134 80000 15136
rect 78029 15131 78095 15134
rect 79200 15104 80000 15134
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 0 14514 800 14544
rect 1485 14514 1551 14517
rect 0 14512 1551 14514
rect 0 14456 1490 14512
rect 1546 14456 1551 14512
rect 0 14454 1551 14456
rect 0 14424 800 14454
rect 1485 14451 1551 14454
rect 77845 14514 77911 14517
rect 79200 14514 80000 14544
rect 77845 14512 80000 14514
rect 77845 14456 77850 14512
rect 77906 14456 80000 14512
rect 77845 14454 80000 14456
rect 77845 14451 77911 14454
rect 79200 14424 80000 14454
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 0 13834 800 13864
rect 1485 13834 1551 13837
rect 0 13832 1551 13834
rect 0 13776 1490 13832
rect 1546 13776 1551 13832
rect 0 13774 1551 13776
rect 0 13744 800 13774
rect 1485 13771 1551 13774
rect 77845 13834 77911 13837
rect 79200 13834 80000 13864
rect 77845 13832 80000 13834
rect 77845 13776 77850 13832
rect 77906 13776 80000 13832
rect 77845 13774 80000 13776
rect 77845 13771 77911 13774
rect 79200 13744 80000 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 0 13154 800 13184
rect 1485 13154 1551 13157
rect 0 13152 1551 13154
rect 0 13096 1490 13152
rect 1546 13096 1551 13152
rect 0 13094 1551 13096
rect 0 13064 800 13094
rect 1485 13091 1551 13094
rect 78029 13154 78095 13157
rect 79200 13154 80000 13184
rect 78029 13152 80000 13154
rect 78029 13096 78034 13152
rect 78090 13096 80000 13152
rect 78029 13094 80000 13096
rect 78029 13091 78095 13094
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 79200 13064 80000 13094
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 0 12474 800 12504
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 1485 12474 1551 12477
rect 0 12472 1551 12474
rect 0 12416 1490 12472
rect 1546 12416 1551 12472
rect 0 12414 1551 12416
rect 0 12384 800 12414
rect 1485 12411 1551 12414
rect 77845 12474 77911 12477
rect 79200 12474 80000 12504
rect 77845 12472 80000 12474
rect 77845 12416 77850 12472
rect 77906 12416 80000 12472
rect 77845 12414 80000 12416
rect 77845 12411 77911 12414
rect 79200 12384 80000 12414
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 0 11794 800 11824
rect 1485 11794 1551 11797
rect 0 11792 1551 11794
rect 0 11736 1490 11792
rect 1546 11736 1551 11792
rect 0 11734 1551 11736
rect 0 11704 800 11734
rect 1485 11731 1551 11734
rect 78029 11794 78095 11797
rect 79200 11794 80000 11824
rect 78029 11792 80000 11794
rect 78029 11736 78034 11792
rect 78090 11736 80000 11792
rect 78029 11734 80000 11736
rect 78029 11731 78095 11734
rect 79200 11704 80000 11734
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 0 11114 800 11144
rect 1485 11114 1551 11117
rect 0 11112 1551 11114
rect 0 11056 1490 11112
rect 1546 11056 1551 11112
rect 0 11054 1551 11056
rect 0 11024 800 11054
rect 1485 11051 1551 11054
rect 78029 11114 78095 11117
rect 79200 11114 80000 11144
rect 78029 11112 80000 11114
rect 78029 11056 78034 11112
rect 78090 11056 80000 11112
rect 78029 11054 80000 11056
rect 78029 11051 78095 11054
rect 79200 11024 80000 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 0 10434 800 10464
rect 1485 10434 1551 10437
rect 0 10432 1551 10434
rect 0 10376 1490 10432
rect 1546 10376 1551 10432
rect 0 10374 1551 10376
rect 0 10344 800 10374
rect 1485 10371 1551 10374
rect 77845 10434 77911 10437
rect 79200 10434 80000 10464
rect 77845 10432 80000 10434
rect 77845 10376 77850 10432
rect 77906 10376 80000 10432
rect 77845 10374 80000 10376
rect 77845 10371 77911 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 79200 10344 80000 10374
rect 65650 10303 65966 10304
rect 19570 9824 19886 9825
rect 0 9754 800 9784
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 1485 9754 1551 9757
rect 0 9752 1551 9754
rect 0 9696 1490 9752
rect 1546 9696 1551 9752
rect 0 9694 1551 9696
rect 0 9664 800 9694
rect 1485 9691 1551 9694
rect 78029 9754 78095 9757
rect 79200 9754 80000 9784
rect 78029 9752 80000 9754
rect 78029 9696 78034 9752
rect 78090 9696 80000 9752
rect 78029 9694 80000 9696
rect 78029 9691 78095 9694
rect 79200 9664 80000 9694
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 0 9074 800 9104
rect 1485 9074 1551 9077
rect 0 9072 1551 9074
rect 0 9016 1490 9072
rect 1546 9016 1551 9072
rect 0 9014 1551 9016
rect 0 8984 800 9014
rect 1485 9011 1551 9014
rect 77845 9074 77911 9077
rect 79200 9074 80000 9104
rect 77845 9072 80000 9074
rect 77845 9016 77850 9072
rect 77906 9016 80000 9072
rect 77845 9014 80000 9016
rect 77845 9011 77911 9014
rect 79200 8984 80000 9014
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 0 8394 800 8424
rect 1485 8394 1551 8397
rect 0 8392 1551 8394
rect 0 8336 1490 8392
rect 1546 8336 1551 8392
rect 0 8334 1551 8336
rect 0 8304 800 8334
rect 1485 8331 1551 8334
rect 77845 8394 77911 8397
rect 79200 8394 80000 8424
rect 77845 8392 80000 8394
rect 77845 8336 77850 8392
rect 77906 8336 80000 8392
rect 77845 8334 80000 8336
rect 77845 8331 77911 8334
rect 79200 8304 80000 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 0 7714 800 7744
rect 1485 7714 1551 7717
rect 0 7712 1551 7714
rect 0 7656 1490 7712
rect 1546 7656 1551 7712
rect 0 7654 1551 7656
rect 0 7624 800 7654
rect 1485 7651 1551 7654
rect 78029 7714 78095 7717
rect 79200 7714 80000 7744
rect 78029 7712 80000 7714
rect 78029 7656 78034 7712
rect 78090 7656 80000 7712
rect 78029 7654 80000 7656
rect 78029 7651 78095 7654
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 79200 7624 80000 7654
rect 50290 7583 50606 7584
rect 4210 7104 4526 7105
rect 0 7034 800 7064
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 1485 7034 1551 7037
rect 0 7032 1551 7034
rect 0 6976 1490 7032
rect 1546 6976 1551 7032
rect 0 6974 1551 6976
rect 0 6944 800 6974
rect 1485 6971 1551 6974
rect 77845 7034 77911 7037
rect 79200 7034 80000 7064
rect 77845 7032 80000 7034
rect 77845 6976 77850 7032
rect 77906 6976 80000 7032
rect 77845 6974 80000 6976
rect 77845 6971 77911 6974
rect 79200 6944 80000 6974
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 0 6354 800 6384
rect 1485 6354 1551 6357
rect 0 6352 1551 6354
rect 0 6296 1490 6352
rect 1546 6296 1551 6352
rect 0 6294 1551 6296
rect 0 6264 800 6294
rect 1485 6291 1551 6294
rect 78029 6354 78095 6357
rect 79200 6354 80000 6384
rect 78029 6352 80000 6354
rect 78029 6296 78034 6352
rect 78090 6296 80000 6352
rect 78029 6294 80000 6296
rect 78029 6291 78095 6294
rect 79200 6264 80000 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 0 5674 800 5704
rect 1485 5674 1551 5677
rect 0 5672 1551 5674
rect 0 5616 1490 5672
rect 1546 5616 1551 5672
rect 0 5614 1551 5616
rect 0 5584 800 5614
rect 1485 5611 1551 5614
rect 78029 5674 78095 5677
rect 79200 5674 80000 5704
rect 78029 5672 80000 5674
rect 78029 5616 78034 5672
rect 78090 5616 80000 5672
rect 78029 5614 80000 5616
rect 78029 5611 78095 5614
rect 79200 5584 80000 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 0 4994 800 5024
rect 1485 4994 1551 4997
rect 0 4992 1551 4994
rect 0 4936 1490 4992
rect 1546 4936 1551 4992
rect 0 4934 1551 4936
rect 0 4904 800 4934
rect 1485 4931 1551 4934
rect 77845 4994 77911 4997
rect 79200 4994 80000 5024
rect 77845 4992 80000 4994
rect 77845 4936 77850 4992
rect 77906 4936 80000 4992
rect 77845 4934 80000 4936
rect 77845 4931 77911 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 79200 4904 80000 4934
rect 65650 4863 65966 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 64965 3362 65031 3365
rect 72049 3362 72115 3365
rect 64965 3360 72115 3362
rect 64965 3304 64970 3360
rect 65026 3304 72054 3360
rect 72110 3304 72115 3360
rect 64965 3302 72115 3304
rect 64965 3299 65031 3302
rect 72049 3299 72115 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 65977 3226 66043 3229
rect 69289 3226 69355 3229
rect 65977 3224 69355 3226
rect 65977 3168 65982 3224
rect 66038 3168 69294 3224
rect 69350 3168 69355 3224
rect 65977 3166 69355 3168
rect 65977 3163 66043 3166
rect 69289 3163 69355 3166
rect 53373 2954 53439 2957
rect 77109 2954 77175 2957
rect 53373 2952 77175 2954
rect 53373 2896 53378 2952
rect 53434 2896 77114 2952
rect 77170 2896 77175 2952
rect 53373 2894 77175 2896
rect 53373 2891 53439 2894
rect 77109 2891 77175 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 4216 77820 4280 77824
rect 4216 77764 4220 77820
rect 4220 77764 4276 77820
rect 4276 77764 4280 77820
rect 4216 77760 4280 77764
rect 4296 77820 4360 77824
rect 4296 77764 4300 77820
rect 4300 77764 4356 77820
rect 4356 77764 4360 77820
rect 4296 77760 4360 77764
rect 4376 77820 4440 77824
rect 4376 77764 4380 77820
rect 4380 77764 4436 77820
rect 4436 77764 4440 77820
rect 4376 77760 4440 77764
rect 4456 77820 4520 77824
rect 4456 77764 4460 77820
rect 4460 77764 4516 77820
rect 4516 77764 4520 77820
rect 4456 77760 4520 77764
rect 34936 77820 35000 77824
rect 34936 77764 34940 77820
rect 34940 77764 34996 77820
rect 34996 77764 35000 77820
rect 34936 77760 35000 77764
rect 35016 77820 35080 77824
rect 35016 77764 35020 77820
rect 35020 77764 35076 77820
rect 35076 77764 35080 77820
rect 35016 77760 35080 77764
rect 35096 77820 35160 77824
rect 35096 77764 35100 77820
rect 35100 77764 35156 77820
rect 35156 77764 35160 77820
rect 35096 77760 35160 77764
rect 35176 77820 35240 77824
rect 35176 77764 35180 77820
rect 35180 77764 35236 77820
rect 35236 77764 35240 77820
rect 35176 77760 35240 77764
rect 65656 77820 65720 77824
rect 65656 77764 65660 77820
rect 65660 77764 65716 77820
rect 65716 77764 65720 77820
rect 65656 77760 65720 77764
rect 65736 77820 65800 77824
rect 65736 77764 65740 77820
rect 65740 77764 65796 77820
rect 65796 77764 65800 77820
rect 65736 77760 65800 77764
rect 65816 77820 65880 77824
rect 65816 77764 65820 77820
rect 65820 77764 65876 77820
rect 65876 77764 65880 77820
rect 65816 77760 65880 77764
rect 65896 77820 65960 77824
rect 65896 77764 65900 77820
rect 65900 77764 65956 77820
rect 65956 77764 65960 77820
rect 65896 77760 65960 77764
rect 19576 77276 19640 77280
rect 19576 77220 19580 77276
rect 19580 77220 19636 77276
rect 19636 77220 19640 77276
rect 19576 77216 19640 77220
rect 19656 77276 19720 77280
rect 19656 77220 19660 77276
rect 19660 77220 19716 77276
rect 19716 77220 19720 77276
rect 19656 77216 19720 77220
rect 19736 77276 19800 77280
rect 19736 77220 19740 77276
rect 19740 77220 19796 77276
rect 19796 77220 19800 77276
rect 19736 77216 19800 77220
rect 19816 77276 19880 77280
rect 19816 77220 19820 77276
rect 19820 77220 19876 77276
rect 19876 77220 19880 77276
rect 19816 77216 19880 77220
rect 50296 77276 50360 77280
rect 50296 77220 50300 77276
rect 50300 77220 50356 77276
rect 50356 77220 50360 77276
rect 50296 77216 50360 77220
rect 50376 77276 50440 77280
rect 50376 77220 50380 77276
rect 50380 77220 50436 77276
rect 50436 77220 50440 77276
rect 50376 77216 50440 77220
rect 50456 77276 50520 77280
rect 50456 77220 50460 77276
rect 50460 77220 50516 77276
rect 50516 77220 50520 77276
rect 50456 77216 50520 77220
rect 50536 77276 50600 77280
rect 50536 77220 50540 77276
rect 50540 77220 50596 77276
rect 50596 77220 50600 77276
rect 50536 77216 50600 77220
rect 4216 76732 4280 76736
rect 4216 76676 4220 76732
rect 4220 76676 4276 76732
rect 4276 76676 4280 76732
rect 4216 76672 4280 76676
rect 4296 76732 4360 76736
rect 4296 76676 4300 76732
rect 4300 76676 4356 76732
rect 4356 76676 4360 76732
rect 4296 76672 4360 76676
rect 4376 76732 4440 76736
rect 4376 76676 4380 76732
rect 4380 76676 4436 76732
rect 4436 76676 4440 76732
rect 4376 76672 4440 76676
rect 4456 76732 4520 76736
rect 4456 76676 4460 76732
rect 4460 76676 4516 76732
rect 4516 76676 4520 76732
rect 4456 76672 4520 76676
rect 34936 76732 35000 76736
rect 34936 76676 34940 76732
rect 34940 76676 34996 76732
rect 34996 76676 35000 76732
rect 34936 76672 35000 76676
rect 35016 76732 35080 76736
rect 35016 76676 35020 76732
rect 35020 76676 35076 76732
rect 35076 76676 35080 76732
rect 35016 76672 35080 76676
rect 35096 76732 35160 76736
rect 35096 76676 35100 76732
rect 35100 76676 35156 76732
rect 35156 76676 35160 76732
rect 35096 76672 35160 76676
rect 35176 76732 35240 76736
rect 35176 76676 35180 76732
rect 35180 76676 35236 76732
rect 35236 76676 35240 76732
rect 35176 76672 35240 76676
rect 65656 76732 65720 76736
rect 65656 76676 65660 76732
rect 65660 76676 65716 76732
rect 65716 76676 65720 76732
rect 65656 76672 65720 76676
rect 65736 76732 65800 76736
rect 65736 76676 65740 76732
rect 65740 76676 65796 76732
rect 65796 76676 65800 76732
rect 65736 76672 65800 76676
rect 65816 76732 65880 76736
rect 65816 76676 65820 76732
rect 65820 76676 65876 76732
rect 65876 76676 65880 76732
rect 65816 76672 65880 76676
rect 65896 76732 65960 76736
rect 65896 76676 65900 76732
rect 65900 76676 65956 76732
rect 65956 76676 65960 76732
rect 65896 76672 65960 76676
rect 19576 76188 19640 76192
rect 19576 76132 19580 76188
rect 19580 76132 19636 76188
rect 19636 76132 19640 76188
rect 19576 76128 19640 76132
rect 19656 76188 19720 76192
rect 19656 76132 19660 76188
rect 19660 76132 19716 76188
rect 19716 76132 19720 76188
rect 19656 76128 19720 76132
rect 19736 76188 19800 76192
rect 19736 76132 19740 76188
rect 19740 76132 19796 76188
rect 19796 76132 19800 76188
rect 19736 76128 19800 76132
rect 19816 76188 19880 76192
rect 19816 76132 19820 76188
rect 19820 76132 19876 76188
rect 19876 76132 19880 76188
rect 19816 76128 19880 76132
rect 50296 76188 50360 76192
rect 50296 76132 50300 76188
rect 50300 76132 50356 76188
rect 50356 76132 50360 76188
rect 50296 76128 50360 76132
rect 50376 76188 50440 76192
rect 50376 76132 50380 76188
rect 50380 76132 50436 76188
rect 50436 76132 50440 76188
rect 50376 76128 50440 76132
rect 50456 76188 50520 76192
rect 50456 76132 50460 76188
rect 50460 76132 50516 76188
rect 50516 76132 50520 76188
rect 50456 76128 50520 76132
rect 50536 76188 50600 76192
rect 50536 76132 50540 76188
rect 50540 76132 50596 76188
rect 50596 76132 50600 76188
rect 50536 76128 50600 76132
rect 4216 75644 4280 75648
rect 4216 75588 4220 75644
rect 4220 75588 4276 75644
rect 4276 75588 4280 75644
rect 4216 75584 4280 75588
rect 4296 75644 4360 75648
rect 4296 75588 4300 75644
rect 4300 75588 4356 75644
rect 4356 75588 4360 75644
rect 4296 75584 4360 75588
rect 4376 75644 4440 75648
rect 4376 75588 4380 75644
rect 4380 75588 4436 75644
rect 4436 75588 4440 75644
rect 4376 75584 4440 75588
rect 4456 75644 4520 75648
rect 4456 75588 4460 75644
rect 4460 75588 4516 75644
rect 4516 75588 4520 75644
rect 4456 75584 4520 75588
rect 34936 75644 35000 75648
rect 34936 75588 34940 75644
rect 34940 75588 34996 75644
rect 34996 75588 35000 75644
rect 34936 75584 35000 75588
rect 35016 75644 35080 75648
rect 35016 75588 35020 75644
rect 35020 75588 35076 75644
rect 35076 75588 35080 75644
rect 35016 75584 35080 75588
rect 35096 75644 35160 75648
rect 35096 75588 35100 75644
rect 35100 75588 35156 75644
rect 35156 75588 35160 75644
rect 35096 75584 35160 75588
rect 35176 75644 35240 75648
rect 35176 75588 35180 75644
rect 35180 75588 35236 75644
rect 35236 75588 35240 75644
rect 35176 75584 35240 75588
rect 65656 75644 65720 75648
rect 65656 75588 65660 75644
rect 65660 75588 65716 75644
rect 65716 75588 65720 75644
rect 65656 75584 65720 75588
rect 65736 75644 65800 75648
rect 65736 75588 65740 75644
rect 65740 75588 65796 75644
rect 65796 75588 65800 75644
rect 65736 75584 65800 75588
rect 65816 75644 65880 75648
rect 65816 75588 65820 75644
rect 65820 75588 65876 75644
rect 65876 75588 65880 75644
rect 65816 75584 65880 75588
rect 65896 75644 65960 75648
rect 65896 75588 65900 75644
rect 65900 75588 65956 75644
rect 65956 75588 65960 75644
rect 65896 75584 65960 75588
rect 1716 75304 1780 75308
rect 1716 75248 1730 75304
rect 1730 75248 1780 75304
rect 1716 75244 1780 75248
rect 19576 75100 19640 75104
rect 19576 75044 19580 75100
rect 19580 75044 19636 75100
rect 19636 75044 19640 75100
rect 19576 75040 19640 75044
rect 19656 75100 19720 75104
rect 19656 75044 19660 75100
rect 19660 75044 19716 75100
rect 19716 75044 19720 75100
rect 19656 75040 19720 75044
rect 19736 75100 19800 75104
rect 19736 75044 19740 75100
rect 19740 75044 19796 75100
rect 19796 75044 19800 75100
rect 19736 75040 19800 75044
rect 19816 75100 19880 75104
rect 19816 75044 19820 75100
rect 19820 75044 19876 75100
rect 19876 75044 19880 75100
rect 19816 75040 19880 75044
rect 50296 75100 50360 75104
rect 50296 75044 50300 75100
rect 50300 75044 50356 75100
rect 50356 75044 50360 75100
rect 50296 75040 50360 75044
rect 50376 75100 50440 75104
rect 50376 75044 50380 75100
rect 50380 75044 50436 75100
rect 50436 75044 50440 75100
rect 50376 75040 50440 75044
rect 50456 75100 50520 75104
rect 50456 75044 50460 75100
rect 50460 75044 50516 75100
rect 50516 75044 50520 75100
rect 50456 75040 50520 75044
rect 50536 75100 50600 75104
rect 50536 75044 50540 75100
rect 50540 75044 50596 75100
rect 50596 75044 50600 75100
rect 50536 75040 50600 75044
rect 4216 74556 4280 74560
rect 4216 74500 4220 74556
rect 4220 74500 4276 74556
rect 4276 74500 4280 74556
rect 4216 74496 4280 74500
rect 4296 74556 4360 74560
rect 4296 74500 4300 74556
rect 4300 74500 4356 74556
rect 4356 74500 4360 74556
rect 4296 74496 4360 74500
rect 4376 74556 4440 74560
rect 4376 74500 4380 74556
rect 4380 74500 4436 74556
rect 4436 74500 4440 74556
rect 4376 74496 4440 74500
rect 4456 74556 4520 74560
rect 4456 74500 4460 74556
rect 4460 74500 4516 74556
rect 4516 74500 4520 74556
rect 4456 74496 4520 74500
rect 34936 74556 35000 74560
rect 34936 74500 34940 74556
rect 34940 74500 34996 74556
rect 34996 74500 35000 74556
rect 34936 74496 35000 74500
rect 35016 74556 35080 74560
rect 35016 74500 35020 74556
rect 35020 74500 35076 74556
rect 35076 74500 35080 74556
rect 35016 74496 35080 74500
rect 35096 74556 35160 74560
rect 35096 74500 35100 74556
rect 35100 74500 35156 74556
rect 35156 74500 35160 74556
rect 35096 74496 35160 74500
rect 35176 74556 35240 74560
rect 35176 74500 35180 74556
rect 35180 74500 35236 74556
rect 35236 74500 35240 74556
rect 35176 74496 35240 74500
rect 65656 74556 65720 74560
rect 65656 74500 65660 74556
rect 65660 74500 65716 74556
rect 65716 74500 65720 74556
rect 65656 74496 65720 74500
rect 65736 74556 65800 74560
rect 65736 74500 65740 74556
rect 65740 74500 65796 74556
rect 65796 74500 65800 74556
rect 65736 74496 65800 74500
rect 65816 74556 65880 74560
rect 65816 74500 65820 74556
rect 65820 74500 65876 74556
rect 65876 74500 65880 74556
rect 65816 74496 65880 74500
rect 65896 74556 65960 74560
rect 65896 74500 65900 74556
rect 65900 74500 65956 74556
rect 65956 74500 65960 74556
rect 65896 74496 65960 74500
rect 19576 74012 19640 74016
rect 19576 73956 19580 74012
rect 19580 73956 19636 74012
rect 19636 73956 19640 74012
rect 19576 73952 19640 73956
rect 19656 74012 19720 74016
rect 19656 73956 19660 74012
rect 19660 73956 19716 74012
rect 19716 73956 19720 74012
rect 19656 73952 19720 73956
rect 19736 74012 19800 74016
rect 19736 73956 19740 74012
rect 19740 73956 19796 74012
rect 19796 73956 19800 74012
rect 19736 73952 19800 73956
rect 19816 74012 19880 74016
rect 19816 73956 19820 74012
rect 19820 73956 19876 74012
rect 19876 73956 19880 74012
rect 19816 73952 19880 73956
rect 50296 74012 50360 74016
rect 50296 73956 50300 74012
rect 50300 73956 50356 74012
rect 50356 73956 50360 74012
rect 50296 73952 50360 73956
rect 50376 74012 50440 74016
rect 50376 73956 50380 74012
rect 50380 73956 50436 74012
rect 50436 73956 50440 74012
rect 50376 73952 50440 73956
rect 50456 74012 50520 74016
rect 50456 73956 50460 74012
rect 50460 73956 50516 74012
rect 50516 73956 50520 74012
rect 50456 73952 50520 73956
rect 50536 74012 50600 74016
rect 50536 73956 50540 74012
rect 50540 73956 50596 74012
rect 50596 73956 50600 74012
rect 50536 73952 50600 73956
rect 4216 73468 4280 73472
rect 4216 73412 4220 73468
rect 4220 73412 4276 73468
rect 4276 73412 4280 73468
rect 4216 73408 4280 73412
rect 4296 73468 4360 73472
rect 4296 73412 4300 73468
rect 4300 73412 4356 73468
rect 4356 73412 4360 73468
rect 4296 73408 4360 73412
rect 4376 73468 4440 73472
rect 4376 73412 4380 73468
rect 4380 73412 4436 73468
rect 4436 73412 4440 73468
rect 4376 73408 4440 73412
rect 4456 73468 4520 73472
rect 4456 73412 4460 73468
rect 4460 73412 4516 73468
rect 4516 73412 4520 73468
rect 4456 73408 4520 73412
rect 34936 73468 35000 73472
rect 34936 73412 34940 73468
rect 34940 73412 34996 73468
rect 34996 73412 35000 73468
rect 34936 73408 35000 73412
rect 35016 73468 35080 73472
rect 35016 73412 35020 73468
rect 35020 73412 35076 73468
rect 35076 73412 35080 73468
rect 35016 73408 35080 73412
rect 35096 73468 35160 73472
rect 35096 73412 35100 73468
rect 35100 73412 35156 73468
rect 35156 73412 35160 73468
rect 35096 73408 35160 73412
rect 35176 73468 35240 73472
rect 35176 73412 35180 73468
rect 35180 73412 35236 73468
rect 35236 73412 35240 73468
rect 35176 73408 35240 73412
rect 65656 73468 65720 73472
rect 65656 73412 65660 73468
rect 65660 73412 65716 73468
rect 65716 73412 65720 73468
rect 65656 73408 65720 73412
rect 65736 73468 65800 73472
rect 65736 73412 65740 73468
rect 65740 73412 65796 73468
rect 65796 73412 65800 73468
rect 65736 73408 65800 73412
rect 65816 73468 65880 73472
rect 65816 73412 65820 73468
rect 65820 73412 65876 73468
rect 65876 73412 65880 73468
rect 65816 73408 65880 73412
rect 65896 73468 65960 73472
rect 65896 73412 65900 73468
rect 65900 73412 65956 73468
rect 65956 73412 65960 73468
rect 65896 73408 65960 73412
rect 19576 72924 19640 72928
rect 19576 72868 19580 72924
rect 19580 72868 19636 72924
rect 19636 72868 19640 72924
rect 19576 72864 19640 72868
rect 19656 72924 19720 72928
rect 19656 72868 19660 72924
rect 19660 72868 19716 72924
rect 19716 72868 19720 72924
rect 19656 72864 19720 72868
rect 19736 72924 19800 72928
rect 19736 72868 19740 72924
rect 19740 72868 19796 72924
rect 19796 72868 19800 72924
rect 19736 72864 19800 72868
rect 19816 72924 19880 72928
rect 19816 72868 19820 72924
rect 19820 72868 19876 72924
rect 19876 72868 19880 72924
rect 19816 72864 19880 72868
rect 50296 72924 50360 72928
rect 50296 72868 50300 72924
rect 50300 72868 50356 72924
rect 50356 72868 50360 72924
rect 50296 72864 50360 72868
rect 50376 72924 50440 72928
rect 50376 72868 50380 72924
rect 50380 72868 50436 72924
rect 50436 72868 50440 72924
rect 50376 72864 50440 72868
rect 50456 72924 50520 72928
rect 50456 72868 50460 72924
rect 50460 72868 50516 72924
rect 50516 72868 50520 72924
rect 50456 72864 50520 72868
rect 50536 72924 50600 72928
rect 50536 72868 50540 72924
rect 50540 72868 50596 72924
rect 50596 72868 50600 72924
rect 50536 72864 50600 72868
rect 4216 72380 4280 72384
rect 4216 72324 4220 72380
rect 4220 72324 4276 72380
rect 4276 72324 4280 72380
rect 4216 72320 4280 72324
rect 4296 72380 4360 72384
rect 4296 72324 4300 72380
rect 4300 72324 4356 72380
rect 4356 72324 4360 72380
rect 4296 72320 4360 72324
rect 4376 72380 4440 72384
rect 4376 72324 4380 72380
rect 4380 72324 4436 72380
rect 4436 72324 4440 72380
rect 4376 72320 4440 72324
rect 4456 72380 4520 72384
rect 4456 72324 4460 72380
rect 4460 72324 4516 72380
rect 4516 72324 4520 72380
rect 4456 72320 4520 72324
rect 34936 72380 35000 72384
rect 34936 72324 34940 72380
rect 34940 72324 34996 72380
rect 34996 72324 35000 72380
rect 34936 72320 35000 72324
rect 35016 72380 35080 72384
rect 35016 72324 35020 72380
rect 35020 72324 35076 72380
rect 35076 72324 35080 72380
rect 35016 72320 35080 72324
rect 35096 72380 35160 72384
rect 35096 72324 35100 72380
rect 35100 72324 35156 72380
rect 35156 72324 35160 72380
rect 35096 72320 35160 72324
rect 35176 72380 35240 72384
rect 35176 72324 35180 72380
rect 35180 72324 35236 72380
rect 35236 72324 35240 72380
rect 35176 72320 35240 72324
rect 65656 72380 65720 72384
rect 65656 72324 65660 72380
rect 65660 72324 65716 72380
rect 65716 72324 65720 72380
rect 65656 72320 65720 72324
rect 65736 72380 65800 72384
rect 65736 72324 65740 72380
rect 65740 72324 65796 72380
rect 65796 72324 65800 72380
rect 65736 72320 65800 72324
rect 65816 72380 65880 72384
rect 65816 72324 65820 72380
rect 65820 72324 65876 72380
rect 65876 72324 65880 72380
rect 65816 72320 65880 72324
rect 65896 72380 65960 72384
rect 65896 72324 65900 72380
rect 65900 72324 65956 72380
rect 65956 72324 65960 72380
rect 65896 72320 65960 72324
rect 19576 71836 19640 71840
rect 19576 71780 19580 71836
rect 19580 71780 19636 71836
rect 19636 71780 19640 71836
rect 19576 71776 19640 71780
rect 19656 71836 19720 71840
rect 19656 71780 19660 71836
rect 19660 71780 19716 71836
rect 19716 71780 19720 71836
rect 19656 71776 19720 71780
rect 19736 71836 19800 71840
rect 19736 71780 19740 71836
rect 19740 71780 19796 71836
rect 19796 71780 19800 71836
rect 19736 71776 19800 71780
rect 19816 71836 19880 71840
rect 19816 71780 19820 71836
rect 19820 71780 19876 71836
rect 19876 71780 19880 71836
rect 19816 71776 19880 71780
rect 50296 71836 50360 71840
rect 50296 71780 50300 71836
rect 50300 71780 50356 71836
rect 50356 71780 50360 71836
rect 50296 71776 50360 71780
rect 50376 71836 50440 71840
rect 50376 71780 50380 71836
rect 50380 71780 50436 71836
rect 50436 71780 50440 71836
rect 50376 71776 50440 71780
rect 50456 71836 50520 71840
rect 50456 71780 50460 71836
rect 50460 71780 50516 71836
rect 50516 71780 50520 71836
rect 50456 71776 50520 71780
rect 50536 71836 50600 71840
rect 50536 71780 50540 71836
rect 50540 71780 50596 71836
rect 50596 71780 50600 71836
rect 50536 71776 50600 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 34936 71292 35000 71296
rect 34936 71236 34940 71292
rect 34940 71236 34996 71292
rect 34996 71236 35000 71292
rect 34936 71232 35000 71236
rect 35016 71292 35080 71296
rect 35016 71236 35020 71292
rect 35020 71236 35076 71292
rect 35076 71236 35080 71292
rect 35016 71232 35080 71236
rect 35096 71292 35160 71296
rect 35096 71236 35100 71292
rect 35100 71236 35156 71292
rect 35156 71236 35160 71292
rect 35096 71232 35160 71236
rect 35176 71292 35240 71296
rect 35176 71236 35180 71292
rect 35180 71236 35236 71292
rect 35236 71236 35240 71292
rect 35176 71232 35240 71236
rect 65656 71292 65720 71296
rect 65656 71236 65660 71292
rect 65660 71236 65716 71292
rect 65716 71236 65720 71292
rect 65656 71232 65720 71236
rect 65736 71292 65800 71296
rect 65736 71236 65740 71292
rect 65740 71236 65796 71292
rect 65796 71236 65800 71292
rect 65736 71232 65800 71236
rect 65816 71292 65880 71296
rect 65816 71236 65820 71292
rect 65820 71236 65876 71292
rect 65876 71236 65880 71292
rect 65816 71232 65880 71236
rect 65896 71292 65960 71296
rect 65896 71236 65900 71292
rect 65900 71236 65956 71292
rect 65956 71236 65960 71292
rect 65896 71232 65960 71236
rect 19576 70748 19640 70752
rect 19576 70692 19580 70748
rect 19580 70692 19636 70748
rect 19636 70692 19640 70748
rect 19576 70688 19640 70692
rect 19656 70748 19720 70752
rect 19656 70692 19660 70748
rect 19660 70692 19716 70748
rect 19716 70692 19720 70748
rect 19656 70688 19720 70692
rect 19736 70748 19800 70752
rect 19736 70692 19740 70748
rect 19740 70692 19796 70748
rect 19796 70692 19800 70748
rect 19736 70688 19800 70692
rect 19816 70748 19880 70752
rect 19816 70692 19820 70748
rect 19820 70692 19876 70748
rect 19876 70692 19880 70748
rect 19816 70688 19880 70692
rect 50296 70748 50360 70752
rect 50296 70692 50300 70748
rect 50300 70692 50356 70748
rect 50356 70692 50360 70748
rect 50296 70688 50360 70692
rect 50376 70748 50440 70752
rect 50376 70692 50380 70748
rect 50380 70692 50436 70748
rect 50436 70692 50440 70748
rect 50376 70688 50440 70692
rect 50456 70748 50520 70752
rect 50456 70692 50460 70748
rect 50460 70692 50516 70748
rect 50516 70692 50520 70748
rect 50456 70688 50520 70692
rect 50536 70748 50600 70752
rect 50536 70692 50540 70748
rect 50540 70692 50596 70748
rect 50596 70692 50600 70748
rect 50536 70688 50600 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 34936 70204 35000 70208
rect 34936 70148 34940 70204
rect 34940 70148 34996 70204
rect 34996 70148 35000 70204
rect 34936 70144 35000 70148
rect 35016 70204 35080 70208
rect 35016 70148 35020 70204
rect 35020 70148 35076 70204
rect 35076 70148 35080 70204
rect 35016 70144 35080 70148
rect 35096 70204 35160 70208
rect 35096 70148 35100 70204
rect 35100 70148 35156 70204
rect 35156 70148 35160 70204
rect 35096 70144 35160 70148
rect 35176 70204 35240 70208
rect 35176 70148 35180 70204
rect 35180 70148 35236 70204
rect 35236 70148 35240 70204
rect 35176 70144 35240 70148
rect 65656 70204 65720 70208
rect 65656 70148 65660 70204
rect 65660 70148 65716 70204
rect 65716 70148 65720 70204
rect 65656 70144 65720 70148
rect 65736 70204 65800 70208
rect 65736 70148 65740 70204
rect 65740 70148 65796 70204
rect 65796 70148 65800 70204
rect 65736 70144 65800 70148
rect 65816 70204 65880 70208
rect 65816 70148 65820 70204
rect 65820 70148 65876 70204
rect 65876 70148 65880 70204
rect 65816 70144 65880 70148
rect 65896 70204 65960 70208
rect 65896 70148 65900 70204
rect 65900 70148 65956 70204
rect 65956 70148 65960 70204
rect 65896 70144 65960 70148
rect 19576 69660 19640 69664
rect 19576 69604 19580 69660
rect 19580 69604 19636 69660
rect 19636 69604 19640 69660
rect 19576 69600 19640 69604
rect 19656 69660 19720 69664
rect 19656 69604 19660 69660
rect 19660 69604 19716 69660
rect 19716 69604 19720 69660
rect 19656 69600 19720 69604
rect 19736 69660 19800 69664
rect 19736 69604 19740 69660
rect 19740 69604 19796 69660
rect 19796 69604 19800 69660
rect 19736 69600 19800 69604
rect 19816 69660 19880 69664
rect 19816 69604 19820 69660
rect 19820 69604 19876 69660
rect 19876 69604 19880 69660
rect 19816 69600 19880 69604
rect 50296 69660 50360 69664
rect 50296 69604 50300 69660
rect 50300 69604 50356 69660
rect 50356 69604 50360 69660
rect 50296 69600 50360 69604
rect 50376 69660 50440 69664
rect 50376 69604 50380 69660
rect 50380 69604 50436 69660
rect 50436 69604 50440 69660
rect 50376 69600 50440 69604
rect 50456 69660 50520 69664
rect 50456 69604 50460 69660
rect 50460 69604 50516 69660
rect 50516 69604 50520 69660
rect 50456 69600 50520 69604
rect 50536 69660 50600 69664
rect 50536 69604 50540 69660
rect 50540 69604 50596 69660
rect 50596 69604 50600 69660
rect 50536 69600 50600 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 34936 69116 35000 69120
rect 34936 69060 34940 69116
rect 34940 69060 34996 69116
rect 34996 69060 35000 69116
rect 34936 69056 35000 69060
rect 35016 69116 35080 69120
rect 35016 69060 35020 69116
rect 35020 69060 35076 69116
rect 35076 69060 35080 69116
rect 35016 69056 35080 69060
rect 35096 69116 35160 69120
rect 35096 69060 35100 69116
rect 35100 69060 35156 69116
rect 35156 69060 35160 69116
rect 35096 69056 35160 69060
rect 35176 69116 35240 69120
rect 35176 69060 35180 69116
rect 35180 69060 35236 69116
rect 35236 69060 35240 69116
rect 35176 69056 35240 69060
rect 65656 69116 65720 69120
rect 65656 69060 65660 69116
rect 65660 69060 65716 69116
rect 65716 69060 65720 69116
rect 65656 69056 65720 69060
rect 65736 69116 65800 69120
rect 65736 69060 65740 69116
rect 65740 69060 65796 69116
rect 65796 69060 65800 69116
rect 65736 69056 65800 69060
rect 65816 69116 65880 69120
rect 65816 69060 65820 69116
rect 65820 69060 65876 69116
rect 65876 69060 65880 69116
rect 65816 69056 65880 69060
rect 65896 69116 65960 69120
rect 65896 69060 65900 69116
rect 65900 69060 65956 69116
rect 65956 69060 65960 69116
rect 65896 69056 65960 69060
rect 19576 68572 19640 68576
rect 19576 68516 19580 68572
rect 19580 68516 19636 68572
rect 19636 68516 19640 68572
rect 19576 68512 19640 68516
rect 19656 68572 19720 68576
rect 19656 68516 19660 68572
rect 19660 68516 19716 68572
rect 19716 68516 19720 68572
rect 19656 68512 19720 68516
rect 19736 68572 19800 68576
rect 19736 68516 19740 68572
rect 19740 68516 19796 68572
rect 19796 68516 19800 68572
rect 19736 68512 19800 68516
rect 19816 68572 19880 68576
rect 19816 68516 19820 68572
rect 19820 68516 19876 68572
rect 19876 68516 19880 68572
rect 19816 68512 19880 68516
rect 50296 68572 50360 68576
rect 50296 68516 50300 68572
rect 50300 68516 50356 68572
rect 50356 68516 50360 68572
rect 50296 68512 50360 68516
rect 50376 68572 50440 68576
rect 50376 68516 50380 68572
rect 50380 68516 50436 68572
rect 50436 68516 50440 68572
rect 50376 68512 50440 68516
rect 50456 68572 50520 68576
rect 50456 68516 50460 68572
rect 50460 68516 50516 68572
rect 50516 68516 50520 68572
rect 50456 68512 50520 68516
rect 50536 68572 50600 68576
rect 50536 68516 50540 68572
rect 50540 68516 50596 68572
rect 50596 68516 50600 68572
rect 50536 68512 50600 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 34936 68028 35000 68032
rect 34936 67972 34940 68028
rect 34940 67972 34996 68028
rect 34996 67972 35000 68028
rect 34936 67968 35000 67972
rect 35016 68028 35080 68032
rect 35016 67972 35020 68028
rect 35020 67972 35076 68028
rect 35076 67972 35080 68028
rect 35016 67968 35080 67972
rect 35096 68028 35160 68032
rect 35096 67972 35100 68028
rect 35100 67972 35156 68028
rect 35156 67972 35160 68028
rect 35096 67968 35160 67972
rect 35176 68028 35240 68032
rect 35176 67972 35180 68028
rect 35180 67972 35236 68028
rect 35236 67972 35240 68028
rect 35176 67968 35240 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 19576 67484 19640 67488
rect 19576 67428 19580 67484
rect 19580 67428 19636 67484
rect 19636 67428 19640 67484
rect 19576 67424 19640 67428
rect 19656 67484 19720 67488
rect 19656 67428 19660 67484
rect 19660 67428 19716 67484
rect 19716 67428 19720 67484
rect 19656 67424 19720 67428
rect 19736 67484 19800 67488
rect 19736 67428 19740 67484
rect 19740 67428 19796 67484
rect 19796 67428 19800 67484
rect 19736 67424 19800 67428
rect 19816 67484 19880 67488
rect 19816 67428 19820 67484
rect 19820 67428 19876 67484
rect 19876 67428 19880 67484
rect 19816 67424 19880 67428
rect 50296 67484 50360 67488
rect 50296 67428 50300 67484
rect 50300 67428 50356 67484
rect 50356 67428 50360 67484
rect 50296 67424 50360 67428
rect 50376 67484 50440 67488
rect 50376 67428 50380 67484
rect 50380 67428 50436 67484
rect 50436 67428 50440 67484
rect 50376 67424 50440 67428
rect 50456 67484 50520 67488
rect 50456 67428 50460 67484
rect 50460 67428 50516 67484
rect 50516 67428 50520 67484
rect 50456 67424 50520 67428
rect 50536 67484 50600 67488
rect 50536 67428 50540 67484
rect 50540 67428 50596 67484
rect 50596 67428 50600 67484
rect 50536 67424 50600 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 19576 66396 19640 66400
rect 19576 66340 19580 66396
rect 19580 66340 19636 66396
rect 19636 66340 19640 66396
rect 19576 66336 19640 66340
rect 19656 66396 19720 66400
rect 19656 66340 19660 66396
rect 19660 66340 19716 66396
rect 19716 66340 19720 66396
rect 19656 66336 19720 66340
rect 19736 66396 19800 66400
rect 19736 66340 19740 66396
rect 19740 66340 19796 66396
rect 19796 66340 19800 66396
rect 19736 66336 19800 66340
rect 19816 66396 19880 66400
rect 19816 66340 19820 66396
rect 19820 66340 19876 66396
rect 19876 66340 19880 66396
rect 19816 66336 19880 66340
rect 50296 66396 50360 66400
rect 50296 66340 50300 66396
rect 50300 66340 50356 66396
rect 50356 66340 50360 66396
rect 50296 66336 50360 66340
rect 50376 66396 50440 66400
rect 50376 66340 50380 66396
rect 50380 66340 50436 66396
rect 50436 66340 50440 66396
rect 50376 66336 50440 66340
rect 50456 66396 50520 66400
rect 50456 66340 50460 66396
rect 50460 66340 50516 66396
rect 50516 66340 50520 66396
rect 50456 66336 50520 66340
rect 50536 66396 50600 66400
rect 50536 66340 50540 66396
rect 50540 66340 50596 66396
rect 50596 66340 50600 66396
rect 50536 66336 50600 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 19576 65308 19640 65312
rect 19576 65252 19580 65308
rect 19580 65252 19636 65308
rect 19636 65252 19640 65308
rect 19576 65248 19640 65252
rect 19656 65308 19720 65312
rect 19656 65252 19660 65308
rect 19660 65252 19716 65308
rect 19716 65252 19720 65308
rect 19656 65248 19720 65252
rect 19736 65308 19800 65312
rect 19736 65252 19740 65308
rect 19740 65252 19796 65308
rect 19796 65252 19800 65308
rect 19736 65248 19800 65252
rect 19816 65308 19880 65312
rect 19816 65252 19820 65308
rect 19820 65252 19876 65308
rect 19876 65252 19880 65308
rect 19816 65248 19880 65252
rect 50296 65308 50360 65312
rect 50296 65252 50300 65308
rect 50300 65252 50356 65308
rect 50356 65252 50360 65308
rect 50296 65248 50360 65252
rect 50376 65308 50440 65312
rect 50376 65252 50380 65308
rect 50380 65252 50436 65308
rect 50436 65252 50440 65308
rect 50376 65248 50440 65252
rect 50456 65308 50520 65312
rect 50456 65252 50460 65308
rect 50460 65252 50516 65308
rect 50516 65252 50520 65308
rect 50456 65248 50520 65252
rect 50536 65308 50600 65312
rect 50536 65252 50540 65308
rect 50540 65252 50596 65308
rect 50596 65252 50600 65308
rect 50536 65248 50600 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 34936 64764 35000 64768
rect 34936 64708 34940 64764
rect 34940 64708 34996 64764
rect 34996 64708 35000 64764
rect 34936 64704 35000 64708
rect 35016 64764 35080 64768
rect 35016 64708 35020 64764
rect 35020 64708 35076 64764
rect 35076 64708 35080 64764
rect 35016 64704 35080 64708
rect 35096 64764 35160 64768
rect 35096 64708 35100 64764
rect 35100 64708 35156 64764
rect 35156 64708 35160 64764
rect 35096 64704 35160 64708
rect 35176 64764 35240 64768
rect 35176 64708 35180 64764
rect 35180 64708 35236 64764
rect 35236 64708 35240 64764
rect 35176 64704 35240 64708
rect 65656 64764 65720 64768
rect 65656 64708 65660 64764
rect 65660 64708 65716 64764
rect 65716 64708 65720 64764
rect 65656 64704 65720 64708
rect 65736 64764 65800 64768
rect 65736 64708 65740 64764
rect 65740 64708 65796 64764
rect 65796 64708 65800 64764
rect 65736 64704 65800 64708
rect 65816 64764 65880 64768
rect 65816 64708 65820 64764
rect 65820 64708 65876 64764
rect 65876 64708 65880 64764
rect 65816 64704 65880 64708
rect 65896 64764 65960 64768
rect 65896 64708 65900 64764
rect 65900 64708 65956 64764
rect 65956 64708 65960 64764
rect 65896 64704 65960 64708
rect 19576 64220 19640 64224
rect 19576 64164 19580 64220
rect 19580 64164 19636 64220
rect 19636 64164 19640 64220
rect 19576 64160 19640 64164
rect 19656 64220 19720 64224
rect 19656 64164 19660 64220
rect 19660 64164 19716 64220
rect 19716 64164 19720 64220
rect 19656 64160 19720 64164
rect 19736 64220 19800 64224
rect 19736 64164 19740 64220
rect 19740 64164 19796 64220
rect 19796 64164 19800 64220
rect 19736 64160 19800 64164
rect 19816 64220 19880 64224
rect 19816 64164 19820 64220
rect 19820 64164 19876 64220
rect 19876 64164 19880 64220
rect 19816 64160 19880 64164
rect 50296 64220 50360 64224
rect 50296 64164 50300 64220
rect 50300 64164 50356 64220
rect 50356 64164 50360 64220
rect 50296 64160 50360 64164
rect 50376 64220 50440 64224
rect 50376 64164 50380 64220
rect 50380 64164 50436 64220
rect 50436 64164 50440 64220
rect 50376 64160 50440 64164
rect 50456 64220 50520 64224
rect 50456 64164 50460 64220
rect 50460 64164 50516 64220
rect 50516 64164 50520 64220
rect 50456 64160 50520 64164
rect 50536 64220 50600 64224
rect 50536 64164 50540 64220
rect 50540 64164 50596 64220
rect 50596 64164 50600 64220
rect 50536 64160 50600 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 34936 63676 35000 63680
rect 34936 63620 34940 63676
rect 34940 63620 34996 63676
rect 34996 63620 35000 63676
rect 34936 63616 35000 63620
rect 35016 63676 35080 63680
rect 35016 63620 35020 63676
rect 35020 63620 35076 63676
rect 35076 63620 35080 63676
rect 35016 63616 35080 63620
rect 35096 63676 35160 63680
rect 35096 63620 35100 63676
rect 35100 63620 35156 63676
rect 35156 63620 35160 63676
rect 35096 63616 35160 63620
rect 35176 63676 35240 63680
rect 35176 63620 35180 63676
rect 35180 63620 35236 63676
rect 35236 63620 35240 63676
rect 35176 63616 35240 63620
rect 65656 63676 65720 63680
rect 65656 63620 65660 63676
rect 65660 63620 65716 63676
rect 65716 63620 65720 63676
rect 65656 63616 65720 63620
rect 65736 63676 65800 63680
rect 65736 63620 65740 63676
rect 65740 63620 65796 63676
rect 65796 63620 65800 63676
rect 65736 63616 65800 63620
rect 65816 63676 65880 63680
rect 65816 63620 65820 63676
rect 65820 63620 65876 63676
rect 65876 63620 65880 63676
rect 65816 63616 65880 63620
rect 65896 63676 65960 63680
rect 65896 63620 65900 63676
rect 65900 63620 65956 63676
rect 65956 63620 65960 63676
rect 65896 63616 65960 63620
rect 19576 63132 19640 63136
rect 19576 63076 19580 63132
rect 19580 63076 19636 63132
rect 19636 63076 19640 63132
rect 19576 63072 19640 63076
rect 19656 63132 19720 63136
rect 19656 63076 19660 63132
rect 19660 63076 19716 63132
rect 19716 63076 19720 63132
rect 19656 63072 19720 63076
rect 19736 63132 19800 63136
rect 19736 63076 19740 63132
rect 19740 63076 19796 63132
rect 19796 63076 19800 63132
rect 19736 63072 19800 63076
rect 19816 63132 19880 63136
rect 19816 63076 19820 63132
rect 19820 63076 19876 63132
rect 19876 63076 19880 63132
rect 19816 63072 19880 63076
rect 50296 63132 50360 63136
rect 50296 63076 50300 63132
rect 50300 63076 50356 63132
rect 50356 63076 50360 63132
rect 50296 63072 50360 63076
rect 50376 63132 50440 63136
rect 50376 63076 50380 63132
rect 50380 63076 50436 63132
rect 50436 63076 50440 63132
rect 50376 63072 50440 63076
rect 50456 63132 50520 63136
rect 50456 63076 50460 63132
rect 50460 63076 50516 63132
rect 50516 63076 50520 63132
rect 50456 63072 50520 63076
rect 50536 63132 50600 63136
rect 50536 63076 50540 63132
rect 50540 63076 50596 63132
rect 50596 63076 50600 63132
rect 50536 63072 50600 63076
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 34936 62588 35000 62592
rect 34936 62532 34940 62588
rect 34940 62532 34996 62588
rect 34996 62532 35000 62588
rect 34936 62528 35000 62532
rect 35016 62588 35080 62592
rect 35016 62532 35020 62588
rect 35020 62532 35076 62588
rect 35076 62532 35080 62588
rect 35016 62528 35080 62532
rect 35096 62588 35160 62592
rect 35096 62532 35100 62588
rect 35100 62532 35156 62588
rect 35156 62532 35160 62588
rect 35096 62528 35160 62532
rect 35176 62588 35240 62592
rect 35176 62532 35180 62588
rect 35180 62532 35236 62588
rect 35236 62532 35240 62588
rect 35176 62528 35240 62532
rect 65656 62588 65720 62592
rect 65656 62532 65660 62588
rect 65660 62532 65716 62588
rect 65716 62532 65720 62588
rect 65656 62528 65720 62532
rect 65736 62588 65800 62592
rect 65736 62532 65740 62588
rect 65740 62532 65796 62588
rect 65796 62532 65800 62588
rect 65736 62528 65800 62532
rect 65816 62588 65880 62592
rect 65816 62532 65820 62588
rect 65820 62532 65876 62588
rect 65876 62532 65880 62588
rect 65816 62528 65880 62532
rect 65896 62588 65960 62592
rect 65896 62532 65900 62588
rect 65900 62532 65956 62588
rect 65956 62532 65960 62588
rect 65896 62528 65960 62532
rect 19576 62044 19640 62048
rect 19576 61988 19580 62044
rect 19580 61988 19636 62044
rect 19636 61988 19640 62044
rect 19576 61984 19640 61988
rect 19656 62044 19720 62048
rect 19656 61988 19660 62044
rect 19660 61988 19716 62044
rect 19716 61988 19720 62044
rect 19656 61984 19720 61988
rect 19736 62044 19800 62048
rect 19736 61988 19740 62044
rect 19740 61988 19796 62044
rect 19796 61988 19800 62044
rect 19736 61984 19800 61988
rect 19816 62044 19880 62048
rect 19816 61988 19820 62044
rect 19820 61988 19876 62044
rect 19876 61988 19880 62044
rect 19816 61984 19880 61988
rect 50296 62044 50360 62048
rect 50296 61988 50300 62044
rect 50300 61988 50356 62044
rect 50356 61988 50360 62044
rect 50296 61984 50360 61988
rect 50376 62044 50440 62048
rect 50376 61988 50380 62044
rect 50380 61988 50436 62044
rect 50436 61988 50440 62044
rect 50376 61984 50440 61988
rect 50456 62044 50520 62048
rect 50456 61988 50460 62044
rect 50460 61988 50516 62044
rect 50516 61988 50520 62044
rect 50456 61984 50520 61988
rect 50536 62044 50600 62048
rect 50536 61988 50540 62044
rect 50540 61988 50596 62044
rect 50596 61988 50600 62044
rect 50536 61984 50600 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 65656 61500 65720 61504
rect 65656 61444 65660 61500
rect 65660 61444 65716 61500
rect 65716 61444 65720 61500
rect 65656 61440 65720 61444
rect 65736 61500 65800 61504
rect 65736 61444 65740 61500
rect 65740 61444 65796 61500
rect 65796 61444 65800 61500
rect 65736 61440 65800 61444
rect 65816 61500 65880 61504
rect 65816 61444 65820 61500
rect 65820 61444 65876 61500
rect 65876 61444 65880 61500
rect 65816 61440 65880 61444
rect 65896 61500 65960 61504
rect 65896 61444 65900 61500
rect 65900 61444 65956 61500
rect 65956 61444 65960 61500
rect 65896 61440 65960 61444
rect 1716 61100 1780 61164
rect 19576 60956 19640 60960
rect 19576 60900 19580 60956
rect 19580 60900 19636 60956
rect 19636 60900 19640 60956
rect 19576 60896 19640 60900
rect 19656 60956 19720 60960
rect 19656 60900 19660 60956
rect 19660 60900 19716 60956
rect 19716 60900 19720 60956
rect 19656 60896 19720 60900
rect 19736 60956 19800 60960
rect 19736 60900 19740 60956
rect 19740 60900 19796 60956
rect 19796 60900 19800 60956
rect 19736 60896 19800 60900
rect 19816 60956 19880 60960
rect 19816 60900 19820 60956
rect 19820 60900 19876 60956
rect 19876 60900 19880 60956
rect 19816 60896 19880 60900
rect 50296 60956 50360 60960
rect 50296 60900 50300 60956
rect 50300 60900 50356 60956
rect 50356 60900 50360 60956
rect 50296 60896 50360 60900
rect 50376 60956 50440 60960
rect 50376 60900 50380 60956
rect 50380 60900 50436 60956
rect 50436 60900 50440 60956
rect 50376 60896 50440 60900
rect 50456 60956 50520 60960
rect 50456 60900 50460 60956
rect 50460 60900 50516 60956
rect 50516 60900 50520 60956
rect 50456 60896 50520 60900
rect 50536 60956 50600 60960
rect 50536 60900 50540 60956
rect 50540 60900 50596 60956
rect 50596 60900 50600 60956
rect 50536 60896 50600 60900
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 65656 60412 65720 60416
rect 65656 60356 65660 60412
rect 65660 60356 65716 60412
rect 65716 60356 65720 60412
rect 65656 60352 65720 60356
rect 65736 60412 65800 60416
rect 65736 60356 65740 60412
rect 65740 60356 65796 60412
rect 65796 60356 65800 60412
rect 65736 60352 65800 60356
rect 65816 60412 65880 60416
rect 65816 60356 65820 60412
rect 65820 60356 65876 60412
rect 65876 60356 65880 60412
rect 65816 60352 65880 60356
rect 65896 60412 65960 60416
rect 65896 60356 65900 60412
rect 65900 60356 65956 60412
rect 65956 60356 65960 60412
rect 65896 60352 65960 60356
rect 19576 59868 19640 59872
rect 19576 59812 19580 59868
rect 19580 59812 19636 59868
rect 19636 59812 19640 59868
rect 19576 59808 19640 59812
rect 19656 59868 19720 59872
rect 19656 59812 19660 59868
rect 19660 59812 19716 59868
rect 19716 59812 19720 59868
rect 19656 59808 19720 59812
rect 19736 59868 19800 59872
rect 19736 59812 19740 59868
rect 19740 59812 19796 59868
rect 19796 59812 19800 59868
rect 19736 59808 19800 59812
rect 19816 59868 19880 59872
rect 19816 59812 19820 59868
rect 19820 59812 19876 59868
rect 19876 59812 19880 59868
rect 19816 59808 19880 59812
rect 50296 59868 50360 59872
rect 50296 59812 50300 59868
rect 50300 59812 50356 59868
rect 50356 59812 50360 59868
rect 50296 59808 50360 59812
rect 50376 59868 50440 59872
rect 50376 59812 50380 59868
rect 50380 59812 50436 59868
rect 50436 59812 50440 59868
rect 50376 59808 50440 59812
rect 50456 59868 50520 59872
rect 50456 59812 50460 59868
rect 50460 59812 50516 59868
rect 50516 59812 50520 59868
rect 50456 59808 50520 59812
rect 50536 59868 50600 59872
rect 50536 59812 50540 59868
rect 50540 59812 50596 59868
rect 50596 59812 50600 59868
rect 50536 59808 50600 59812
rect 4216 59324 4280 59328
rect 4216 59268 4220 59324
rect 4220 59268 4276 59324
rect 4276 59268 4280 59324
rect 4216 59264 4280 59268
rect 4296 59324 4360 59328
rect 4296 59268 4300 59324
rect 4300 59268 4356 59324
rect 4356 59268 4360 59324
rect 4296 59264 4360 59268
rect 4376 59324 4440 59328
rect 4376 59268 4380 59324
rect 4380 59268 4436 59324
rect 4436 59268 4440 59324
rect 4376 59264 4440 59268
rect 4456 59324 4520 59328
rect 4456 59268 4460 59324
rect 4460 59268 4516 59324
rect 4516 59268 4520 59324
rect 4456 59264 4520 59268
rect 34936 59324 35000 59328
rect 34936 59268 34940 59324
rect 34940 59268 34996 59324
rect 34996 59268 35000 59324
rect 34936 59264 35000 59268
rect 35016 59324 35080 59328
rect 35016 59268 35020 59324
rect 35020 59268 35076 59324
rect 35076 59268 35080 59324
rect 35016 59264 35080 59268
rect 35096 59324 35160 59328
rect 35096 59268 35100 59324
rect 35100 59268 35156 59324
rect 35156 59268 35160 59324
rect 35096 59264 35160 59268
rect 35176 59324 35240 59328
rect 35176 59268 35180 59324
rect 35180 59268 35236 59324
rect 35236 59268 35240 59324
rect 35176 59264 35240 59268
rect 65656 59324 65720 59328
rect 65656 59268 65660 59324
rect 65660 59268 65716 59324
rect 65716 59268 65720 59324
rect 65656 59264 65720 59268
rect 65736 59324 65800 59328
rect 65736 59268 65740 59324
rect 65740 59268 65796 59324
rect 65796 59268 65800 59324
rect 65736 59264 65800 59268
rect 65816 59324 65880 59328
rect 65816 59268 65820 59324
rect 65820 59268 65876 59324
rect 65876 59268 65880 59324
rect 65816 59264 65880 59268
rect 65896 59324 65960 59328
rect 65896 59268 65900 59324
rect 65900 59268 65956 59324
rect 65956 59268 65960 59324
rect 65896 59264 65960 59268
rect 19576 58780 19640 58784
rect 19576 58724 19580 58780
rect 19580 58724 19636 58780
rect 19636 58724 19640 58780
rect 19576 58720 19640 58724
rect 19656 58780 19720 58784
rect 19656 58724 19660 58780
rect 19660 58724 19716 58780
rect 19716 58724 19720 58780
rect 19656 58720 19720 58724
rect 19736 58780 19800 58784
rect 19736 58724 19740 58780
rect 19740 58724 19796 58780
rect 19796 58724 19800 58780
rect 19736 58720 19800 58724
rect 19816 58780 19880 58784
rect 19816 58724 19820 58780
rect 19820 58724 19876 58780
rect 19876 58724 19880 58780
rect 19816 58720 19880 58724
rect 50296 58780 50360 58784
rect 50296 58724 50300 58780
rect 50300 58724 50356 58780
rect 50356 58724 50360 58780
rect 50296 58720 50360 58724
rect 50376 58780 50440 58784
rect 50376 58724 50380 58780
rect 50380 58724 50436 58780
rect 50436 58724 50440 58780
rect 50376 58720 50440 58724
rect 50456 58780 50520 58784
rect 50456 58724 50460 58780
rect 50460 58724 50516 58780
rect 50516 58724 50520 58780
rect 50456 58720 50520 58724
rect 50536 58780 50600 58784
rect 50536 58724 50540 58780
rect 50540 58724 50596 58780
rect 50596 58724 50600 58780
rect 50536 58720 50600 58724
rect 4216 58236 4280 58240
rect 4216 58180 4220 58236
rect 4220 58180 4276 58236
rect 4276 58180 4280 58236
rect 4216 58176 4280 58180
rect 4296 58236 4360 58240
rect 4296 58180 4300 58236
rect 4300 58180 4356 58236
rect 4356 58180 4360 58236
rect 4296 58176 4360 58180
rect 4376 58236 4440 58240
rect 4376 58180 4380 58236
rect 4380 58180 4436 58236
rect 4436 58180 4440 58236
rect 4376 58176 4440 58180
rect 4456 58236 4520 58240
rect 4456 58180 4460 58236
rect 4460 58180 4516 58236
rect 4516 58180 4520 58236
rect 4456 58176 4520 58180
rect 34936 58236 35000 58240
rect 34936 58180 34940 58236
rect 34940 58180 34996 58236
rect 34996 58180 35000 58236
rect 34936 58176 35000 58180
rect 35016 58236 35080 58240
rect 35016 58180 35020 58236
rect 35020 58180 35076 58236
rect 35076 58180 35080 58236
rect 35016 58176 35080 58180
rect 35096 58236 35160 58240
rect 35096 58180 35100 58236
rect 35100 58180 35156 58236
rect 35156 58180 35160 58236
rect 35096 58176 35160 58180
rect 35176 58236 35240 58240
rect 35176 58180 35180 58236
rect 35180 58180 35236 58236
rect 35236 58180 35240 58236
rect 35176 58176 35240 58180
rect 65656 58236 65720 58240
rect 65656 58180 65660 58236
rect 65660 58180 65716 58236
rect 65716 58180 65720 58236
rect 65656 58176 65720 58180
rect 65736 58236 65800 58240
rect 65736 58180 65740 58236
rect 65740 58180 65796 58236
rect 65796 58180 65800 58236
rect 65736 58176 65800 58180
rect 65816 58236 65880 58240
rect 65816 58180 65820 58236
rect 65820 58180 65876 58236
rect 65876 58180 65880 58236
rect 65816 58176 65880 58180
rect 65896 58236 65960 58240
rect 65896 58180 65900 58236
rect 65900 58180 65956 58236
rect 65956 58180 65960 58236
rect 65896 58176 65960 58180
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 77824 4528 77840
rect 4208 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4528 77824
rect 4208 76736 4528 77760
rect 4208 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4528 76736
rect 4208 75648 4528 76672
rect 4208 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4528 75648
rect 1715 75308 1781 75309
rect 1715 75244 1716 75308
rect 1780 75244 1781 75308
rect 1715 75243 1781 75244
rect 1718 61165 1778 75243
rect 4208 74560 4528 75584
rect 4208 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4528 74560
rect 4208 73472 4528 74496
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 72384 4528 73408
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 71296 4528 72320
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4528 66944
rect 4208 65856 4528 66880
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 1715 61164 1781 61165
rect 1715 61100 1716 61164
rect 1780 61100 1781 61164
rect 1715 61099 1781 61100
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59328 4528 60352
rect 4208 59264 4216 59328
rect 4280 59264 4296 59328
rect 4360 59264 4376 59328
rect 4440 59264 4456 59328
rect 4520 59264 4528 59328
rect 4208 58240 4528 59264
rect 4208 58176 4216 58240
rect 4280 58176 4296 58240
rect 4360 58176 4376 58240
rect 4440 58176 4456 58240
rect 4520 58176 4528 58240
rect 4208 57152 4528 58176
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 77280 19888 77840
rect 19568 77216 19576 77280
rect 19640 77216 19656 77280
rect 19720 77216 19736 77280
rect 19800 77216 19816 77280
rect 19880 77216 19888 77280
rect 19568 76192 19888 77216
rect 19568 76128 19576 76192
rect 19640 76128 19656 76192
rect 19720 76128 19736 76192
rect 19800 76128 19816 76192
rect 19880 76128 19888 76192
rect 19568 75104 19888 76128
rect 19568 75040 19576 75104
rect 19640 75040 19656 75104
rect 19720 75040 19736 75104
rect 19800 75040 19816 75104
rect 19880 75040 19888 75104
rect 19568 74016 19888 75040
rect 19568 73952 19576 74016
rect 19640 73952 19656 74016
rect 19720 73952 19736 74016
rect 19800 73952 19816 74016
rect 19880 73952 19888 74016
rect 19568 72928 19888 73952
rect 19568 72864 19576 72928
rect 19640 72864 19656 72928
rect 19720 72864 19736 72928
rect 19800 72864 19816 72928
rect 19880 72864 19888 72928
rect 19568 71840 19888 72864
rect 19568 71776 19576 71840
rect 19640 71776 19656 71840
rect 19720 71776 19736 71840
rect 19800 71776 19816 71840
rect 19880 71776 19888 71840
rect 19568 70752 19888 71776
rect 19568 70688 19576 70752
rect 19640 70688 19656 70752
rect 19720 70688 19736 70752
rect 19800 70688 19816 70752
rect 19880 70688 19888 70752
rect 19568 69664 19888 70688
rect 19568 69600 19576 69664
rect 19640 69600 19656 69664
rect 19720 69600 19736 69664
rect 19800 69600 19816 69664
rect 19880 69600 19888 69664
rect 19568 68576 19888 69600
rect 19568 68512 19576 68576
rect 19640 68512 19656 68576
rect 19720 68512 19736 68576
rect 19800 68512 19816 68576
rect 19880 68512 19888 68576
rect 19568 67488 19888 68512
rect 19568 67424 19576 67488
rect 19640 67424 19656 67488
rect 19720 67424 19736 67488
rect 19800 67424 19816 67488
rect 19880 67424 19888 67488
rect 19568 66400 19888 67424
rect 19568 66336 19576 66400
rect 19640 66336 19656 66400
rect 19720 66336 19736 66400
rect 19800 66336 19816 66400
rect 19880 66336 19888 66400
rect 19568 65312 19888 66336
rect 19568 65248 19576 65312
rect 19640 65248 19656 65312
rect 19720 65248 19736 65312
rect 19800 65248 19816 65312
rect 19880 65248 19888 65312
rect 19568 64224 19888 65248
rect 19568 64160 19576 64224
rect 19640 64160 19656 64224
rect 19720 64160 19736 64224
rect 19800 64160 19816 64224
rect 19880 64160 19888 64224
rect 19568 63136 19888 64160
rect 19568 63072 19576 63136
rect 19640 63072 19656 63136
rect 19720 63072 19736 63136
rect 19800 63072 19816 63136
rect 19880 63072 19888 63136
rect 19568 62048 19888 63072
rect 19568 61984 19576 62048
rect 19640 61984 19656 62048
rect 19720 61984 19736 62048
rect 19800 61984 19816 62048
rect 19880 61984 19888 62048
rect 19568 60960 19888 61984
rect 19568 60896 19576 60960
rect 19640 60896 19656 60960
rect 19720 60896 19736 60960
rect 19800 60896 19816 60960
rect 19880 60896 19888 60960
rect 19568 59872 19888 60896
rect 19568 59808 19576 59872
rect 19640 59808 19656 59872
rect 19720 59808 19736 59872
rect 19800 59808 19816 59872
rect 19880 59808 19888 59872
rect 19568 58784 19888 59808
rect 19568 58720 19576 58784
rect 19640 58720 19656 58784
rect 19720 58720 19736 58784
rect 19800 58720 19816 58784
rect 19880 58720 19888 58784
rect 19568 57696 19888 58720
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 77824 35248 77840
rect 34928 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35248 77824
rect 34928 76736 35248 77760
rect 34928 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35248 76736
rect 34928 75648 35248 76672
rect 34928 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35248 75648
rect 34928 74560 35248 75584
rect 34928 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35248 74560
rect 34928 73472 35248 74496
rect 34928 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35248 73472
rect 34928 72384 35248 73408
rect 34928 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35248 72384
rect 34928 71296 35248 72320
rect 34928 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35248 71296
rect 34928 70208 35248 71232
rect 34928 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35248 70208
rect 34928 69120 35248 70144
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 68032 35248 69056
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 66944 35248 67968
rect 34928 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35248 66944
rect 34928 65856 35248 66880
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 64768 35248 65792
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 63680 35248 64704
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 62592 35248 63616
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 61504 35248 62528
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59328 35248 60352
rect 34928 59264 34936 59328
rect 35000 59264 35016 59328
rect 35080 59264 35096 59328
rect 35160 59264 35176 59328
rect 35240 59264 35248 59328
rect 34928 58240 35248 59264
rect 34928 58176 34936 58240
rect 35000 58176 35016 58240
rect 35080 58176 35096 58240
rect 35160 58176 35176 58240
rect 35240 58176 35248 58240
rect 34928 57152 35248 58176
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 77280 50608 77840
rect 50288 77216 50296 77280
rect 50360 77216 50376 77280
rect 50440 77216 50456 77280
rect 50520 77216 50536 77280
rect 50600 77216 50608 77280
rect 50288 76192 50608 77216
rect 50288 76128 50296 76192
rect 50360 76128 50376 76192
rect 50440 76128 50456 76192
rect 50520 76128 50536 76192
rect 50600 76128 50608 76192
rect 50288 75104 50608 76128
rect 50288 75040 50296 75104
rect 50360 75040 50376 75104
rect 50440 75040 50456 75104
rect 50520 75040 50536 75104
rect 50600 75040 50608 75104
rect 50288 74016 50608 75040
rect 50288 73952 50296 74016
rect 50360 73952 50376 74016
rect 50440 73952 50456 74016
rect 50520 73952 50536 74016
rect 50600 73952 50608 74016
rect 50288 72928 50608 73952
rect 50288 72864 50296 72928
rect 50360 72864 50376 72928
rect 50440 72864 50456 72928
rect 50520 72864 50536 72928
rect 50600 72864 50608 72928
rect 50288 71840 50608 72864
rect 50288 71776 50296 71840
rect 50360 71776 50376 71840
rect 50440 71776 50456 71840
rect 50520 71776 50536 71840
rect 50600 71776 50608 71840
rect 50288 70752 50608 71776
rect 50288 70688 50296 70752
rect 50360 70688 50376 70752
rect 50440 70688 50456 70752
rect 50520 70688 50536 70752
rect 50600 70688 50608 70752
rect 50288 69664 50608 70688
rect 50288 69600 50296 69664
rect 50360 69600 50376 69664
rect 50440 69600 50456 69664
rect 50520 69600 50536 69664
rect 50600 69600 50608 69664
rect 50288 68576 50608 69600
rect 50288 68512 50296 68576
rect 50360 68512 50376 68576
rect 50440 68512 50456 68576
rect 50520 68512 50536 68576
rect 50600 68512 50608 68576
rect 50288 67488 50608 68512
rect 50288 67424 50296 67488
rect 50360 67424 50376 67488
rect 50440 67424 50456 67488
rect 50520 67424 50536 67488
rect 50600 67424 50608 67488
rect 50288 66400 50608 67424
rect 50288 66336 50296 66400
rect 50360 66336 50376 66400
rect 50440 66336 50456 66400
rect 50520 66336 50536 66400
rect 50600 66336 50608 66400
rect 50288 65312 50608 66336
rect 50288 65248 50296 65312
rect 50360 65248 50376 65312
rect 50440 65248 50456 65312
rect 50520 65248 50536 65312
rect 50600 65248 50608 65312
rect 50288 64224 50608 65248
rect 50288 64160 50296 64224
rect 50360 64160 50376 64224
rect 50440 64160 50456 64224
rect 50520 64160 50536 64224
rect 50600 64160 50608 64224
rect 50288 63136 50608 64160
rect 50288 63072 50296 63136
rect 50360 63072 50376 63136
rect 50440 63072 50456 63136
rect 50520 63072 50536 63136
rect 50600 63072 50608 63136
rect 50288 62048 50608 63072
rect 50288 61984 50296 62048
rect 50360 61984 50376 62048
rect 50440 61984 50456 62048
rect 50520 61984 50536 62048
rect 50600 61984 50608 62048
rect 50288 60960 50608 61984
rect 50288 60896 50296 60960
rect 50360 60896 50376 60960
rect 50440 60896 50456 60960
rect 50520 60896 50536 60960
rect 50600 60896 50608 60960
rect 50288 59872 50608 60896
rect 50288 59808 50296 59872
rect 50360 59808 50376 59872
rect 50440 59808 50456 59872
rect 50520 59808 50536 59872
rect 50600 59808 50608 59872
rect 50288 58784 50608 59808
rect 50288 58720 50296 58784
rect 50360 58720 50376 58784
rect 50440 58720 50456 58784
rect 50520 58720 50536 58784
rect 50600 58720 50608 58784
rect 50288 57696 50608 58720
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 77824 65968 77840
rect 65648 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65968 77824
rect 65648 76736 65968 77760
rect 65648 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65968 76736
rect 65648 75648 65968 76672
rect 65648 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65968 75648
rect 65648 74560 65968 75584
rect 65648 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65968 74560
rect 65648 73472 65968 74496
rect 65648 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65968 73472
rect 65648 72384 65968 73408
rect 65648 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65968 72384
rect 65648 71296 65968 72320
rect 65648 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65968 71296
rect 65648 70208 65968 71232
rect 65648 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65968 70208
rect 65648 69120 65968 70144
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 68032 65968 69056
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65968 66944
rect 65648 65856 65968 66880
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 64768 65968 65792
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 63680 65968 64704
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 62592 65968 63616
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 61504 65968 62528
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 60416 65968 61440
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 59328 65968 60352
rect 65648 59264 65656 59328
rect 65720 59264 65736 59328
rect 65800 59264 65816 59328
rect 65880 59264 65896 59328
rect 65960 59264 65968 59328
rect 65648 58240 65968 59264
rect 65648 58176 65656 58240
rect 65720 58176 65736 58240
rect 65800 58176 65816 58240
rect 65880 58176 65896 58240
rect 65960 58176 65968 58240
rect 65648 57152 65968 58176
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__029__A pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30728 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__029__B
timestamp 1649977179
transform 1 0 30544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__029__C
timestamp 1649977179
transform 1 0 29992 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__029__D
timestamp 1649977179
transform 1 0 30544 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__030__A
timestamp 1649977179
transform 1 0 30268 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__030__B
timestamp 1649977179
transform 1 0 30820 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__030__C_N
timestamp 1649977179
transform 1 0 31004 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__030__D_N
timestamp 1649977179
transform 1 0 30820 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__032__A
timestamp 1649977179
transform 1 0 25760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__032__B
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__032__C
timestamp 1649977179
transform 1 0 26312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__033__A
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__033__B
timestamp 1649977179
transform 1 0 26312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__033__C
timestamp 1649977179
transform 1 0 26128 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__033__D
timestamp 1649977179
transform 1 0 25760 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__034__A
timestamp 1649977179
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__034__B
timestamp 1649977179
transform 1 0 26864 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__034__C
timestamp 1649977179
transform 1 0 26312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__034__D
timestamp 1649977179
transform 1 0 26496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__036__A_N
timestamp 1649977179
transform 1 0 40848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__036__C
timestamp 1649977179
transform 1 0 40664 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__037__A
timestamp 1649977179
transform 1 0 60536 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__039__A
timestamp 1649977179
transform 1 0 41124 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__039__C
timestamp 1649977179
transform -1 0 41860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__040__A
timestamp 1649977179
transform 1 0 61088 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__042__A1
timestamp 1649977179
transform 1 0 53912 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__042__B2
timestamp 1649977179
transform -1 0 52900 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__043__A1
timestamp 1649977179
transform -1 0 51428 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__043__B2
timestamp 1649977179
transform -1 0 49772 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__044__A1
timestamp 1649977179
transform -1 0 51428 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__044__B2
timestamp 1649977179
transform -1 0 49680 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__045__A1
timestamp 1649977179
transform -1 0 51612 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__045__B2
timestamp 1649977179
transform -1 0 49956 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__046__A1
timestamp 1649977179
transform 1 0 51888 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__046__B2
timestamp 1649977179
transform 1 0 50232 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__049__A1
timestamp 1649977179
transform -1 0 54372 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__049__B2
timestamp 1649977179
transform -1 0 51428 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__050__A1
timestamp 1649977179
transform -1 0 55660 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__050__B2
timestamp 1649977179
transform -1 0 54832 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__051__A1
timestamp 1649977179
transform -1 0 53912 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__051__B2
timestamp 1649977179
transform -1 0 52992 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__052__A1
timestamp 1649977179
transform 1 0 52256 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__052__B2
timestamp 1649977179
transform -1 0 51152 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__053__A1
timestamp 1649977179
transform -1 0 55384 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__053__B2
timestamp 1649977179
transform -1 0 54464 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A1
timestamp 1649977179
transform -1 0 57316 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__B2
timestamp 1649977179
transform -1 0 55660 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__A1
timestamp 1649977179
transform -1 0 57132 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__B2
timestamp 1649977179
transform -1 0 55844 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A1
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__B2
timestamp 1649977179
transform 1 0 55936 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A1
timestamp 1649977179
transform 1 0 58420 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__B2
timestamp 1649977179
transform -1 0 58880 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A1
timestamp 1649977179
transform -1 0 59064 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__B2
timestamp 1649977179
transform -1 0 59156 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A1
timestamp 1649977179
transform -1 0 58420 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__B2
timestamp 1649977179
transform -1 0 58972 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A1
timestamp 1649977179
transform -1 0 61364 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__B2
timestamp 1649977179
transform -1 0 61272 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A1
timestamp 1649977179
transform 1 0 60628 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__B2
timestamp 1649977179
transform 1 0 59800 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A1
timestamp 1649977179
transform -1 0 59616 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__B2
timestamp 1649977179
transform 1 0 58696 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A1
timestamp 1649977179
transform -1 0 59524 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__B2
timestamp 1649977179
transform 1 0 58696 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A1
timestamp 1649977179
transform 1 0 62376 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__B2
timestamp 1649977179
transform -1 0 63204 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A1
timestamp 1649977179
transform -1 0 64308 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__B2
timestamp 1649977179
transform -1 0 63204 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A1
timestamp 1649977179
transform 1 0 64492 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__B2
timestamp 1649977179
transform -1 0 63756 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A1
timestamp 1649977179
transform 1 0 62560 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__B2
timestamp 1649977179
transform 1 0 61640 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A1
timestamp 1649977179
transform 1 0 63940 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__B2
timestamp 1649977179
transform -1 0 62284 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform 1 0 65412 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1649977179
transform -1 0 66424 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A1
timestamp 1649977179
transform -1 0 67344 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__B2
timestamp 1649977179
transform -1 0 66148 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A1
timestamp 1649977179
transform 1 0 67528 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__B2
timestamp 1649977179
transform -1 0 64676 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A1
timestamp 1649977179
transform 1 0 65596 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__B2
timestamp 1649977179
transform -1 0 65228 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A1
timestamp 1649977179
transform -1 0 66792 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__B2
timestamp 1649977179
transform 1 0 63112 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A1
timestamp 1649977179
transform -1 0 66700 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B2
timestamp 1649977179
transform -1 0 65780 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform -1 0 66976 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform -1 0 63204 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A1
timestamp 1649977179
transform 1 0 67344 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__B2
timestamp 1649977179
transform -1 0 66332 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A1
timestamp 1649977179
transform 1 0 68632 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__B2
timestamp 1649977179
transform -1 0 68264 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A1
timestamp 1649977179
transform 1 0 65596 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B2
timestamp 1649977179
transform 1 0 64216 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform 1 0 67344 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1649977179
transform -1 0 66884 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform -1 0 62560 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform -1 0 62192 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1649977179
transform 1 0 41492 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1649977179
transform 1 0 27600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform -1 0 26864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1649977179
transform 1 0 26312 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1649977179
transform -1 0 28336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform 1 0 26680 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1649977179
transform 1 0 26312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 32292 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1649977179
transform 1 0 31464 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1649977179
transform -1 0 31096 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1649977179
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform -1 0 27324 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1649977179
transform -1 0 27508 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform 1 0 27140 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1649977179
transform -1 0 27324 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform -1 0 33028 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1649977179
transform -1 0 31556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform -1 0 32108 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1649977179
transform -1 0 32568 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1649977179
transform -1 0 12328 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1649977179
transform 1 0 12144 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1649977179
transform 1 0 14076 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1649977179
transform 1 0 12972 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1649977179
transform 1 0 15088 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1649977179
transform -1 0 15640 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A
timestamp 1649977179
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1649977179
transform 1 0 17296 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1649977179
transform -1 0 17848 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1649977179
transform -1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1649977179
transform 1 0 19688 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1649977179
transform 1 0 20608 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1649977179
transform -1 0 20516 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1649977179
transform 1 0 22448 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1649977179
transform -1 0 23092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1649977179
transform -1 0 23092 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1649977179
transform 1 0 23552 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1649977179
transform -1 0 26220 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1649977179
transform 1 0 27324 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A
timestamp 1649977179
transform 1 0 27876 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A
timestamp 1649977179
transform -1 0 28336 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1649977179
transform 1 0 28888 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A
timestamp 1649977179
transform 1 0 30636 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1649977179
transform 1 0 31924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1649977179
transform -1 0 33028 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1649977179
transform -1 0 32844 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A
timestamp 1649977179
transform 1 0 33396 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1649977179
transform -1 0 34224 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A
timestamp 1649977179
transform -1 0 35604 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1649977179
transform -1 0 35696 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1649977179
transform 1 0 36248 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A
timestamp 1649977179
transform 1 0 37168 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 1649977179
transform -1 0 38180 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A
timestamp 1649977179
transform -1 0 38548 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A
timestamp 1649977179
transform 1 0 40020 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 1649977179
transform 1 0 40756 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A
timestamp 1649977179
transform 1 0 41492 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__A
timestamp 1649977179
transform -1 0 42780 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A
timestamp 1649977179
transform -1 0 44068 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__A
timestamp 1649977179
transform -1 0 44528 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1649977179
transform -1 0 44528 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__A
timestamp 1649977179
transform -1 0 46000 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1649977179
transform 1 0 46368 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__187__A
timestamp 1649977179
transform -1 0 47748 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1649977179
transform -1 0 48208 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1649977179
transform -1 0 48944 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1649977179
transform -1 0 49680 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 1649977179
transform 1 0 25484 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A
timestamp 1649977179
transform -1 0 26496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1649977179
transform 1 0 27324 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1649977179
transform -1 0 27048 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1649977179
transform -1 0 27784 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1649977179
transform -1 0 29256 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A
timestamp 1649977179
transform 1 0 29992 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1649977179
transform -1 0 29992 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 1649977179
transform 1 0 31464 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1649977179
transform -1 0 33120 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A
timestamp 1649977179
transform -1 0 34500 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__A
timestamp 1649977179
transform -1 0 32936 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1649977179
transform -1 0 33672 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A
timestamp 1649977179
transform 1 0 35696 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1649977179
transform -1 0 35144 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A
timestamp 1649977179
transform -1 0 35788 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1649977179
transform -1 0 36524 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1649977179
transform 1 0 38548 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A
timestamp 1649977179
transform -1 0 37996 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1649977179
transform -1 0 38640 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1649977179
transform -1 0 39468 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1649977179
transform -1 0 41124 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1649977179
transform 1 0 42964 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A
timestamp 1649977179
transform -1 0 42320 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1649977179
transform -1 0 43976 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1649977179
transform -1 0 43792 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1649977179
transform -1 0 46736 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1649977179
transform -1 0 45172 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1649977179
transform -1 0 46828 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1649977179
transform -1 0 48208 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1649977179
transform -1 0 74704 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A
timestamp 1649977179
transform -1 0 75440 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1649977179
transform -1 0 76728 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1649977179
transform -1 0 76820 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1649977179
transform -1 0 71668 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1649977179
transform 1 0 71852 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1649977179
transform -1 0 72680 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A
timestamp 1649977179
transform 1 0 73324 0 -1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__231__A
timestamp 1649977179
transform -1 0 73968 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__A
timestamp 1649977179
transform -1 0 70932 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 78200 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 1564 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 1748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 9844 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 10488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 12420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 14904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 15640 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 16192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 17572 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 18124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 18676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 20056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 20792 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 21344 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 21988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 22724 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 23276 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 4416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 23828 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 25208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 7268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 7820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 8372 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 78200 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 76728 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 77556 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 77372 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 77556 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 78200 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 77372 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 77556 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 77372 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 77556 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 77556 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 77372 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 78016 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 77556 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 78200 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 77372 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 77556 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 77372 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 77556 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 77556 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 77372 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 77556 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 78200 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 77464 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 77372 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 77556 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 76728 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 76912 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 78200 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 77648 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 76912 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 77556 0 1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 78016 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 2300 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 2300 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 2300 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 2300 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 1564 0 1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 2300 0 -1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 2300 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 2300 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 1564 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 2300 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 2300 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 1564 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 2300 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 1564 0 1 63104
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 2300 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 2300 0 1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 2300 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 1564 0 -1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 2300 0 1 66368
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 2300 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 2300 0 1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1649977179
transform -1 0 1564 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1649977179
transform -1 0 2300 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1649977179
transform -1 0 2300 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1649977179
transform -1 0 2300 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1649977179
transform -1 0 2300 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1649977179
transform -1 0 2300 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1649977179
transform -1 0 1564 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1649977179
transform -1 0 2300 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1649977179
transform -1 0 2300 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1649977179
transform -1 0 2300 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1649977179
transform -1 0 1564 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1649977179
transform -1 0 27140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1649977179
transform -1 0 33028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1649977179
transform -1 0 33764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1649977179
transform -1 0 34132 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1649977179
transform -1 0 35512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1649977179
transform -1 0 36248 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1649977179
transform -1 0 36800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1649977179
transform -1 0 37444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1649977179
transform -1 0 38732 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1649977179
transform -1 0 39284 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1649977179
transform -1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1649977179
transform -1 0 40020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1649977179
transform -1 0 41124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1649977179
transform -1 0 42596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1649977179
transform -1 0 43148 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1649977179
transform -1 0 43884 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1649977179
transform -1 0 43700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1649977179
transform -1 0 44988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1649977179
transform -1 0 45724 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1649977179
transform -1 0 46460 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1649977179
transform -1 0 47748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1649977179
transform -1 0 26772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1649977179
transform -1 0 48300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1649977179
transform -1 0 48852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1649977179
transform -1 0 28612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1649977179
transform -1 0 29716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1649977179
transform -1 0 30636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1649977179
transform -1 0 30084 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1649977179
transform -1 0 30360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1649977179
transform -1 0 31648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1649977179
transform -1 0 32292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1649977179
transform -1 0 74060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1649977179
transform -1 0 74796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1649977179
transform -1 0 74612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1649977179
transform -1 0 75900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1649977179
transform -1 0 76636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input137_A
timestamp 1649977179
transform -1 0 73508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output138_A
timestamp 1649977179
transform 1 0 77096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output139_A
timestamp 1649977179
transform 1 0 77096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output140_A
timestamp 1649977179
transform -1 0 77464 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output141_A
timestamp 1649977179
transform 1 0 77096 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output142_A
timestamp 1649977179
transform -1 0 77464 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output143_A
timestamp 1649977179
transform -1 0 77280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output144_A
timestamp 1649977179
transform 1 0 77096 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output145_A
timestamp 1649977179
transform -1 0 77464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1649977179
transform -1 0 77280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output147_A
timestamp 1649977179
transform -1 0 77464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output148_A
timestamp 1649977179
transform -1 0 77464 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output149_A
timestamp 1649977179
transform 1 0 77096 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output150_A
timestamp 1649977179
transform -1 0 77464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output151_A
timestamp 1649977179
transform -1 0 77464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output152_A
timestamp 1649977179
transform -1 0 77280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output153_A
timestamp 1649977179
transform 1 0 77096 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output154_A
timestamp 1649977179
transform -1 0 77464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output155_A
timestamp 1649977179
transform 1 0 77096 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output156_A
timestamp 1649977179
transform -1 0 77464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output157_A
timestamp 1649977179
transform -1 0 77464 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output158_A
timestamp 1649977179
transform 1 0 77096 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output159_A
timestamp 1649977179
transform -1 0 77464 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output160_A
timestamp 1649977179
transform 1 0 77096 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output161_A
timestamp 1649977179
transform -1 0 77464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output162_A
timestamp 1649977179
transform 1 0 77096 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output163_A
timestamp 1649977179
transform -1 0 77464 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output164_A
timestamp 1649977179
transform 1 0 77096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output165_A
timestamp 1649977179
transform -1 0 77464 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output166_A
timestamp 1649977179
transform 1 0 77096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output167_A
timestamp 1649977179
transform 1 0 77096 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output168_A
timestamp 1649977179
transform -1 0 77464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output169_A
timestamp 1649977179
transform 1 0 77096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output170_A
timestamp 1649977179
transform -1 0 77464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output189_A
timestamp 1649977179
transform -1 0 2300 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output190_A
timestamp 1649977179
transform 1 0 2116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output191_A
timestamp 1649977179
transform -1 0 2300 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output192_A
timestamp 1649977179
transform 1 0 2116 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output194_A
timestamp 1649977179
transform 1 0 2116 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output195_A
timestamp 1649977179
transform -1 0 2300 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output203_A
timestamp 1649977179
transform -1 0 77464 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output204_A
timestamp 1649977179
transform -1 0 2300 0 1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output205_A
timestamp 1649977179
transform -1 0 50140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output206_A
timestamp 1649977179
transform -1 0 57316 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output207_A
timestamp 1649977179
transform -1 0 58052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output208_A
timestamp 1649977179
transform 1 0 58420 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output209_A
timestamp 1649977179
transform 1 0 58972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output210_A
timestamp 1649977179
transform -1 0 60444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output211_A
timestamp 1649977179
transform 1 0 60812 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output212_A
timestamp 1649977179
transform -1 0 61548 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output213_A
timestamp 1649977179
transform -1 0 62100 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output214_A
timestamp 1649977179
transform -1 0 63204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output215_A
timestamp 1649977179
transform 1 0 63572 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output216_A
timestamp 1649977179
transform 1 0 50508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output217_A
timestamp 1649977179
transform 1 0 64308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output218_A
timestamp 1649977179
transform -1 0 64308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output219_A
timestamp 1649977179
transform 1 0 65412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output220_A
timestamp 1649977179
transform 1 0 66148 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output221_A
timestamp 1649977179
transform 1 0 66884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output222_A
timestamp 1649977179
transform -1 0 68356 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output223_A
timestamp 1649977179
transform 1 0 68724 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output224_A
timestamp 1649977179
transform 1 0 69460 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output225_A
timestamp 1649977179
transform -1 0 69460 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output226_A
timestamp 1649977179
transform 1 0 70564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output227_A
timestamp 1649977179
transform -1 0 51428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output228_A
timestamp 1649977179
transform 1 0 71300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output229_A
timestamp 1649977179
transform 1 0 72036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output230_A
timestamp 1649977179
transform -1 0 51980 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output231_A
timestamp 1649977179
transform -1 0 52900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output232_A
timestamp 1649977179
transform 1 0 53820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output233_A
timestamp 1649977179
transform -1 0 53452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output234_A
timestamp 1649977179
transform -1 0 54004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output235_A
timestamp 1649977179
transform 1 0 55108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output236_A
timestamp 1649977179
transform 1 0 56396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output237_A
timestamp 1649977179
transform 1 0 77096 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output238_A
timestamp 1649977179
transform -1 0 77464 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output239_A
timestamp 1649977179
transform 1 0 77096 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output240_A
timestamp 1649977179
transform -1 0 77464 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output241_A
timestamp 1649977179
transform 1 0 77096 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output242_A
timestamp 1649977179
transform 1 0 77096 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output243_A
timestamp 1649977179
transform -1 0 77464 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output244_A
timestamp 1649977179
transform 1 0 77096 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output245_A
timestamp 1649977179
transform -1 0 77464 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output246_A
timestamp 1649977179
transform -1 0 77464 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output247_A
timestamp 1649977179
transform 1 0 77096 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output248_A
timestamp 1649977179
transform -1 0 77464 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output249_A
timestamp 1649977179
transform -1 0 77464 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output250_A
timestamp 1649977179
transform 1 0 77096 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output251_A
timestamp 1649977179
transform 1 0 77096 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output252_A
timestamp 1649977179
transform -1 0 77464 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output253_A
timestamp 1649977179
transform 1 0 77096 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output254_A
timestamp 1649977179
transform -1 0 77464 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output255_A
timestamp 1649977179
transform -1 0 77464 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output256_A
timestamp 1649977179
transform 1 0 77096 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output257_A
timestamp 1649977179
transform -1 0 77464 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output258_A
timestamp 1649977179
transform 1 0 77096 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output259_A
timestamp 1649977179
transform -1 0 77464 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output260_A
timestamp 1649977179
transform 1 0 77096 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output261_A
timestamp 1649977179
transform -1 0 77464 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output262_A
timestamp 1649977179
transform 1 0 77096 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output263_A
timestamp 1649977179
transform -1 0 77464 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output264_A
timestamp 1649977179
transform 1 0 77096 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output265_A
timestamp 1649977179
transform 1 0 77096 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output266_A
timestamp 1649977179
transform -1 0 77464 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output267_A
timestamp 1649977179
transform 1 0 77096 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output268_A
timestamp 1649977179
transform -1 0 77464 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output269_A
timestamp 1649977179
transform 1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output270_A
timestamp 1649977179
transform -1 0 2300 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output271_A
timestamp 1649977179
transform 1 0 2116 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output272_A
timestamp 1649977179
transform -1 0 2300 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output273_A
timestamp 1649977179
transform 1 0 2116 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output274_A
timestamp 1649977179
transform 1 0 2116 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output275_A
timestamp 1649977179
transform -1 0 2300 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output276_A
timestamp 1649977179
transform 1 0 2116 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output277_A
timestamp 1649977179
transform -1 0 2300 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output278_A
timestamp 1649977179
transform -1 0 2300 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output279_A
timestamp 1649977179
transform 1 0 2116 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output280_A
timestamp 1649977179
transform -1 0 2300 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output281_A
timestamp 1649977179
transform -1 0 2300 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output282_A
timestamp 1649977179
transform 1 0 2116 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output283_A
timestamp 1649977179
transform 1 0 2116 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output284_A
timestamp 1649977179
transform -1 0 2300 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output285_A
timestamp 1649977179
transform 1 0 2116 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output286_A
timestamp 1649977179
transform -1 0 2300 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output287_A
timestamp 1649977179
transform -1 0 2300 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output288_A
timestamp 1649977179
transform 1 0 2116 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output289_A
timestamp 1649977179
transform -1 0 2300 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output290_A
timestamp 1649977179
transform 1 0 2116 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output291_A
timestamp 1649977179
transform -1 0 2300 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output292_A
timestamp 1649977179
transform 1 0 2116 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output293_A
timestamp 1649977179
transform -1 0 2300 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output294_A
timestamp 1649977179
transform 1 0 2116 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output295_A
timestamp 1649977179
transform -1 0 2300 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output296_A
timestamp 1649977179
transform 1 0 2116 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output297_A
timestamp 1649977179
transform 1 0 2116 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output298_A
timestamp 1649977179
transform -1 0 2300 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output299_A
timestamp 1649977179
transform 1 0 2116 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output300_A
timestamp 1649977179
transform -1 0 2300 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output305_A
timestamp 1649977179
transform -1 0 2300 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output306_A
timestamp 1649977179
transform -1 0 2300 0 1 71808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output307_A
timestamp 1649977179
transform 1 0 2116 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output308_A
timestamp 1649977179
transform -1 0 2300 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output309_A
timestamp 1649977179
transform 1 0 77096 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output310_A
timestamp 1649977179
transform 1 0 2116 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output312_A
timestamp 1649977179
transform 1 0 2116 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14
timestamp 1649977179
transform 1 0 2392 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31
timestamp 1649977179
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1649977179
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1649977179
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70
timestamp 1649977179
transform 1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1649977179
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 1649977179
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1649977179
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1649977179
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_183
timestamp 1649977179
transform 1 0 17940 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1649977179
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1649977179
transform 1 0 19872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_231
timestamp 1649977179
transform 1 0 22356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_239
timestamp 1649977179
transform 1 0 23092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1649977179
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1649977179
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_257
timestamp 1649977179
transform 1 0 24748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_283 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27140 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_291
timestamp 1649977179
transform 1 0 27876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_311
timestamp 1649977179
transform 1 0 29716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_315
timestamp 1649977179
transform 1 0 30084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_318
timestamp 1649977179
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_347
timestamp 1649977179
transform 1 0 33028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1649977179
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1649977179
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_372
timestamp 1649977179
transform 1 0 35328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_380
timestamp 1649977179
transform 1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1649977179
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_399
timestamp 1649977179
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_407
timestamp 1649977179
transform 1 0 38548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_415
timestamp 1649977179
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1649977179
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_423
timestamp 1649977179
transform 1 0 40020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_439
timestamp 1649977179
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1649977179
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_453
timestamp 1649977179
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1649977179
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_469
timestamp 1649977179
transform 1 0 44252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1649977179
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_481
timestamp 1649977179
transform 1 0 45356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1649977179
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_497
timestamp 1649977179
transform 1 0 46828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1649977179
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_509
timestamp 1649977179
transform 1 0 47932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_517
timestamp 1649977179
transform 1 0 48668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_525
timestamp 1649977179
transform 1 0 49404 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1649977179
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_537
timestamp 1649977179
transform 1 0 50508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_545
timestamp 1649977179
transform 1 0 51244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_553
timestamp 1649977179
transform 1 0 51980 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_559
timestamp 1649977179
transform 1 0 52532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_565
timestamp 1649977179
transform 1 0 53084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_573
timestamp 1649977179
transform 1 0 53820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_581
timestamp 1649977179
transform 1 0 54556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1649977179
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_593
timestamp 1649977179
transform 1 0 55660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_601
timestamp 1649977179
transform 1 0 56396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_609
timestamp 1649977179
transform 1 0 57132 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1649977179
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1649977179
transform 1 0 58236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_629
timestamp 1649977179
transform 1 0 58972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_637
timestamp 1649977179
transform 1 0 59708 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_643
timestamp 1649977179
transform 1 0 60260 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_649
timestamp 1649977179
transform 1 0 60812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_657
timestamp 1649977179
transform 1 0 61548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_665
timestamp 1649977179
transform 1 0 62284 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_671
timestamp 1649977179
transform 1 0 62836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_677
timestamp 1649977179
transform 1 0 63388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_685
timestamp 1649977179
transform 1 0 64124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_693
timestamp 1649977179
transform 1 0 64860 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_699
timestamp 1649977179
transform 1 0 65412 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_705
timestamp 1649977179
transform 1 0 65964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_713
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_721
timestamp 1649977179
transform 1 0 67436 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_727
timestamp 1649977179
transform 1 0 67988 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_733
timestamp 1649977179
transform 1 0 68540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_741
timestamp 1649977179
transform 1 0 69276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_749
timestamp 1649977179
transform 1 0 70012 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_755
timestamp 1649977179
transform 1 0 70564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_761
timestamp 1649977179
transform 1 0 71116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_769
timestamp 1649977179
transform 1 0 71852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_777
timestamp 1649977179
transform 1 0 72588 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_783
timestamp 1649977179
transform 1 0 73140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_789
timestamp 1649977179
transform 1 0 73692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_797
timestamp 1649977179
transform 1 0 74428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_805
timestamp 1649977179
transform 1 0 75164 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_811
timestamp 1649977179
transform 1 0 75716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_817
timestamp 1649977179
transform 1 0 76268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_825
timestamp 1649977179
transform 1 0 77004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_833
timestamp 1649977179
transform 1 0 77740 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_839
timestamp 1649977179
transform 1 0 78292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_841
timestamp 1649977179
transform 1 0 78476 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_36
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1649977179
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_59
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_67
timestamp 1649977179
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1649977179
transform 1 0 8372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_86
timestamp 1649977179
transform 1 0 9016 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_92
timestamp 1649977179
transform 1 0 9568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_95
timestamp 1649977179
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_99
timestamp 1649977179
transform 1 0 10212 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_115
timestamp 1649977179
transform 1 0 11684 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1649977179
transform 1 0 12420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_147
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_150
timestamp 1649977179
transform 1 0 14904 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_171
timestamp 1649977179
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_179
timestamp 1649977179
transform 1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_191
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_203
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_214
timestamp 1649977179
transform 1 0 20792 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_227
timestamp 1649977179
transform 1 0 21988 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_235
timestamp 1649977179
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1649977179
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_259
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_283
timestamp 1649977179
transform 1 0 27140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_297
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_311
timestamp 1649977179
transform 1 0 29716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_325
timestamp 1649977179
transform 1 0 31004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_329
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_343
timestamp 1649977179
transform 1 0 32660 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_351
timestamp 1649977179
transform 1 0 33396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_359
timestamp 1649977179
transform 1 0 34132 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_367
timestamp 1649977179
transform 1 0 34868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_371
timestamp 1649977179
transform 1 0 35236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_374
timestamp 1649977179
transform 1 0 35512 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_382
timestamp 1649977179
transform 1 0 36248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1649977179
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_395
timestamp 1649977179
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_409
timestamp 1649977179
transform 1 0 38732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_415
timestamp 1649977179
transform 1 0 39284 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_423
timestamp 1649977179
transform 1 0 40020 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_435
timestamp 1649977179
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1649977179
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_451
timestamp 1649977179
transform 1 0 42596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_457
timestamp 1649977179
transform 1 0 43148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_463
timestamp 1649977179
transform 1 0 43700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_471
timestamp 1649977179
transform 1 0 44436 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_477
timestamp 1649977179
transform 1 0 44988 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_485
timestamp 1649977179
transform 1 0 45724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_493
timestamp 1649977179
transform 1 0 46460 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_501
timestamp 1649977179
transform 1 0 47196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_507
timestamp 1649977179
transform 1 0 47748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_513
timestamp 1649977179
transform 1 0 48300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_519
timestamp 1649977179
transform 1 0 48852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_527
timestamp 1649977179
transform 1 0 49588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_533
timestamp 1649977179
transform 1 0 50140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_539
timestamp 1649977179
transform 1 0 50692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_547
timestamp 1649977179
transform 1 0 51428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 1649977179
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1649977179
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_563
timestamp 1649977179
transform 1 0 52900 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_569
timestamp 1649977179
transform 1 0 53452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_575
timestamp 1649977179
transform 1 0 54004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_583
timestamp 1649977179
transform 1 0 54740 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_589
timestamp 1649977179
transform 1 0 55292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_603
timestamp 1649977179
transform 1 0 56580 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_611
timestamp 1649977179
transform 1 0 57316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1649977179
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_619
timestamp 1649977179
transform 1 0 58052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_625
timestamp 1649977179
transform 1 0 58604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_631
timestamp 1649977179
transform 1 0 59156 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_639
timestamp 1649977179
transform 1 0 59892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_645
timestamp 1649977179
transform 1 0 60444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_651
timestamp 1649977179
transform 1 0 60996 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_657
timestamp 1649977179
transform 1 0 61548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_663
timestamp 1649977179
transform 1 0 62100 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1649977179
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_675
timestamp 1649977179
transform 1 0 63204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_681
timestamp 1649977179
transform 1 0 63756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_687
timestamp 1649977179
transform 1 0 64308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_695
timestamp 1649977179
transform 1 0 65044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_701
timestamp 1649977179
transform 1 0 65596 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_709
timestamp 1649977179
transform 1 0 66332 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_717
timestamp 1649977179
transform 1 0 67068 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_725
timestamp 1649977179
transform 1 0 67804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_731
timestamp 1649977179
transform 1 0 68356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_737
timestamp 1649977179
transform 1 0 68908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_743
timestamp 1649977179
transform 1 0 69460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_751
timestamp 1649977179
transform 1 0 70196 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_757
timestamp 1649977179
transform 1 0 70748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_765
timestamp 1649977179
transform 1 0 71484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_773
timestamp 1649977179
transform 1 0 72220 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_781
timestamp 1649977179
transform 1 0 72956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_787
timestamp 1649977179
transform 1 0 73508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_793
timestamp 1649977179
transform 1 0 74060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_799
timestamp 1649977179
transform 1 0 74612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_807
timestamp 1649977179
transform 1 0 75348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_813
timestamp 1649977179
transform 1 0 75900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_821
timestamp 1649977179
transform 1 0 76636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_825
timestamp 1649977179
transform 1 0 77004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_828
timestamp 1649977179
transform 1 0 77280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_836
timestamp 1649977179
transform 1 0 78016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_841
timestamp 1649977179
transform 1 0 78476 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_279
timestamp 1649977179
transform 1 0 26772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_293
timestamp 1649977179
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_299
timestamp 1649977179
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_315
timestamp 1649977179
transform 1 0 30084 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_339
timestamp 1649977179
transform 1 0 32292 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_347
timestamp 1649977179
transform 1 0 33028 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_355
timestamp 1649977179
transform 1 0 33764 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1649977179
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1649977179
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_457
timestamp 1649977179
transform 1 0 43148 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_465
timestamp 1649977179
transform 1 0 43884 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_473
timestamp 1649977179
transform 1 0 44620 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1649977179
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1649977179
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1649977179
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1649977179
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_569
timestamp 1649977179
transform 1 0 53452 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_575
timestamp 1649977179
transform 1 0 54004 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1649977179
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1649977179
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1649977179
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1649977179
transform 1 0 58604 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 1649977179
transform 1 0 59708 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1649977179
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1649977179
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1649977179
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1649977179
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_681
timestamp 1649977179
transform 1 0 63756 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_689
timestamp 1649977179
transform 1 0 64492 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_697
timestamp 1649977179
transform 1 0 65228 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1649977179
transform 1 0 67804 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_737
timestamp 1649977179
transform 1 0 68908 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_745
timestamp 1649977179
transform 1 0 69644 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_753
timestamp 1649977179
transform 1 0 70380 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1649977179
transform 1 0 70748 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1649977179
transform 1 0 71852 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1649977179
transform 1 0 72956 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_793
timestamp 1649977179
transform 1 0 74060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_801
timestamp 1649977179
transform 1 0 74796 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_809
timestamp 1649977179
transform 1 0 75532 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1649977179
transform 1 0 75900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_825
timestamp 1649977179
transform 1 0 77004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_833
timestamp 1649977179
transform 1 0 77740 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_838
timestamp 1649977179
transform 1 0 78200 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1649977179
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1649977179
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1649977179
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1649977179
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1649977179
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1649977179
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1649977179
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 1649977179
transform 1 0 67436 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 1649977179
transform 1 0 67988 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1649977179
transform 1 0 69276 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1649977179
transform 1 0 70380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1649977179
transform 1 0 71484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 1649977179
transform 1 0 72588 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 1649977179
transform 1 0 73140 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1649977179
transform 1 0 73324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1649977179
transform 1 0 74428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1649977179
transform 1 0 75532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1649977179
transform 1 0 76636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 1649977179
transform 1 0 77740 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 1649977179
transform 1 0 78292 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_841
timestamp 1649977179
transform 1 0 78476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp 1649977179
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_57
timestamp 1649977179
transform 1 0 6348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_69
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_569
timestamp 1649977179
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1649977179
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_613
timestamp 1649977179
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_625
timestamp 1649977179
transform 1 0 58604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_637
timestamp 1649977179
transform 1 0 59708 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_643
timestamp 1649977179
transform 1 0 60260 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1649977179
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1649977179
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1649977179
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1649977179
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1649977179
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1649977179
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_737
timestamp 1649977179
transform 1 0 68908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_749
timestamp 1649977179
transform 1 0 70012 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_755
timestamp 1649977179
transform 1 0 70564 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1649977179
transform 1 0 70748 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1649977179
transform 1 0 71852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_781
timestamp 1649977179
transform 1 0 72956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_793
timestamp 1649977179
transform 1 0 74060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_805
timestamp 1649977179
transform 1 0 75164 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_811
timestamp 1649977179
transform 1 0 75716 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1649977179
transform 1 0 75900 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1649977179
transform 1 0 77004 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_837
timestamp 1649977179
transform 1 0 78108 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_841
timestamp 1649977179
transform 1 0 78476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_62
timestamp 1649977179
transform 1 0 6808 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_74
timestamp 1649977179
transform 1 0 7912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_86
timestamp 1649977179
transform 1 0 9016 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_98
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_573
timestamp 1649977179
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_585
timestamp 1649977179
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_597
timestamp 1649977179
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_609
timestamp 1649977179
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_615
timestamp 1649977179
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1649977179
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1649977179
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1649977179
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1649977179
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1649977179
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1649977179
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_741
timestamp 1649977179
transform 1 0 69276 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_753
timestamp 1649977179
transform 1 0 70380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_765
timestamp 1649977179
transform 1 0 71484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_777
timestamp 1649977179
transform 1 0 72588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_783
timestamp 1649977179
transform 1 0 73140 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_785
timestamp 1649977179
transform 1 0 73324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_797
timestamp 1649977179
transform 1 0 74428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_809
timestamp 1649977179
transform 1 0 75532 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_821
timestamp 1649977179
transform 1 0 76636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_825
timestamp 1649977179
transform 1 0 77004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_828
timestamp 1649977179
transform 1 0 77280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_836
timestamp 1649977179
transform 1 0 78016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_841
timestamp 1649977179
transform 1 0 78476 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1649977179
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1649977179
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1649977179
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_737
timestamp 1649977179
transform 1 0 68908 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_749
timestamp 1649977179
transform 1 0 70012 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_755
timestamp 1649977179
transform 1 0 70564 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_757
timestamp 1649977179
transform 1 0 70748 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_769
timestamp 1649977179
transform 1 0 71852 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_781
timestamp 1649977179
transform 1 0 72956 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_793
timestamp 1649977179
transform 1 0 74060 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_805
timestamp 1649977179
transform 1 0 75164 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_811
timestamp 1649977179
transform 1 0 75716 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_813
timestamp 1649977179
transform 1 0 75900 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_825
timestamp 1649977179
transform 1 0 77004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_830
timestamp 1649977179
transform 1 0 77464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_838
timestamp 1649977179
transform 1 0 78200 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_26
timestamp 1649977179
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_38
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1649977179
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_67
timestamp 1649977179
transform 1 0 7268 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_79
timestamp 1649977179
transform 1 0 8372 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_91
timestamp 1649977179
transform 1 0 9476 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1649977179
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1649977179
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_741
timestamp 1649977179
transform 1 0 69276 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_753
timestamp 1649977179
transform 1 0 70380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_765
timestamp 1649977179
transform 1 0 71484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_777
timestamp 1649977179
transform 1 0 72588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_783
timestamp 1649977179
transform 1 0 73140 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_785
timestamp 1649977179
transform 1 0 73324 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_797
timestamp 1649977179
transform 1 0 74428 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_809
timestamp 1649977179
transform 1 0 75532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_821
timestamp 1649977179
transform 1 0 76636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_833
timestamp 1649977179
transform 1 0 77740 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_839
timestamp 1649977179
transform 1 0 78292 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_841
timestamp 1649977179
transform 1 0 78476 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_7
timestamp 1649977179
transform 1 0 1748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_33
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_45
timestamp 1649977179
transform 1 0 5244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_57
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_73
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1649977179
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1649977179
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1649977179
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1649977179
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_737
timestamp 1649977179
transform 1 0 68908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_749
timestamp 1649977179
transform 1 0 70012 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_755
timestamp 1649977179
transform 1 0 70564 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_757
timestamp 1649977179
transform 1 0 70748 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_769
timestamp 1649977179
transform 1 0 71852 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_781
timestamp 1649977179
transform 1 0 72956 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_793
timestamp 1649977179
transform 1 0 74060 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_805
timestamp 1649977179
transform 1 0 75164 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_811
timestamp 1649977179
transform 1 0 75716 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_813
timestamp 1649977179
transform 1 0 75900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_825
timestamp 1649977179
transform 1 0 77004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_830
timestamp 1649977179
transform 1 0 77464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_838
timestamp 1649977179
transform 1 0 78200 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_19
timestamp 1649977179
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_31
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_40
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_79
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_91
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1649977179
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1649977179
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_741
timestamp 1649977179
transform 1 0 69276 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_753
timestamp 1649977179
transform 1 0 70380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_765
timestamp 1649977179
transform 1 0 71484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_777
timestamp 1649977179
transform 1 0 72588 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_783
timestamp 1649977179
transform 1 0 73140 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_785
timestamp 1649977179
transform 1 0 73324 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_797
timestamp 1649977179
transform 1 0 74428 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_809
timestamp 1649977179
transform 1 0 75532 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_821
timestamp 1649977179
transform 1 0 76636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_825
timestamp 1649977179
transform 1 0 77004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_828
timestamp 1649977179
transform 1 0 77280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_836
timestamp 1649977179
transform 1 0 78016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_841
timestamp 1649977179
transform 1 0 78476 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_7
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_48
timestamp 1649977179
transform 1 0 5520 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_60
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_72
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_113
timestamp 1649977179
transform 1 0 11500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_125
timestamp 1649977179
transform 1 0 12604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1649977179
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1649977179
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_737
timestamp 1649977179
transform 1 0 68908 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_749
timestamp 1649977179
transform 1 0 70012 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_755
timestamp 1649977179
transform 1 0 70564 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_757
timestamp 1649977179
transform 1 0 70748 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_769
timestamp 1649977179
transform 1 0 71852 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_781
timestamp 1649977179
transform 1 0 72956 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_793
timestamp 1649977179
transform 1 0 74060 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_805
timestamp 1649977179
transform 1 0 75164 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_811
timestamp 1649977179
transform 1 0 75716 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_813
timestamp 1649977179
transform 1 0 75900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_825
timestamp 1649977179
transform 1 0 77004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_830
timestamp 1649977179
transform 1 0 77464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_838
timestamp 1649977179
transform 1 0 78200 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1649977179
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_741
timestamp 1649977179
transform 1 0 69276 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_753
timestamp 1649977179
transform 1 0 70380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_765
timestamp 1649977179
transform 1 0 71484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_777
timestamp 1649977179
transform 1 0 72588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_783
timestamp 1649977179
transform 1 0 73140 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_785
timestamp 1649977179
transform 1 0 73324 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_797
timestamp 1649977179
transform 1 0 74428 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_809
timestamp 1649977179
transform 1 0 75532 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_821
timestamp 1649977179
transform 1 0 76636 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_825
timestamp 1649977179
transform 1 0 77004 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_828
timestamp 1649977179
transform 1 0 77280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_836
timestamp 1649977179
transform 1 0 78016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_841
timestamp 1649977179
transform 1 0 78476 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_56
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_68
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_93
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_105
timestamp 1649977179
transform 1 0 10764 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_117
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_129
timestamp 1649977179
transform 1 0 12972 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1649977179
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1649977179
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1649977179
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1649977179
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_737
timestamp 1649977179
transform 1 0 68908 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_749
timestamp 1649977179
transform 1 0 70012 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_755
timestamp 1649977179
transform 1 0 70564 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_757
timestamp 1649977179
transform 1 0 70748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_769
timestamp 1649977179
transform 1 0 71852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_781
timestamp 1649977179
transform 1 0 72956 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_793
timestamp 1649977179
transform 1 0 74060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_805
timestamp 1649977179
transform 1 0 75164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_811
timestamp 1649977179
transform 1 0 75716 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_813
timestamp 1649977179
transform 1 0 75900 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_825
timestamp 1649977179
transform 1 0 77004 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_837
timestamp 1649977179
transform 1 0 78108 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_841
timestamp 1649977179
transform 1 0 78476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_7
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_19
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_31
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_43
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_64
timestamp 1649977179
transform 1 0 6992 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_76
timestamp 1649977179
transform 1 0 8096 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_88
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_100
timestamp 1649977179
transform 1 0 10304 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1649977179
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1649977179
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1649977179
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1649977179
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1649977179
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1649977179
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1649977179
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1649977179
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1649977179
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_729
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_741
timestamp 1649977179
transform 1 0 69276 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_753
timestamp 1649977179
transform 1 0 70380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_765
timestamp 1649977179
transform 1 0 71484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_777
timestamp 1649977179
transform 1 0 72588 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_783
timestamp 1649977179
transform 1 0 73140 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_785
timestamp 1649977179
transform 1 0 73324 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_797
timestamp 1649977179
transform 1 0 74428 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_809
timestamp 1649977179
transform 1 0 75532 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_821
timestamp 1649977179
transform 1 0 76636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_825
timestamp 1649977179
transform 1 0 77004 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_828
timestamp 1649977179
transform 1 0 77280 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_836
timestamp 1649977179
transform 1 0 78016 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_841
timestamp 1649977179
transform 1 0 78476 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_7
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_69
timestamp 1649977179
transform 1 0 7452 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_73
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_81
timestamp 1649977179
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_103
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_108
timestamp 1649977179
transform 1 0 11040 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_120
timestamp 1649977179
transform 1 0 12144 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1649977179
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1649977179
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1649977179
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1649977179
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1649977179
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1649977179
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1649977179
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1649977179
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_737
timestamp 1649977179
transform 1 0 68908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_749
timestamp 1649977179
transform 1 0 70012 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_755
timestamp 1649977179
transform 1 0 70564 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_757
timestamp 1649977179
transform 1 0 70748 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_769
timestamp 1649977179
transform 1 0 71852 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_781
timestamp 1649977179
transform 1 0 72956 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_793
timestamp 1649977179
transform 1 0 74060 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_805
timestamp 1649977179
transform 1 0 75164 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_811
timestamp 1649977179
transform 1 0 75716 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_813
timestamp 1649977179
transform 1 0 75900 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_825
timestamp 1649977179
transform 1 0 77004 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_830
timestamp 1649977179
transform 1 0 77464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_838
timestamp 1649977179
transform 1 0 78200 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_7
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_19
timestamp 1649977179
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_31
timestamp 1649977179
transform 1 0 3956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_77
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_117
timestamp 1649977179
transform 1 0 11868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_129
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_141
timestamp 1649977179
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_153
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1649977179
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1649977179
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1649977179
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1649977179
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1649977179
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1649977179
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1649977179
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1649977179
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1649977179
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1649977179
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1649977179
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1649977179
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1649977179
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_741
timestamp 1649977179
transform 1 0 69276 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_753
timestamp 1649977179
transform 1 0 70380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_765
timestamp 1649977179
transform 1 0 71484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_777
timestamp 1649977179
transform 1 0 72588 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_783
timestamp 1649977179
transform 1 0 73140 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_785
timestamp 1649977179
transform 1 0 73324 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_797
timestamp 1649977179
transform 1 0 74428 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_809
timestamp 1649977179
transform 1 0 75532 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_821
timestamp 1649977179
transform 1 0 76636 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_825
timestamp 1649977179
transform 1 0 77004 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_828
timestamp 1649977179
transform 1 0 77280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_836
timestamp 1649977179
transform 1 0 78016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_841
timestamp 1649977179
transform 1 0 78476 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1649977179
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1649977179
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1649977179
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1649977179
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1649977179
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1649977179
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1649977179
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1649977179
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1649977179
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1649977179
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_725
timestamp 1649977179
transform 1 0 67804 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_737
timestamp 1649977179
transform 1 0 68908 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_749
timestamp 1649977179
transform 1 0 70012 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_755
timestamp 1649977179
transform 1 0 70564 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_757
timestamp 1649977179
transform 1 0 70748 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_769
timestamp 1649977179
transform 1 0 71852 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_781
timestamp 1649977179
transform 1 0 72956 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_793
timestamp 1649977179
transform 1 0 74060 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_805
timestamp 1649977179
transform 1 0 75164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_811
timestamp 1649977179
transform 1 0 75716 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_813
timestamp 1649977179
transform 1 0 75900 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_825
timestamp 1649977179
transform 1 0 77004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_830
timestamp 1649977179
transform 1 0 77464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_838
timestamp 1649977179
transform 1 0 78200 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_85
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_89
timestamp 1649977179
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1649977179
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_117
timestamp 1649977179
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_122
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_134
timestamp 1649977179
transform 1 0 13432 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_146
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1649977179
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1649977179
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1649977179
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1649977179
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1649977179
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1649977179
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1649977179
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1649977179
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1649977179
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_709
timestamp 1649977179
transform 1 0 66332 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_721
timestamp 1649977179
transform 1 0 67436 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_727
timestamp 1649977179
transform 1 0 67988 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_729
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_741
timestamp 1649977179
transform 1 0 69276 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_753
timestamp 1649977179
transform 1 0 70380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_765
timestamp 1649977179
transform 1 0 71484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_777
timestamp 1649977179
transform 1 0 72588 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_783
timestamp 1649977179
transform 1 0 73140 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_785
timestamp 1649977179
transform 1 0 73324 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_797
timestamp 1649977179
transform 1 0 74428 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_809
timestamp 1649977179
transform 1 0 75532 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_821
timestamp 1649977179
transform 1 0 76636 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_833
timestamp 1649977179
transform 1 0 77740 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_839
timestamp 1649977179
transform 1 0 78292 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_841
timestamp 1649977179
transform 1 0 78476 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_7
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_19
timestamp 1649977179
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_96
timestamp 1649977179
transform 1 0 9936 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_108
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1649977179
transform 1 0 12144 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_124
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_129
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1649977179
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1649977179
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1649977179
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1649977179
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1649977179
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1649977179
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1649977179
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1649977179
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1649977179
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1649977179
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_725
timestamp 1649977179
transform 1 0 67804 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_737
timestamp 1649977179
transform 1 0 68908 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_749
timestamp 1649977179
transform 1 0 70012 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_755
timestamp 1649977179
transform 1 0 70564 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_757
timestamp 1649977179
transform 1 0 70748 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_769
timestamp 1649977179
transform 1 0 71852 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_781
timestamp 1649977179
transform 1 0 72956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_793
timestamp 1649977179
transform 1 0 74060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_805
timestamp 1649977179
transform 1 0 75164 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_811
timestamp 1649977179
transform 1 0 75716 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_813
timestamp 1649977179
transform 1 0 75900 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_825
timestamp 1649977179
transform 1 0 77004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_830
timestamp 1649977179
transform 1 0 77464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_838
timestamp 1649977179
transform 1 0 78200 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_19
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_31
timestamp 1649977179
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_43
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1649977179
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1649977179
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1649977179
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1649977179
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1649977179
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1649977179
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1649977179
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1649977179
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1649977179
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1649977179
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1649977179
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1649977179
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_729
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_741
timestamp 1649977179
transform 1 0 69276 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_753
timestamp 1649977179
transform 1 0 70380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_765
timestamp 1649977179
transform 1 0 71484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_777
timestamp 1649977179
transform 1 0 72588 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_783
timestamp 1649977179
transform 1 0 73140 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_785
timestamp 1649977179
transform 1 0 73324 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_797
timestamp 1649977179
transform 1 0 74428 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_809
timestamp 1649977179
transform 1 0 75532 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_821
timestamp 1649977179
transform 1 0 76636 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_825
timestamp 1649977179
transform 1 0 77004 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_828
timestamp 1649977179
transform 1 0 77280 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_836
timestamp 1649977179
transform 1 0 78016 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_841
timestamp 1649977179
transform 1 0 78476 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_7
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_19
timestamp 1649977179
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1649977179
transform 1 0 9660 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_99
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_111
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_123
timestamp 1649977179
transform 1 0 12420 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1649977179
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_279
timestamp 1649977179
transform 1 0 26772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_287
timestamp 1649977179
transform 1 0 27508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_290
timestamp 1649977179
transform 1 0 27784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_302
timestamp 1649977179
transform 1 0 28888 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1649977179
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_441
timestamp 1649977179
transform 1 0 41676 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_449
timestamp 1649977179
transform 1 0 42412 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_461
timestamp 1649977179
transform 1 0 43516 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_473
timestamp 1649977179
transform 1 0 44620 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1649977179
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1649977179
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1649977179
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1649977179
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1649977179
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1649977179
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1649977179
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1649977179
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1649977179
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_725
timestamp 1649977179
transform 1 0 67804 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_737
timestamp 1649977179
transform 1 0 68908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_749
timestamp 1649977179
transform 1 0 70012 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_755
timestamp 1649977179
transform 1 0 70564 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_757
timestamp 1649977179
transform 1 0 70748 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_769
timestamp 1649977179
transform 1 0 71852 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_781
timestamp 1649977179
transform 1 0 72956 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_793
timestamp 1649977179
transform 1 0 74060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_805
timestamp 1649977179
transform 1 0 75164 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_811
timestamp 1649977179
transform 1 0 75716 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_813
timestamp 1649977179
transform 1 0 75900 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_825
timestamp 1649977179
transform 1 0 77004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_830
timestamp 1649977179
transform 1 0 77464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_838
timestamp 1649977179
transform 1 0 78200 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_19
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_31
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_43
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_127
timestamp 1649977179
transform 1 0 12788 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_139
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_151
timestamp 1649977179
transform 1 0 14996 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1649977179
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_267
timestamp 1649977179
transform 1 0 25668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_270
timestamp 1649977179
transform 1 0 25944 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1649977179
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_286
timestamp 1649977179
transform 1 0 27416 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_294
timestamp 1649977179
transform 1 0 28152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_306
timestamp 1649977179
transform 1 0 29256 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_318
timestamp 1649977179
transform 1 0 30360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1649977179
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1649977179
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1649977179
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1649977179
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1649977179
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1649977179
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1649977179
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1649977179
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1649977179
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1649977179
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1649977179
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1649977179
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_729
timestamp 1649977179
transform 1 0 68172 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_741
timestamp 1649977179
transform 1 0 69276 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_753
timestamp 1649977179
transform 1 0 70380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_765
timestamp 1649977179
transform 1 0 71484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_777
timestamp 1649977179
transform 1 0 72588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_783
timestamp 1649977179
transform 1 0 73140 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_785
timestamp 1649977179
transform 1 0 73324 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_797
timestamp 1649977179
transform 1 0 74428 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_809
timestamp 1649977179
transform 1 0 75532 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_821
timestamp 1649977179
transform 1 0 76636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_825
timestamp 1649977179
transform 1 0 77004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_828
timestamp 1649977179
transform 1 0 77280 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_836
timestamp 1649977179
transform 1 0 78016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_841
timestamp 1649977179
transform 1 0 78476 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_116
timestamp 1649977179
transform 1 0 11776 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_122
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_134
timestamp 1649977179
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1649977179
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_288
timestamp 1649977179
transform 1 0 27600 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_300
timestamp 1649977179
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1649977179
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1649977179
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1649977179
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1649977179
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1649977179
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1649977179
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1649977179
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1649977179
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1649977179
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1649977179
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1649977179
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1649977179
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1649977179
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1649977179
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1649977179
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_725
timestamp 1649977179
transform 1 0 67804 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_737
timestamp 1649977179
transform 1 0 68908 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_749
timestamp 1649977179
transform 1 0 70012 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_755
timestamp 1649977179
transform 1 0 70564 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_757
timestamp 1649977179
transform 1 0 70748 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_769
timestamp 1649977179
transform 1 0 71852 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_781
timestamp 1649977179
transform 1 0 72956 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_793
timestamp 1649977179
transform 1 0 74060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_805
timestamp 1649977179
transform 1 0 75164 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_811
timestamp 1649977179
transform 1 0 75716 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_813
timestamp 1649977179
transform 1 0 75900 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_825
timestamp 1649977179
transform 1 0 77004 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_837
timestamp 1649977179
transform 1 0 78108 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_841
timestamp 1649977179
transform 1 0 78476 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_19
timestamp 1649977179
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_31
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_116
timestamp 1649977179
transform 1 0 11776 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_122
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_134
timestamp 1649977179
transform 1 0 13432 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_146
timestamp 1649977179
transform 1 0 14536 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_158
timestamp 1649977179
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1649977179
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1649977179
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_285
timestamp 1649977179
transform 1 0 27324 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_290
timestamp 1649977179
transform 1 0 27784 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_302
timestamp 1649977179
transform 1 0 28888 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_314
timestamp 1649977179
transform 1 0 29992 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_326
timestamp 1649977179
transform 1 0 31096 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1649977179
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1649977179
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1649977179
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1649977179
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1649977179
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1649977179
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1649977179
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1649977179
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1649977179
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1649977179
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1649977179
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1649977179
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1649977179
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1649977179
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1649977179
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_729
timestamp 1649977179
transform 1 0 68172 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_741
timestamp 1649977179
transform 1 0 69276 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_753
timestamp 1649977179
transform 1 0 70380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_765
timestamp 1649977179
transform 1 0 71484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_777
timestamp 1649977179
transform 1 0 72588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_783
timestamp 1649977179
transform 1 0 73140 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_785
timestamp 1649977179
transform 1 0 73324 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_797
timestamp 1649977179
transform 1 0 74428 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_809
timestamp 1649977179
transform 1 0 75532 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_821
timestamp 1649977179
transform 1 0 76636 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_825
timestamp 1649977179
transform 1 0 77004 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_828
timestamp 1649977179
transform 1 0 77280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_836
timestamp 1649977179
transform 1 0 78016 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_841
timestamp 1649977179
transform 1 0 78476 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1649977179
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_131
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_279
timestamp 1649977179
transform 1 0 26772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_287
timestamp 1649977179
transform 1 0 27508 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_291
timestamp 1649977179
transform 1 0 27876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_303
timestamp 1649977179
transform 1 0 28980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1649977179
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1649977179
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1649977179
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1649977179
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1649977179
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1649977179
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1649977179
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1649977179
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1649977179
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1649977179
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1649977179
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_725
timestamp 1649977179
transform 1 0 67804 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_737
timestamp 1649977179
transform 1 0 68908 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_749
timestamp 1649977179
transform 1 0 70012 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_755
timestamp 1649977179
transform 1 0 70564 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_757
timestamp 1649977179
transform 1 0 70748 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_769
timestamp 1649977179
transform 1 0 71852 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_781
timestamp 1649977179
transform 1 0 72956 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_793
timestamp 1649977179
transform 1 0 74060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_805
timestamp 1649977179
transform 1 0 75164 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_811
timestamp 1649977179
transform 1 0 75716 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_813
timestamp 1649977179
transform 1 0 75900 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_825
timestamp 1649977179
transform 1 0 77004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_830
timestamp 1649977179
transform 1 0 77464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_838
timestamp 1649977179
transform 1 0 78200 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_19
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_31
timestamp 1649977179
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_43
timestamp 1649977179
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_133
timestamp 1649977179
transform 1 0 13340 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_143
timestamp 1649977179
transform 1 0 14260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_155
timestamp 1649977179
transform 1 0 15364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_267
timestamp 1649977179
transform 1 0 25668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_270
timestamp 1649977179
transform 1 0 25944 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1649977179
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_287
timestamp 1649977179
transform 1 0 27508 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_295
timestamp 1649977179
transform 1 0 28244 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_307
timestamp 1649977179
transform 1 0 29348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_319
timestamp 1649977179
transform 1 0 30452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1649977179
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1649977179
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1649977179
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1649977179
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1649977179
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1649977179
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1649977179
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1649977179
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1649977179
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1649977179
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1649977179
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1649977179
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_729
timestamp 1649977179
transform 1 0 68172 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_741
timestamp 1649977179
transform 1 0 69276 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_753
timestamp 1649977179
transform 1 0 70380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_765
timestamp 1649977179
transform 1 0 71484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_777
timestamp 1649977179
transform 1 0 72588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_783
timestamp 1649977179
transform 1 0 73140 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_785
timestamp 1649977179
transform 1 0 73324 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_797
timestamp 1649977179
transform 1 0 74428 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_809
timestamp 1649977179
transform 1 0 75532 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_821
timestamp 1649977179
transform 1 0 76636 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_825
timestamp 1649977179
transform 1 0 77004 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_828
timestamp 1649977179
transform 1 0 77280 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_836
timestamp 1649977179
transform 1 0 78016 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_841
timestamp 1649977179
transform 1 0 78476 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1649977179
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_271
timestamp 1649977179
transform 1 0 26036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_274
timestamp 1649977179
transform 1 0 26312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_280
timestamp 1649977179
transform 1 0 26864 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_288
timestamp 1649977179
transform 1 0 27600 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_296
timestamp 1649977179
transform 1 0 28336 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1649977179
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1649977179
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1649977179
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1649977179
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1649977179
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1649977179
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1649977179
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1649977179
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1649977179
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1649977179
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1649977179
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_725
timestamp 1649977179
transform 1 0 67804 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_737
timestamp 1649977179
transform 1 0 68908 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_749
timestamp 1649977179
transform 1 0 70012 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_755
timestamp 1649977179
transform 1 0 70564 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_757
timestamp 1649977179
transform 1 0 70748 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_769
timestamp 1649977179
transform 1 0 71852 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_781
timestamp 1649977179
transform 1 0 72956 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_793
timestamp 1649977179
transform 1 0 74060 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_805
timestamp 1649977179
transform 1 0 75164 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_811
timestamp 1649977179
transform 1 0 75716 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_813
timestamp 1649977179
transform 1 0 75900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_825
timestamp 1649977179
transform 1 0 77004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_830
timestamp 1649977179
transform 1 0 77464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_838
timestamp 1649977179
transform 1 0 78200 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1649977179
transform 1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_154
timestamp 1649977179
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1649977179
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_285
timestamp 1649977179
transform 1 0 27324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_290
timestamp 1649977179
transform 1 0 27784 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_296
timestamp 1649977179
transform 1 0 28336 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_308
timestamp 1649977179
transform 1 0 29440 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_320
timestamp 1649977179
transform 1 0 30544 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1649977179
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1649977179
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1649977179
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1649977179
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1649977179
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1649977179
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1649977179
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1649977179
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1649977179
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1649977179
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1649977179
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1649977179
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1649977179
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1649977179
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1649977179
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_729
timestamp 1649977179
transform 1 0 68172 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_741
timestamp 1649977179
transform 1 0 69276 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_753
timestamp 1649977179
transform 1 0 70380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_765
timestamp 1649977179
transform 1 0 71484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_777
timestamp 1649977179
transform 1 0 72588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_783
timestamp 1649977179
transform 1 0 73140 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_785
timestamp 1649977179
transform 1 0 73324 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_797
timestamp 1649977179
transform 1 0 74428 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_809
timestamp 1649977179
transform 1 0 75532 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_821
timestamp 1649977179
transform 1 0 76636 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_833
timestamp 1649977179
transform 1 0 77740 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_839
timestamp 1649977179
transform 1 0 78292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_841
timestamp 1649977179
transform 1 0 78476 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_152
timestamp 1649977179
transform 1 0 15088 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_158
timestamp 1649977179
transform 1 0 15640 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_170
timestamp 1649977179
transform 1 0 16744 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_182
timestamp 1649977179
transform 1 0 17848 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_273
timestamp 1649977179
transform 1 0 26220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_278
timestamp 1649977179
transform 1 0 26680 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_292
timestamp 1649977179
transform 1 0 27968 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_304
timestamp 1649977179
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1649977179
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1649977179
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1649977179
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1649977179
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1649977179
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1649977179
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_625
timestamp 1649977179
transform 1 0 58604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_637
timestamp 1649977179
transform 1 0 59708 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_643
timestamp 1649977179
transform 1 0 60260 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1649977179
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1649977179
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1649977179
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1649977179
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1649977179
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1649977179
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1649977179
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1649977179
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_725
timestamp 1649977179
transform 1 0 67804 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_737
timestamp 1649977179
transform 1 0 68908 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_749
timestamp 1649977179
transform 1 0 70012 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_755
timestamp 1649977179
transform 1 0 70564 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_757
timestamp 1649977179
transform 1 0 70748 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_769
timestamp 1649977179
transform 1 0 71852 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_781
timestamp 1649977179
transform 1 0 72956 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_793
timestamp 1649977179
transform 1 0 74060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_805
timestamp 1649977179
transform 1 0 75164 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_811
timestamp 1649977179
transform 1 0 75716 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_813
timestamp 1649977179
transform 1 0 75900 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_825
timestamp 1649977179
transform 1 0 77004 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_830
timestamp 1649977179
transform 1 0 77464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_838
timestamp 1649977179
transform 1 0 78200 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_19
timestamp 1649977179
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_31
timestamp 1649977179
transform 1 0 3956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1649977179
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_288
timestamp 1649977179
transform 1 0 27600 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_300
timestamp 1649977179
transform 1 0 28704 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_312
timestamp 1649977179
transform 1 0 29808 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_320
timestamp 1649977179
transform 1 0 30544 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_324
timestamp 1649977179
transform 1 0 30912 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_339
timestamp 1649977179
transform 1 0 32292 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_351
timestamp 1649977179
transform 1 0 33396 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_363
timestamp 1649977179
transform 1 0 34500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_375
timestamp 1649977179
transform 1 0 35604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_387
timestamp 1649977179
transform 1 0 36708 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1649977179
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1649977179
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1649977179
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1649977179
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1649977179
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1649977179
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1649977179
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1649977179
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1649977179
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1649977179
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1649977179
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1649977179
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1649977179
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_729
timestamp 1649977179
transform 1 0 68172 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_741
timestamp 1649977179
transform 1 0 69276 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_753
timestamp 1649977179
transform 1 0 70380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_765
timestamp 1649977179
transform 1 0 71484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_777
timestamp 1649977179
transform 1 0 72588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_783
timestamp 1649977179
transform 1 0 73140 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_785
timestamp 1649977179
transform 1 0 73324 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_797
timestamp 1649977179
transform 1 0 74428 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_809
timestamp 1649977179
transform 1 0 75532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_821
timestamp 1649977179
transform 1 0 76636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_825
timestamp 1649977179
transform 1 0 77004 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_828
timestamp 1649977179
transform 1 0 77280 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_836
timestamp 1649977179
transform 1 0 78016 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_841
timestamp 1649977179
transform 1 0 78476 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_19
timestamp 1649977179
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_161
timestamp 1649977179
transform 1 0 15916 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_166
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_172
timestamp 1649977179
transform 1 0 16928 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_184
timestamp 1649977179
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_273
timestamp 1649977179
transform 1 0 26220 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_276
timestamp 1649977179
transform 1 0 26496 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_282
timestamp 1649977179
transform 1 0 27048 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_294
timestamp 1649977179
transform 1 0 28152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1649977179
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_313
timestamp 1649977179
transform 1 0 29900 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_316
timestamp 1649977179
transform 1 0 30176 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_322
timestamp 1649977179
transform 1 0 30728 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_332
timestamp 1649977179
transform 1 0 31648 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_340
timestamp 1649977179
transform 1 0 32384 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_352
timestamp 1649977179
transform 1 0 33488 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1649977179
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1649977179
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1649977179
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1649977179
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1649977179
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1649977179
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1649977179
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1649977179
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1649977179
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1649977179
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1649977179
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1649977179
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1649977179
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1649977179
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1649977179
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1649977179
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_725
timestamp 1649977179
transform 1 0 67804 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_737
timestamp 1649977179
transform 1 0 68908 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_749
timestamp 1649977179
transform 1 0 70012 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_755
timestamp 1649977179
transform 1 0 70564 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_757
timestamp 1649977179
transform 1 0 70748 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_769
timestamp 1649977179
transform 1 0 71852 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_781
timestamp 1649977179
transform 1 0 72956 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_793
timestamp 1649977179
transform 1 0 74060 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_805
timestamp 1649977179
transform 1 0 75164 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_811
timestamp 1649977179
transform 1 0 75716 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_813
timestamp 1649977179
transform 1 0 75900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_825
timestamp 1649977179
transform 1 0 77004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_830
timestamp 1649977179
transform 1 0 77464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_838
timestamp 1649977179
transform 1 0 78200 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_31
timestamp 1649977179
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_43
timestamp 1649977179
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1649977179
transform 1 0 16928 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_178
timestamp 1649977179
transform 1 0 17480 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_190
timestamp 1649977179
transform 1 0 18584 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_202
timestamp 1649977179
transform 1 0 19688 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_214
timestamp 1649977179
transform 1 0 20792 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1649977179
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_322
timestamp 1649977179
transform 1 0 30728 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1649977179
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_341
timestamp 1649977179
transform 1 0 32476 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_353
timestamp 1649977179
transform 1 0 33580 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_365
timestamp 1649977179
transform 1 0 34684 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_377
timestamp 1649977179
transform 1 0 35788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1649977179
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1649977179
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1649977179
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1649977179
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1649977179
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1649977179
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1649977179
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1649977179
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1649977179
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1649977179
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1649977179
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1649977179
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1649977179
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_729
timestamp 1649977179
transform 1 0 68172 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_741
timestamp 1649977179
transform 1 0 69276 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_753
timestamp 1649977179
transform 1 0 70380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_765
timestamp 1649977179
transform 1 0 71484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_777
timestamp 1649977179
transform 1 0 72588 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_783
timestamp 1649977179
transform 1 0 73140 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_785
timestamp 1649977179
transform 1 0 73324 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_797
timestamp 1649977179
transform 1 0 74428 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_809
timestamp 1649977179
transform 1 0 75532 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_821
timestamp 1649977179
transform 1 0 76636 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_825
timestamp 1649977179
transform 1 0 77004 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_828
timestamp 1649977179
transform 1 0 77280 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_836
timestamp 1649977179
transform 1 0 78016 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_841
timestamp 1649977179
transform 1 0 78476 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1649977179
transform 1 0 17296 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_182
timestamp 1649977179
transform 1 0 17848 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_326
timestamp 1649977179
transform 1 0 31096 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_334
timestamp 1649977179
transform 1 0 31832 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_346
timestamp 1649977179
transform 1 0 32936 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 1649977179
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1649977179
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1649977179
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1649977179
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1649977179
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1649977179
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1649977179
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1649977179
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1649977179
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1649977179
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1649977179
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1649977179
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1649977179
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1649977179
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_725
timestamp 1649977179
transform 1 0 67804 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_737
timestamp 1649977179
transform 1 0 68908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_749
timestamp 1649977179
transform 1 0 70012 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_755
timestamp 1649977179
transform 1 0 70564 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_757
timestamp 1649977179
transform 1 0 70748 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_769
timestamp 1649977179
transform 1 0 71852 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_781
timestamp 1649977179
transform 1 0 72956 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_793
timestamp 1649977179
transform 1 0 74060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_805
timestamp 1649977179
transform 1 0 75164 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_811
timestamp 1649977179
transform 1 0 75716 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_813
timestamp 1649977179
transform 1 0 75900 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_825
timestamp 1649977179
transform 1 0 77004 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_837
timestamp 1649977179
transform 1 0 78108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_841
timestamp 1649977179
transform 1 0 78476 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_7
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_19
timestamp 1649977179
transform 1 0 2852 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_31
timestamp 1649977179
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_43
timestamp 1649977179
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1649977179
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_198
timestamp 1649977179
transform 1 0 19320 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_210
timestamp 1649977179
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1649977179
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1649977179
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_341
timestamp 1649977179
transform 1 0 32476 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_353
timestamp 1649977179
transform 1 0 33580 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_365
timestamp 1649977179
transform 1 0 34684 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_377
timestamp 1649977179
transform 1 0 35788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1649977179
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1649977179
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1649977179
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1649977179
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1649977179
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1649977179
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1649977179
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1649977179
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1649977179
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1649977179
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1649977179
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1649977179
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_729
timestamp 1649977179
transform 1 0 68172 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_741
timestamp 1649977179
transform 1 0 69276 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_753
timestamp 1649977179
transform 1 0 70380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_765
timestamp 1649977179
transform 1 0 71484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_777
timestamp 1649977179
transform 1 0 72588 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_783
timestamp 1649977179
transform 1 0 73140 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_785
timestamp 1649977179
transform 1 0 73324 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_797
timestamp 1649977179
transform 1 0 74428 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_809
timestamp 1649977179
transform 1 0 75532 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_821
timestamp 1649977179
transform 1 0 76636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_825
timestamp 1649977179
transform 1 0 77004 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_828
timestamp 1649977179
transform 1 0 77280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_836
timestamp 1649977179
transform 1 0 78016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_841
timestamp 1649977179
transform 1 0 78476 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_7
timestamp 1649977179
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1649977179
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_181
timestamp 1649977179
transform 1 0 17756 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_185
timestamp 1649977179
transform 1 0 18124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1649977179
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_285
timestamp 1649977179
transform 1 0 27324 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_293
timestamp 1649977179
transform 1 0 28060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1649977179
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1649977179
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1649977179
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1649977179
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1649977179
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1649977179
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1649977179
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1649977179
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1649977179
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1649977179
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1649977179
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1649977179
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_725
timestamp 1649977179
transform 1 0 67804 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_737
timestamp 1649977179
transform 1 0 68908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_749
timestamp 1649977179
transform 1 0 70012 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_755
timestamp 1649977179
transform 1 0 70564 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_757
timestamp 1649977179
transform 1 0 70748 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_769
timestamp 1649977179
transform 1 0 71852 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_781
timestamp 1649977179
transform 1 0 72956 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_793
timestamp 1649977179
transform 1 0 74060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_805
timestamp 1649977179
transform 1 0 75164 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_811
timestamp 1649977179
transform 1 0 75716 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_813
timestamp 1649977179
transform 1 0 75900 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_825
timestamp 1649977179
transform 1 0 77004 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_830
timestamp 1649977179
transform 1 0 77464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_838
timestamp 1649977179
transform 1 0 78200 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_7
timestamp 1649977179
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_19
timestamp 1649977179
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_31
timestamp 1649977179
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_43
timestamp 1649977179
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_198
timestamp 1649977179
transform 1 0 19320 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_204
timestamp 1649977179
transform 1 0 19872 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1649977179
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1649977179
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1649977179
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1649977179
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1649977179
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1649977179
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1649977179
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1649977179
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1649977179
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1649977179
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1649977179
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1649977179
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1649977179
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1649977179
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1649977179
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_729
timestamp 1649977179
transform 1 0 68172 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_741
timestamp 1649977179
transform 1 0 69276 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_753
timestamp 1649977179
transform 1 0 70380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_765
timestamp 1649977179
transform 1 0 71484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_777
timestamp 1649977179
transform 1 0 72588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_783
timestamp 1649977179
transform 1 0 73140 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_785
timestamp 1649977179
transform 1 0 73324 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_797
timestamp 1649977179
transform 1 0 74428 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_809
timestamp 1649977179
transform 1 0 75532 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_821
timestamp 1649977179
transform 1 0 76636 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_825
timestamp 1649977179
transform 1 0 77004 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_828
timestamp 1649977179
transform 1 0 77280 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_836
timestamp 1649977179
transform 1 0 78016 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_841
timestamp 1649977179
transform 1 0 78476 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_7
timestamp 1649977179
transform 1 0 1748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_19
timestamp 1649977179
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_287
timestamp 1649977179
transform 1 0 27508 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_295
timestamp 1649977179
transform 1 0 28244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1649977179
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1649977179
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1649977179
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1649977179
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1649977179
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1649977179
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1649977179
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1649977179
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1649977179
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1649977179
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1649977179
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1649977179
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1649977179
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_725
timestamp 1649977179
transform 1 0 67804 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_737
timestamp 1649977179
transform 1 0 68908 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_749
timestamp 1649977179
transform 1 0 70012 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_755
timestamp 1649977179
transform 1 0 70564 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_757
timestamp 1649977179
transform 1 0 70748 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_769
timestamp 1649977179
transform 1 0 71852 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_781
timestamp 1649977179
transform 1 0 72956 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_793
timestamp 1649977179
transform 1 0 74060 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_805
timestamp 1649977179
transform 1 0 75164 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_811
timestamp 1649977179
transform 1 0 75716 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_813
timestamp 1649977179
transform 1 0 75900 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_825
timestamp 1649977179
transform 1 0 77004 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_830
timestamp 1649977179
transform 1 0 77464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_838
timestamp 1649977179
transform 1 0 78200 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_208
timestamp 1649977179
transform 1 0 20240 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_214
timestamp 1649977179
transform 1 0 20792 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1649977179
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_285
timestamp 1649977179
transform 1 0 27324 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_327
timestamp 1649977179
transform 1 0 31188 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1649977179
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1649977179
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1649977179
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1649977179
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1649977179
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1649977179
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1649977179
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1649977179
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1649977179
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1649977179
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1649977179
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1649977179
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1649977179
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1649977179
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_729
timestamp 1649977179
transform 1 0 68172 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_741
timestamp 1649977179
transform 1 0 69276 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_753
timestamp 1649977179
transform 1 0 70380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_765
timestamp 1649977179
transform 1 0 71484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_777
timestamp 1649977179
transform 1 0 72588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_783
timestamp 1649977179
transform 1 0 73140 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_785
timestamp 1649977179
transform 1 0 73324 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_797
timestamp 1649977179
transform 1 0 74428 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_809
timestamp 1649977179
transform 1 0 75532 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_821
timestamp 1649977179
transform 1 0 76636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_833
timestamp 1649977179
transform 1 0 77740 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_839
timestamp 1649977179
transform 1 0 78292 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_841
timestamp 1649977179
transform 1 0 78476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 1649977179
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_13
timestamp 1649977179
transform 1 0 2300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1649977179
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_201
timestamp 1649977179
transform 1 0 19596 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_205
timestamp 1649977179
transform 1 0 19964 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_211
timestamp 1649977179
transform 1 0 20516 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_223
timestamp 1649977179
transform 1 0 21620 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_235
timestamp 1649977179
transform 1 0 22724 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1649977179
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_277
timestamp 1649977179
transform 1 0 26588 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_285
timestamp 1649977179
transform 1 0 27324 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_293
timestamp 1649977179
transform 1 0 28060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1649977179
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_319
timestamp 1649977179
transform 1 0 30452 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_325
timestamp 1649977179
transform 1 0 31004 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_338
timestamp 1649977179
transform 1 0 32200 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_350
timestamp 1649977179
transform 1 0 33304 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_362
timestamp 1649977179
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1649977179
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1649977179
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1649977179
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1649977179
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1649977179
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1649977179
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1649977179
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1649977179
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1649977179
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1649977179
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1649977179
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1649977179
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_725
timestamp 1649977179
transform 1 0 67804 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_737
timestamp 1649977179
transform 1 0 68908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_749
timestamp 1649977179
transform 1 0 70012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_755
timestamp 1649977179
transform 1 0 70564 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_757
timestamp 1649977179
transform 1 0 70748 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_769
timestamp 1649977179
transform 1 0 71852 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_781
timestamp 1649977179
transform 1 0 72956 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_793
timestamp 1649977179
transform 1 0 74060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_805
timestamp 1649977179
transform 1 0 75164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_811
timestamp 1649977179
transform 1 0 75716 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_813
timestamp 1649977179
transform 1 0 75900 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_825
timestamp 1649977179
transform 1 0 77004 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_830
timestamp 1649977179
transform 1 0 77464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_838
timestamp 1649977179
transform 1 0 78200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_7
timestamp 1649977179
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_13
timestamp 1649977179
transform 1 0 2300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_25
timestamp 1649977179
transform 1 0 3404 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_37
timestamp 1649977179
transform 1 0 4508 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_49
timestamp 1649977179
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_228
timestamp 1649977179
transform 1 0 22080 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_234
timestamp 1649977179
transform 1 0 22632 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_246
timestamp 1649977179
transform 1 0 23736 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_258
timestamp 1649977179
transform 1 0 24840 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_270
timestamp 1649977179
transform 1 0 25944 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1649977179
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_325
timestamp 1649977179
transform 1 0 31004 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1649977179
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_341
timestamp 1649977179
transform 1 0 32476 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_347
timestamp 1649977179
transform 1 0 33028 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_359
timestamp 1649977179
transform 1 0 34132 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_371
timestamp 1649977179
transform 1 0 35236 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_383
timestamp 1649977179
transform 1 0 36340 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1649977179
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_429
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_437
timestamp 1649977179
transform 1 0 41308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_443
timestamp 1649977179
transform 1 0 41860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1649977179
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1649977179
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1649977179
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1649977179
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1649977179
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1649977179
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1649977179
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1649977179
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1649977179
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1649977179
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1649977179
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_729
timestamp 1649977179
transform 1 0 68172 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_741
timestamp 1649977179
transform 1 0 69276 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_753
timestamp 1649977179
transform 1 0 70380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_765
timestamp 1649977179
transform 1 0 71484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_777
timestamp 1649977179
transform 1 0 72588 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_783
timestamp 1649977179
transform 1 0 73140 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_785
timestamp 1649977179
transform 1 0 73324 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_797
timestamp 1649977179
transform 1 0 74428 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_809
timestamp 1649977179
transform 1 0 75532 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_821
timestamp 1649977179
transform 1 0 76636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_825
timestamp 1649977179
transform 1 0 77004 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_828
timestamp 1649977179
transform 1 0 77280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_836
timestamp 1649977179
transform 1 0 78016 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_841
timestamp 1649977179
transform 1 0 78476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_7
timestamp 1649977179
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_13
timestamp 1649977179
transform 1 0 2300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1649977179
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_229
timestamp 1649977179
transform 1 0 22172 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_239
timestamp 1649977179
transform 1 0 23092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_331
timestamp 1649977179
transform 1 0 31556 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_339
timestamp 1649977179
transform 1 0 32292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_351
timestamp 1649977179
transform 1 0 33396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_429
timestamp 1649977179
transform 1 0 40572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_434
timestamp 1649977179
transform 1 0 41032 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_438
timestamp 1649977179
transform 1 0 41400 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1649977179
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1649977179
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1649977179
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1649977179
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1649977179
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1649977179
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1649977179
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1649977179
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1649977179
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1649977179
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1649977179
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_725
timestamp 1649977179
transform 1 0 67804 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_737
timestamp 1649977179
transform 1 0 68908 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_749
timestamp 1649977179
transform 1 0 70012 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_755
timestamp 1649977179
transform 1 0 70564 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_757
timestamp 1649977179
transform 1 0 70748 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_769
timestamp 1649977179
transform 1 0 71852 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_781
timestamp 1649977179
transform 1 0 72956 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_793
timestamp 1649977179
transform 1 0 74060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_805
timestamp 1649977179
transform 1 0 75164 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_811
timestamp 1649977179
transform 1 0 75716 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_813
timestamp 1649977179
transform 1 0 75900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_825
timestamp 1649977179
transform 1 0 77004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_830
timestamp 1649977179
transform 1 0 77464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_838
timestamp 1649977179
transform 1 0 78200 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_7
timestamp 1649977179
transform 1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_13
timestamp 1649977179
transform 1 0 2300 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_25
timestamp 1649977179
transform 1 0 3404 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_37
timestamp 1649977179
transform 1 0 4508 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_49
timestamp 1649977179
transform 1 0 5612 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_432
timestamp 1649977179
transform 1 0 40848 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_444
timestamp 1649977179
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1649977179
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1649977179
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1649977179
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1649977179
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1649977179
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1649977179
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1649977179
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1649977179
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1649977179
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1649977179
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1649977179
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_729
timestamp 1649977179
transform 1 0 68172 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_741
timestamp 1649977179
transform 1 0 69276 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_753
timestamp 1649977179
transform 1 0 70380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_765
timestamp 1649977179
transform 1 0 71484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_777
timestamp 1649977179
transform 1 0 72588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_783
timestamp 1649977179
transform 1 0 73140 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_785
timestamp 1649977179
transform 1 0 73324 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_797
timestamp 1649977179
transform 1 0 74428 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_809
timestamp 1649977179
transform 1 0 75532 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_821
timestamp 1649977179
transform 1 0 76636 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_825
timestamp 1649977179
transform 1 0 77004 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_828
timestamp 1649977179
transform 1 0 77280 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_836
timestamp 1649977179
transform 1 0 78016 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_841
timestamp 1649977179
transform 1 0 78476 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_229
timestamp 1649977179
transform 1 0 22172 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_239
timestamp 1649977179
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_337
timestamp 1649977179
transform 1 0 32108 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1649977179
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1649977179
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1649977179
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_645
timestamp 1649977179
transform 1 0 60444 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_657
timestamp 1649977179
transform 1 0 61548 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_669
timestamp 1649977179
transform 1 0 62652 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_681
timestamp 1649977179
transform 1 0 63756 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_693
timestamp 1649977179
transform 1 0 64860 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1649977179
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1649977179
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1649977179
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_725
timestamp 1649977179
transform 1 0 67804 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_737
timestamp 1649977179
transform 1 0 68908 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_749
timestamp 1649977179
transform 1 0 70012 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_755
timestamp 1649977179
transform 1 0 70564 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_757
timestamp 1649977179
transform 1 0 70748 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_769
timestamp 1649977179
transform 1 0 71852 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_781
timestamp 1649977179
transform 1 0 72956 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_793
timestamp 1649977179
transform 1 0 74060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_805
timestamp 1649977179
transform 1 0 75164 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_811
timestamp 1649977179
transform 1 0 75716 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_813
timestamp 1649977179
transform 1 0 75900 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_825
timestamp 1649977179
transform 1 0 77004 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_837
timestamp 1649977179
transform 1 0 78108 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_841
timestamp 1649977179
transform 1 0 78476 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_7
timestamp 1649977179
transform 1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_13
timestamp 1649977179
transform 1 0 2300 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_25
timestamp 1649977179
transform 1 0 3404 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_37
timestamp 1649977179
transform 1 0 4508 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_49
timestamp 1649977179
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_233
timestamp 1649977179
transform 1 0 22540 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_240
timestamp 1649977179
transform 1 0 23184 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_246
timestamp 1649977179
transform 1 0 23736 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_258
timestamp 1649977179
transform 1 0 24840 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_264
timestamp 1649977179
transform 1 0 25392 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_267
timestamp 1649977179
transform 1 0 25668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_341
timestamp 1649977179
transform 1 0 32476 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_346
timestamp 1649977179
transform 1 0 32936 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_358
timestamp 1649977179
transform 1 0 34040 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_370
timestamp 1649977179
transform 1 0 35144 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 1649977179
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1649977179
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1649977179
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1649977179
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1649977179
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1649977179
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1649977179
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1649977179
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1649977179
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1649977179
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1649977179
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1649977179
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1649977179
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1649977179
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_729
timestamp 1649977179
transform 1 0 68172 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_741
timestamp 1649977179
transform 1 0 69276 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_753
timestamp 1649977179
transform 1 0 70380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_765
timestamp 1649977179
transform 1 0 71484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_777
timestamp 1649977179
transform 1 0 72588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_783
timestamp 1649977179
transform 1 0 73140 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_785
timestamp 1649977179
transform 1 0 73324 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_797
timestamp 1649977179
transform 1 0 74428 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_809
timestamp 1649977179
transform 1 0 75532 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_821
timestamp 1649977179
transform 1 0 76636 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_825
timestamp 1649977179
transform 1 0 77004 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_828
timestamp 1649977179
transform 1 0 77280 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_836
timestamp 1649977179
transform 1 0 78016 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_841
timestamp 1649977179
transform 1 0 78476 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_7
timestamp 1649977179
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_13
timestamp 1649977179
transform 1 0 2300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_25
timestamp 1649977179
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_273
timestamp 1649977179
transform 1 0 26220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_281
timestamp 1649977179
transform 1 0 26956 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_287
timestamp 1649977179
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1649977179
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_339
timestamp 1649977179
transform 1 0 32292 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_342
timestamp 1649977179
transform 1 0 32568 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_354
timestamp 1649977179
transform 1 0 33672 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_362
timestamp 1649977179
transform 1 0 34408 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1649977179
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1649977179
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1649977179
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1649977179
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1649977179
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1649977179
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1649977179
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1649977179
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1649977179
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1649977179
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1649977179
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1649977179
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1649977179
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_725
timestamp 1649977179
transform 1 0 67804 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_737
timestamp 1649977179
transform 1 0 68908 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_749
timestamp 1649977179
transform 1 0 70012 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_755
timestamp 1649977179
transform 1 0 70564 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_757
timestamp 1649977179
transform 1 0 70748 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_769
timestamp 1649977179
transform 1 0 71852 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_781
timestamp 1649977179
transform 1 0 72956 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_793
timestamp 1649977179
transform 1 0 74060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_805
timestamp 1649977179
transform 1 0 75164 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_811
timestamp 1649977179
transform 1 0 75716 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_813
timestamp 1649977179
transform 1 0 75900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_825
timestamp 1649977179
transform 1 0 77004 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_830
timestamp 1649977179
transform 1 0 77464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_838
timestamp 1649977179
transform 1 0 78200 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_7
timestamp 1649977179
transform 1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_13
timestamp 1649977179
transform 1 0 2300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_25
timestamp 1649977179
transform 1 0 3404 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_37
timestamp 1649977179
transform 1 0 4508 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1649977179
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_269
timestamp 1649977179
transform 1 0 25852 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1649977179
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_289
timestamp 1649977179
transform 1 0 27692 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_301
timestamp 1649977179
transform 1 0 28796 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_313
timestamp 1649977179
transform 1 0 29900 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_325
timestamp 1649977179
transform 1 0 31004 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_333
timestamp 1649977179
transform 1 0 31740 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1649977179
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1649977179
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1649977179
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1649977179
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1649977179
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1649977179
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1649977179
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1649977179
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1649977179
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1649977179
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1649977179
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_729
timestamp 1649977179
transform 1 0 68172 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_741
timestamp 1649977179
transform 1 0 69276 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_753
timestamp 1649977179
transform 1 0 70380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_765
timestamp 1649977179
transform 1 0 71484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_777
timestamp 1649977179
transform 1 0 72588 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_783
timestamp 1649977179
transform 1 0 73140 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_785
timestamp 1649977179
transform 1 0 73324 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_797
timestamp 1649977179
transform 1 0 74428 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_809
timestamp 1649977179
transform 1 0 75532 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_821
timestamp 1649977179
transform 1 0 76636 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_825
timestamp 1649977179
transform 1 0 77004 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_828
timestamp 1649977179
transform 1 0 77280 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_836
timestamp 1649977179
transform 1 0 78016 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_841
timestamp 1649977179
transform 1 0 78476 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_7
timestamp 1649977179
transform 1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_13
timestamp 1649977179
transform 1 0 2300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_25
timestamp 1649977179
transform 1 0 3404 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_273
timestamp 1649977179
transform 1 0 26220 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_276
timestamp 1649977179
transform 1 0 26496 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_284
timestamp 1649977179
transform 1 0 27232 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_287
timestamp 1649977179
transform 1 0 27508 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_293
timestamp 1649977179
transform 1 0 28060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_305
timestamp 1649977179
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1649977179
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1649977179
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1649977179
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1649977179
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1649977179
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1649977179
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1649977179
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1649977179
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1649977179
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1649977179
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1649977179
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1649977179
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1649977179
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_725
timestamp 1649977179
transform 1 0 67804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_737
timestamp 1649977179
transform 1 0 68908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_749
timestamp 1649977179
transform 1 0 70012 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_755
timestamp 1649977179
transform 1 0 70564 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_757
timestamp 1649977179
transform 1 0 70748 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_769
timestamp 1649977179
transform 1 0 71852 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_781
timestamp 1649977179
transform 1 0 72956 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_793
timestamp 1649977179
transform 1 0 74060 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_805
timestamp 1649977179
transform 1 0 75164 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_811
timestamp 1649977179
transform 1 0 75716 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_813
timestamp 1649977179
transform 1 0 75900 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_825
timestamp 1649977179
transform 1 0 77004 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_830
timestamp 1649977179
transform 1 0 77464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_838
timestamp 1649977179
transform 1 0 78200 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1649977179
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1649977179
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_285
timestamp 1649977179
transform 1 0 27324 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_297
timestamp 1649977179
transform 1 0 28428 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_309
timestamp 1649977179
transform 1 0 29532 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_321
timestamp 1649977179
transform 1 0 30636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_333
timestamp 1649977179
transform 1 0 31740 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1649977179
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1649977179
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1649977179
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1649977179
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1649977179
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1649977179
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1649977179
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1649977179
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1649977179
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1649977179
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1649977179
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_729
timestamp 1649977179
transform 1 0 68172 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_741
timestamp 1649977179
transform 1 0 69276 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_753
timestamp 1649977179
transform 1 0 70380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_765
timestamp 1649977179
transform 1 0 71484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_777
timestamp 1649977179
transform 1 0 72588 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_783
timestamp 1649977179
transform 1 0 73140 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_785
timestamp 1649977179
transform 1 0 73324 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_797
timestamp 1649977179
transform 1 0 74428 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_809
timestamp 1649977179
transform 1 0 75532 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_821
timestamp 1649977179
transform 1 0 76636 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_833
timestamp 1649977179
transform 1 0 77740 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_839
timestamp 1649977179
transform 1 0 78292 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_841
timestamp 1649977179
transform 1 0 78476 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_7
timestamp 1649977179
transform 1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_13
timestamp 1649977179
transform 1 0 2300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_25
timestamp 1649977179
transform 1 0 3404 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_282
timestamp 1649977179
transform 1 0 27048 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_290
timestamp 1649977179
transform 1 0 27784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_296
timestamp 1649977179
transform 1 0 28336 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1649977179
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1649977179
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1649977179
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1649977179
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1649977179
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1649977179
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1649977179
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1649977179
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1649977179
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1649977179
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1649977179
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1649977179
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_725
timestamp 1649977179
transform 1 0 67804 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_737
timestamp 1649977179
transform 1 0 68908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_749
timestamp 1649977179
transform 1 0 70012 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_755
timestamp 1649977179
transform 1 0 70564 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_757
timestamp 1649977179
transform 1 0 70748 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_769
timestamp 1649977179
transform 1 0 71852 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_781
timestamp 1649977179
transform 1 0 72956 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_793
timestamp 1649977179
transform 1 0 74060 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_805
timestamp 1649977179
transform 1 0 75164 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_811
timestamp 1649977179
transform 1 0 75716 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_813
timestamp 1649977179
transform 1 0 75900 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_825
timestamp 1649977179
transform 1 0 77004 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_830
timestamp 1649977179
transform 1 0 77464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_838
timestamp 1649977179
transform 1 0 78200 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_7
timestamp 1649977179
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_13
timestamp 1649977179
transform 1 0 2300 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_25
timestamp 1649977179
transform 1 0 3404 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_37
timestamp 1649977179
transform 1 0 4508 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_49
timestamp 1649977179
transform 1 0 5612 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_287
timestamp 1649977179
transform 1 0 27508 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_290
timestamp 1649977179
transform 1 0 27784 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_298
timestamp 1649977179
transform 1 0 28520 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_304
timestamp 1649977179
transform 1 0 29072 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_312
timestamp 1649977179
transform 1 0 29808 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_324
timestamp 1649977179
transform 1 0 30912 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1649977179
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1649977179
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1649977179
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1649977179
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1649977179
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1649977179
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1649977179
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1649977179
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1649977179
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1649977179
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1649977179
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1649977179
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1649977179
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_729
timestamp 1649977179
transform 1 0 68172 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_741
timestamp 1649977179
transform 1 0 69276 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_753
timestamp 1649977179
transform 1 0 70380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_765
timestamp 1649977179
transform 1 0 71484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_777
timestamp 1649977179
transform 1 0 72588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_783
timestamp 1649977179
transform 1 0 73140 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_785
timestamp 1649977179
transform 1 0 73324 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_797
timestamp 1649977179
transform 1 0 74428 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_809
timestamp 1649977179
transform 1 0 75532 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_821
timestamp 1649977179
transform 1 0 76636 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_825
timestamp 1649977179
transform 1 0 77004 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_828
timestamp 1649977179
transform 1 0 77280 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_836
timestamp 1649977179
transform 1 0 78016 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_841
timestamp 1649977179
transform 1 0 78476 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_7
timestamp 1649977179
transform 1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_13
timestamp 1649977179
transform 1 0 2300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_25
timestamp 1649977179
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_297
timestamp 1649977179
transform 1 0 28428 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1649977179
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_311
timestamp 1649977179
transform 1 0 29716 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_319
timestamp 1649977179
transform 1 0 30452 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_331
timestamp 1649977179
transform 1 0 31556 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_343
timestamp 1649977179
transform 1 0 32660 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_355
timestamp 1649977179
transform 1 0 33764 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1649977179
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1649977179
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1649977179
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1649977179
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1649977179
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1649977179
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1649977179
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1649977179
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1649977179
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1649977179
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1649977179
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1649977179
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_713
timestamp 1649977179
transform 1 0 66700 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_725
timestamp 1649977179
transform 1 0 67804 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_737
timestamp 1649977179
transform 1 0 68908 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_749
timestamp 1649977179
transform 1 0 70012 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_755
timestamp 1649977179
transform 1 0 70564 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_757
timestamp 1649977179
transform 1 0 70748 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_769
timestamp 1649977179
transform 1 0 71852 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_781
timestamp 1649977179
transform 1 0 72956 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_793
timestamp 1649977179
transform 1 0 74060 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_805
timestamp 1649977179
transform 1 0 75164 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_811
timestamp 1649977179
transform 1 0 75716 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_813
timestamp 1649977179
transform 1 0 75900 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_825
timestamp 1649977179
transform 1 0 77004 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_830
timestamp 1649977179
transform 1 0 77464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_838
timestamp 1649977179
transform 1 0 78200 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_7
timestamp 1649977179
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_13
timestamp 1649977179
transform 1 0 2300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_25
timestamp 1649977179
transform 1 0 3404 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_37
timestamp 1649977179
transform 1 0 4508 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 1649977179
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_301
timestamp 1649977179
transform 1 0 28796 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_306
timestamp 1649977179
transform 1 0 29256 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_316
timestamp 1649977179
transform 1 0 30176 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_320
timestamp 1649977179
transform 1 0 30544 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_323
timestamp 1649977179
transform 1 0 30820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1649977179
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1649977179
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1649977179
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1649977179
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1649977179
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1649977179
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1649977179
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1649977179
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1649977179
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1649977179
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1649977179
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1649977179
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_729
timestamp 1649977179
transform 1 0 68172 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_741
timestamp 1649977179
transform 1 0 69276 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_753
timestamp 1649977179
transform 1 0 70380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_765
timestamp 1649977179
transform 1 0 71484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_777
timestamp 1649977179
transform 1 0 72588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_783
timestamp 1649977179
transform 1 0 73140 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_785
timestamp 1649977179
transform 1 0 73324 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_797
timestamp 1649977179
transform 1 0 74428 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_809
timestamp 1649977179
transform 1 0 75532 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_821
timestamp 1649977179
transform 1 0 76636 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_825
timestamp 1649977179
transform 1 0 77004 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_828
timestamp 1649977179
transform 1 0 77280 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_836
timestamp 1649977179
transform 1 0 78016 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_841
timestamp 1649977179
transform 1 0 78476 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_314
timestamp 1649977179
transform 1 0 29992 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_322
timestamp 1649977179
transform 1 0 30728 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_327
timestamp 1649977179
transform 1 0 31188 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_337
timestamp 1649977179
transform 1 0 32108 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_349
timestamp 1649977179
transform 1 0 33212 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1649977179
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1649977179
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1649977179
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1649977179
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1649977179
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1649977179
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1649977179
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1649977179
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1649977179
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1649977179
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1649977179
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1649977179
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1649977179
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_725
timestamp 1649977179
transform 1 0 67804 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_737
timestamp 1649977179
transform 1 0 68908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_749
timestamp 1649977179
transform 1 0 70012 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_755
timestamp 1649977179
transform 1 0 70564 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_757
timestamp 1649977179
transform 1 0 70748 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_769
timestamp 1649977179
transform 1 0 71852 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_781
timestamp 1649977179
transform 1 0 72956 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_793
timestamp 1649977179
transform 1 0 74060 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_805
timestamp 1649977179
transform 1 0 75164 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_811
timestamp 1649977179
transform 1 0 75716 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_813
timestamp 1649977179
transform 1 0 75900 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_825
timestamp 1649977179
transform 1 0 77004 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_837
timestamp 1649977179
transform 1 0 78108 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_841
timestamp 1649977179
transform 1 0 78476 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_7
timestamp 1649977179
transform 1 0 1748 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_13
timestamp 1649977179
transform 1 0 2300 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_25
timestamp 1649977179
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_37
timestamp 1649977179
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_49
timestamp 1649977179
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_311
timestamp 1649977179
transform 1 0 29716 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_314
timestamp 1649977179
transform 1 0 29992 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_322
timestamp 1649977179
transform 1 0 30728 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1649977179
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_341
timestamp 1649977179
transform 1 0 32476 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_347
timestamp 1649977179
transform 1 0 33028 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_359
timestamp 1649977179
transform 1 0 34132 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_371
timestamp 1649977179
transform 1 0 35236 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_383
timestamp 1649977179
transform 1 0 36340 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1649977179
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1649977179
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1649977179
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1649977179
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1649977179
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1649977179
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1649977179
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1649977179
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1649977179
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1649977179
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1649977179
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_729
timestamp 1649977179
transform 1 0 68172 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_741
timestamp 1649977179
transform 1 0 69276 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_753
timestamp 1649977179
transform 1 0 70380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_765
timestamp 1649977179
transform 1 0 71484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_777
timestamp 1649977179
transform 1 0 72588 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_783
timestamp 1649977179
transform 1 0 73140 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_785
timestamp 1649977179
transform 1 0 73324 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_797
timestamp 1649977179
transform 1 0 74428 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_809
timestamp 1649977179
transform 1 0 75532 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_821
timestamp 1649977179
transform 1 0 76636 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_825
timestamp 1649977179
transform 1 0 77004 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_828
timestamp 1649977179
transform 1 0 77280 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_836
timestamp 1649977179
transform 1 0 78016 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_841
timestamp 1649977179
transform 1 0 78476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_7
timestamp 1649977179
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_13
timestamp 1649977179
transform 1 0 2300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_25
timestamp 1649977179
transform 1 0 3404 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_325
timestamp 1649977179
transform 1 0 31004 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_330
timestamp 1649977179
transform 1 0 31464 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_342
timestamp 1649977179
transform 1 0 32568 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_348
timestamp 1649977179
transform 1 0 33120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1649977179
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1649977179
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_625
timestamp 1649977179
transform 1 0 58604 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_637
timestamp 1649977179
transform 1 0 59708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_643
timestamp 1649977179
transform 1 0 60260 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1649977179
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1649977179
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1649977179
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1649977179
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1649977179
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1649977179
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1649977179
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1649977179
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_725
timestamp 1649977179
transform 1 0 67804 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_737
timestamp 1649977179
transform 1 0 68908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_749
timestamp 1649977179
transform 1 0 70012 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_755
timestamp 1649977179
transform 1 0 70564 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_757
timestamp 1649977179
transform 1 0 70748 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_769
timestamp 1649977179
transform 1 0 71852 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_781
timestamp 1649977179
transform 1 0 72956 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_793
timestamp 1649977179
transform 1 0 74060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_805
timestamp 1649977179
transform 1 0 75164 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_811
timestamp 1649977179
transform 1 0 75716 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_813
timestamp 1649977179
transform 1 0 75900 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_825
timestamp 1649977179
transform 1 0 77004 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_830
timestamp 1649977179
transform 1 0 77464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_838
timestamp 1649977179
transform 1 0 78200 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_7
timestamp 1649977179
transform 1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_13
timestamp 1649977179
transform 1 0 2300 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_25
timestamp 1649977179
transform 1 0 3404 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_37
timestamp 1649977179
transform 1 0 4508 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_49
timestamp 1649977179
transform 1 0 5612 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_341
timestamp 1649977179
transform 1 0 32476 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1649977179
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1649977179
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1649977179
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1649977179
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1649977179
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1649977179
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1649977179
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1649977179
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1649977179
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 1649977179
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 1649977179
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_729
timestamp 1649977179
transform 1 0 68172 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_741
timestamp 1649977179
transform 1 0 69276 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_753
timestamp 1649977179
transform 1 0 70380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_765
timestamp 1649977179
transform 1 0 71484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_777
timestamp 1649977179
transform 1 0 72588 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_783
timestamp 1649977179
transform 1 0 73140 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_785
timestamp 1649977179
transform 1 0 73324 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_797
timestamp 1649977179
transform 1 0 74428 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_809
timestamp 1649977179
transform 1 0 75532 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_821
timestamp 1649977179
transform 1 0 76636 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_825
timestamp 1649977179
transform 1 0 77004 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_828
timestamp 1649977179
transform 1 0 77280 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_836
timestamp 1649977179
transform 1 0 78016 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_841
timestamp 1649977179
transform 1 0 78476 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_7
timestamp 1649977179
transform 1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_13
timestamp 1649977179
transform 1 0 2300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_25
timestamp 1649977179
transform 1 0 3404 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_341
timestamp 1649977179
transform 1 0 32476 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_353
timestamp 1649977179
transform 1 0 33580 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_361
timestamp 1649977179
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1649977179
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1649977179
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1649977179
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1649977179
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1649977179
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1649977179
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1649977179
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1649977179
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1649977179
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1649977179
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1649977179
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_725
timestamp 1649977179
transform 1 0 67804 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_737
timestamp 1649977179
transform 1 0 68908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_749
timestamp 1649977179
transform 1 0 70012 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_755
timestamp 1649977179
transform 1 0 70564 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_757
timestamp 1649977179
transform 1 0 70748 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_769
timestamp 1649977179
transform 1 0 71852 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_781
timestamp 1649977179
transform 1 0 72956 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_793
timestamp 1649977179
transform 1 0 74060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_805
timestamp 1649977179
transform 1 0 75164 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_811
timestamp 1649977179
transform 1 0 75716 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_813
timestamp 1649977179
transform 1 0 75900 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_825
timestamp 1649977179
transform 1 0 77004 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_830
timestamp 1649977179
transform 1 0 77464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_838
timestamp 1649977179
transform 1 0 78200 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_341
timestamp 1649977179
transform 1 0 32476 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_346
timestamp 1649977179
transform 1 0 32936 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_352
timestamp 1649977179
transform 1 0 33488 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_357
timestamp 1649977179
transform 1 0 33948 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_363
timestamp 1649977179
transform 1 0 34500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_375
timestamp 1649977179
transform 1 0 35604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_387
timestamp 1649977179
transform 1 0 36708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1649977179
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1649977179
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1649977179
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1649977179
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1649977179
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1649977179
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1649977179
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1649977179
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1649977179
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1649977179
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1649977179
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_729
timestamp 1649977179
transform 1 0 68172 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_741
timestamp 1649977179
transform 1 0 69276 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_753
timestamp 1649977179
transform 1 0 70380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_765
timestamp 1649977179
transform 1 0 71484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_777
timestamp 1649977179
transform 1 0 72588 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_783
timestamp 1649977179
transform 1 0 73140 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_785
timestamp 1649977179
transform 1 0 73324 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_797
timestamp 1649977179
transform 1 0 74428 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_809
timestamp 1649977179
transform 1 0 75532 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_821
timestamp 1649977179
transform 1 0 76636 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_833
timestamp 1649977179
transform 1 0 77740 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_839
timestamp 1649977179
transform 1 0 78292 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_841
timestamp 1649977179
transform 1 0 78476 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_7
timestamp 1649977179
transform 1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_13
timestamp 1649977179
transform 1 0 2300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_25
timestamp 1649977179
transform 1 0 3404 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_341
timestamp 1649977179
transform 1 0 32476 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_346
timestamp 1649977179
transform 1 0 32936 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_354
timestamp 1649977179
transform 1 0 33672 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1649977179
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_369
timestamp 1649977179
transform 1 0 35052 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_375
timestamp 1649977179
transform 1 0 35604 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_387
timestamp 1649977179
transform 1 0 36708 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_399
timestamp 1649977179
transform 1 0 37812 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_411
timestamp 1649977179
transform 1 0 38916 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1649977179
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1649977179
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1649977179
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1649977179
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1649977179
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1649977179
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1649977179
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1649977179
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1649977179
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1649977179
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1649977179
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_725
timestamp 1649977179
transform 1 0 67804 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_737
timestamp 1649977179
transform 1 0 68908 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_749
timestamp 1649977179
transform 1 0 70012 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_755
timestamp 1649977179
transform 1 0 70564 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_757
timestamp 1649977179
transform 1 0 70748 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_769
timestamp 1649977179
transform 1 0 71852 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_781
timestamp 1649977179
transform 1 0 72956 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_793
timestamp 1649977179
transform 1 0 74060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_805
timestamp 1649977179
transform 1 0 75164 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_811
timestamp 1649977179
transform 1 0 75716 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_813
timestamp 1649977179
transform 1 0 75900 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_825
timestamp 1649977179
transform 1 0 77004 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_830
timestamp 1649977179
transform 1 0 77464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_838
timestamp 1649977179
transform 1 0 78200 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_7
timestamp 1649977179
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_13
timestamp 1649977179
transform 1 0 2300 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_25
timestamp 1649977179
transform 1 0 3404 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_37
timestamp 1649977179
transform 1 0 4508 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_49
timestamp 1649977179
transform 1 0 5612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_354
timestamp 1649977179
transform 1 0 33672 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_362
timestamp 1649977179
transform 1 0 34408 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_372
timestamp 1649977179
transform 1 0 35328 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_378
timestamp 1649977179
transform 1 0 35880 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1649977179
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1649977179
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1649977179
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1649977179
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1649977179
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1649977179
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1649977179
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1649977179
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1649977179
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1649977179
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1649977179
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1649977179
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_729
timestamp 1649977179
transform 1 0 68172 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_741
timestamp 1649977179
transform 1 0 69276 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_753
timestamp 1649977179
transform 1 0 70380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_765
timestamp 1649977179
transform 1 0 71484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_777
timestamp 1649977179
transform 1 0 72588 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_783
timestamp 1649977179
transform 1 0 73140 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_785
timestamp 1649977179
transform 1 0 73324 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_797
timestamp 1649977179
transform 1 0 74428 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_809
timestamp 1649977179
transform 1 0 75532 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_821
timestamp 1649977179
transform 1 0 76636 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_825
timestamp 1649977179
transform 1 0 77004 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_828
timestamp 1649977179
transform 1 0 77280 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_836
timestamp 1649977179
transform 1 0 78016 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_841
timestamp 1649977179
transform 1 0 78476 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_7
timestamp 1649977179
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_13
timestamp 1649977179
transform 1 0 2300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_25
timestamp 1649977179
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_370
timestamp 1649977179
transform 1 0 35144 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_380
timestamp 1649977179
transform 1 0 36064 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_392
timestamp 1649977179
transform 1 0 37168 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_404
timestamp 1649977179
transform 1 0 38272 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_416
timestamp 1649977179
transform 1 0 39376 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1649977179
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1649977179
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1649977179
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1649977179
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1649977179
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_669
timestamp 1649977179
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_681
timestamp 1649977179
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1649977179
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1649977179
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1649977179
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1649977179
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_725
timestamp 1649977179
transform 1 0 67804 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_737
timestamp 1649977179
transform 1 0 68908 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_749
timestamp 1649977179
transform 1 0 70012 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_755
timestamp 1649977179
transform 1 0 70564 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_757
timestamp 1649977179
transform 1 0 70748 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_769
timestamp 1649977179
transform 1 0 71852 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_781
timestamp 1649977179
transform 1 0 72956 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_793
timestamp 1649977179
transform 1 0 74060 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_805
timestamp 1649977179
transform 1 0 75164 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_811
timestamp 1649977179
transform 1 0 75716 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_813
timestamp 1649977179
transform 1 0 75900 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_825
timestamp 1649977179
transform 1 0 77004 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_830
timestamp 1649977179
transform 1 0 77464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_838
timestamp 1649977179
transform 1 0 78200 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1649977179
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_13
timestamp 1649977179
transform 1 0 2300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_25
timestamp 1649977179
transform 1 0 3404 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_37
timestamp 1649977179
transform 1 0 4508 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_49
timestamp 1649977179
transform 1 0 5612 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_376
timestamp 1649977179
transform 1 0 35696 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_384
timestamp 1649977179
transform 1 0 36432 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_629
timestamp 1649977179
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_641
timestamp 1649977179
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_653
timestamp 1649977179
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1649977179
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1649977179
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_673
timestamp 1649977179
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_685
timestamp 1649977179
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_697
timestamp 1649977179
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_709
timestamp 1649977179
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1649977179
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1649977179
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_729
timestamp 1649977179
transform 1 0 68172 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_741
timestamp 1649977179
transform 1 0 69276 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_753
timestamp 1649977179
transform 1 0 70380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_765
timestamp 1649977179
transform 1 0 71484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_777
timestamp 1649977179
transform 1 0 72588 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_783
timestamp 1649977179
transform 1 0 73140 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_785
timestamp 1649977179
transform 1 0 73324 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_797
timestamp 1649977179
transform 1 0 74428 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_809
timestamp 1649977179
transform 1 0 75532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_821
timestamp 1649977179
transform 1 0 76636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_825
timestamp 1649977179
transform 1 0 77004 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_828
timestamp 1649977179
transform 1 0 77280 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_836
timestamp 1649977179
transform 1 0 78016 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_841
timestamp 1649977179
transform 1 0 78476 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_370
timestamp 1649977179
transform 1 0 35144 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_378
timestamp 1649977179
transform 1 0 35880 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_388
timestamp 1649977179
transform 1 0 36800 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_394
timestamp 1649977179
transform 1 0 37352 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_406
timestamp 1649977179
transform 1 0 38456 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_418
timestamp 1649977179
transform 1 0 39560 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_625
timestamp 1649977179
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1649977179
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1649977179
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1649977179
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1649977179
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1649977179
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1649977179
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1649977179
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1649977179
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_701
timestamp 1649977179
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_713
timestamp 1649977179
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_725
timestamp 1649977179
transform 1 0 67804 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_737
timestamp 1649977179
transform 1 0 68908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_749
timestamp 1649977179
transform 1 0 70012 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_755
timestamp 1649977179
transform 1 0 70564 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_757
timestamp 1649977179
transform 1 0 70748 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_769
timestamp 1649977179
transform 1 0 71852 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_781
timestamp 1649977179
transform 1 0 72956 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_793
timestamp 1649977179
transform 1 0 74060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_805
timestamp 1649977179
transform 1 0 75164 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_811
timestamp 1649977179
transform 1 0 75716 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_813
timestamp 1649977179
transform 1 0 75900 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_825
timestamp 1649977179
transform 1 0 77004 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_837
timestamp 1649977179
transform 1 0 78108 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_841
timestamp 1649977179
transform 1 0 78476 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_7
timestamp 1649977179
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_13
timestamp 1649977179
transform 1 0 2300 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_25
timestamp 1649977179
transform 1 0 3404 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_37
timestamp 1649977179
transform 1 0 4508 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_49
timestamp 1649977179
transform 1 0 5612 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_377
timestamp 1649977179
transform 1 0 35788 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_397
timestamp 1649977179
transform 1 0 37628 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_403
timestamp 1649977179
transform 1 0 38180 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_415
timestamp 1649977179
transform 1 0 39284 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_427
timestamp 1649977179
transform 1 0 40388 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_439
timestamp 1649977179
transform 1 0 41492 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_629
timestamp 1649977179
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_641
timestamp 1649977179
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_653
timestamp 1649977179
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1649977179
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1649977179
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1649977179
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_685
timestamp 1649977179
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_697
timestamp 1649977179
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_709
timestamp 1649977179
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1649977179
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1649977179
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_729
timestamp 1649977179
transform 1 0 68172 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_741
timestamp 1649977179
transform 1 0 69276 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_753
timestamp 1649977179
transform 1 0 70380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_765
timestamp 1649977179
transform 1 0 71484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_777
timestamp 1649977179
transform 1 0 72588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_783
timestamp 1649977179
transform 1 0 73140 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_785
timestamp 1649977179
transform 1 0 73324 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_797
timestamp 1649977179
transform 1 0 74428 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_809
timestamp 1649977179
transform 1 0 75532 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_821
timestamp 1649977179
transform 1 0 76636 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_825
timestamp 1649977179
transform 1 0 77004 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_828
timestamp 1649977179
transform 1 0 77280 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_836
timestamp 1649977179
transform 1 0 78016 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_841
timestamp 1649977179
transform 1 0 78476 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_7
timestamp 1649977179
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_13
timestamp 1649977179
transform 1 0 2300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1649977179
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1649977179
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_385
timestamp 1649977179
transform 1 0 36524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_393
timestamp 1649977179
transform 1 0 37260 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1649977179
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_409
timestamp 1649977179
transform 1 0 38732 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1649977179
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_625
timestamp 1649977179
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1649977179
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1649977179
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1649977179
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1649977179
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_669
timestamp 1649977179
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_681
timestamp 1649977179
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_693
timestamp 1649977179
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1649977179
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_701
timestamp 1649977179
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_713
timestamp 1649977179
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_725
timestamp 1649977179
transform 1 0 67804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_737
timestamp 1649977179
transform 1 0 68908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_749
timestamp 1649977179
transform 1 0 70012 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_755
timestamp 1649977179
transform 1 0 70564 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_757
timestamp 1649977179
transform 1 0 70748 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_769
timestamp 1649977179
transform 1 0 71852 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_781
timestamp 1649977179
transform 1 0 72956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_793
timestamp 1649977179
transform 1 0 74060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_805
timestamp 1649977179
transform 1 0 75164 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_811
timestamp 1649977179
transform 1 0 75716 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_813
timestamp 1649977179
transform 1 0 75900 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_825
timestamp 1649977179
transform 1 0 77004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_830
timestamp 1649977179
transform 1 0 77464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_838
timestamp 1649977179
transform 1 0 78200 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_7
timestamp 1649977179
transform 1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_13
timestamp 1649977179
transform 1 0 2300 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_25
timestamp 1649977179
transform 1 0 3404 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_37
timestamp 1649977179
transform 1 0 4508 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_49
timestamp 1649977179
transform 1 0 5612 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1649977179
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1649977179
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_401
timestamp 1649977179
transform 1 0 37996 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_411
timestamp 1649977179
transform 1 0 38916 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_423
timestamp 1649977179
transform 1 0 40020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_435
timestamp 1649977179
transform 1 0 41124 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_629
timestamp 1649977179
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_641
timestamp 1649977179
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_653
timestamp 1649977179
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1649977179
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1649977179
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_673
timestamp 1649977179
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_685
timestamp 1649977179
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_697
timestamp 1649977179
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_709
timestamp 1649977179
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_721
timestamp 1649977179
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_727
timestamp 1649977179
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_729
timestamp 1649977179
transform 1 0 68172 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_741
timestamp 1649977179
transform 1 0 69276 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_753
timestamp 1649977179
transform 1 0 70380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_765
timestamp 1649977179
transform 1 0 71484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_777
timestamp 1649977179
transform 1 0 72588 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_783
timestamp 1649977179
transform 1 0 73140 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_785
timestamp 1649977179
transform 1 0 73324 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_797
timestamp 1649977179
transform 1 0 74428 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_809
timestamp 1649977179
transform 1 0 75532 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_821
timestamp 1649977179
transform 1 0 76636 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_825
timestamp 1649977179
transform 1 0 77004 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_828
timestamp 1649977179
transform 1 0 77280 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_836
timestamp 1649977179
transform 1 0 78016 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_841
timestamp 1649977179
transform 1 0 78476 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_7
timestamp 1649977179
transform 1 0 1748 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_13
timestamp 1649977179
transform 1 0 2300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_25
timestamp 1649977179
transform 1 0 3404 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1649977179
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_407
timestamp 1649977179
transform 1 0 38548 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_415
timestamp 1649977179
transform 1 0 39284 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_625
timestamp 1649977179
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1649977179
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1649977179
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_645
timestamp 1649977179
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_657
timestamp 1649977179
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_669
timestamp 1649977179
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_681
timestamp 1649977179
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1649977179
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1649977179
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_701
timestamp 1649977179
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_713
timestamp 1649977179
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_725
timestamp 1649977179
transform 1 0 67804 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_737
timestamp 1649977179
transform 1 0 68908 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_749
timestamp 1649977179
transform 1 0 70012 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_755
timestamp 1649977179
transform 1 0 70564 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_757
timestamp 1649977179
transform 1 0 70748 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_769
timestamp 1649977179
transform 1 0 71852 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_781
timestamp 1649977179
transform 1 0 72956 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_793
timestamp 1649977179
transform 1 0 74060 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_805
timestamp 1649977179
transform 1 0 75164 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_811
timestamp 1649977179
transform 1 0 75716 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_813
timestamp 1649977179
transform 1 0 75900 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_825
timestamp 1649977179
transform 1 0 77004 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_830
timestamp 1649977179
transform 1 0 77464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_838
timestamp 1649977179
transform 1 0 78200 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_401
timestamp 1649977179
transform 1 0 37996 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_409
timestamp 1649977179
transform 1 0 38732 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_419
timestamp 1649977179
transform 1 0 39652 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_425
timestamp 1649977179
transform 1 0 40204 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_437
timestamp 1649977179
transform 1 0 41308 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_445
timestamp 1649977179
transform 1 0 42044 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_629
timestamp 1649977179
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_641
timestamp 1649977179
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_653
timestamp 1649977179
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1649977179
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1649977179
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_673
timestamp 1649977179
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_685
timestamp 1649977179
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_697
timestamp 1649977179
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_709
timestamp 1649977179
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_721
timestamp 1649977179
transform 1 0 67436 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_727
timestamp 1649977179
transform 1 0 67988 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_729
timestamp 1649977179
transform 1 0 68172 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_741
timestamp 1649977179
transform 1 0 69276 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_753
timestamp 1649977179
transform 1 0 70380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_765
timestamp 1649977179
transform 1 0 71484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_777
timestamp 1649977179
transform 1 0 72588 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_783
timestamp 1649977179
transform 1 0 73140 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_785
timestamp 1649977179
transform 1 0 73324 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_797
timestamp 1649977179
transform 1 0 74428 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_809
timestamp 1649977179
transform 1 0 75532 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_821
timestamp 1649977179
transform 1 0 76636 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_833
timestamp 1649977179
transform 1 0 77740 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_839
timestamp 1649977179
transform 1 0 78292 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_841
timestamp 1649977179
transform 1 0 78476 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_7
timestamp 1649977179
transform 1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_13
timestamp 1649977179
transform 1 0 2300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_25
timestamp 1649977179
transform 1 0 3404 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1649977179
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_405
timestamp 1649977179
transform 1 0 38364 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_408
timestamp 1649977179
transform 1 0 38640 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_416
timestamp 1649977179
transform 1 0 39376 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_427
timestamp 1649977179
transform 1 0 40388 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_625
timestamp 1649977179
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1649977179
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1649977179
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_645
timestamp 1649977179
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_657
timestamp 1649977179
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_669
timestamp 1649977179
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_681
timestamp 1649977179
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1649977179
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1649977179
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_701
timestamp 1649977179
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_713
timestamp 1649977179
transform 1 0 66700 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_725
timestamp 1649977179
transform 1 0 67804 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_737
timestamp 1649977179
transform 1 0 68908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_749
timestamp 1649977179
transform 1 0 70012 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_755
timestamp 1649977179
transform 1 0 70564 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_757
timestamp 1649977179
transform 1 0 70748 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_769
timestamp 1649977179
transform 1 0 71852 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_781
timestamp 1649977179
transform 1 0 72956 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_793
timestamp 1649977179
transform 1 0 74060 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_805
timestamp 1649977179
transform 1 0 75164 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_811
timestamp 1649977179
transform 1 0 75716 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_813
timestamp 1649977179
transform 1 0 75900 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_825
timestamp 1649977179
transform 1 0 77004 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_830
timestamp 1649977179
transform 1 0 77464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_838
timestamp 1649977179
transform 1 0 78200 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_7
timestamp 1649977179
transform 1 0 1748 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_13
timestamp 1649977179
transform 1 0 2300 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_25
timestamp 1649977179
transform 1 0 3404 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_37
timestamp 1649977179
transform 1 0 4508 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_49
timestamp 1649977179
transform 1 0 5612 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_413
timestamp 1649977179
transform 1 0 39100 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_425
timestamp 1649977179
transform 1 0 40204 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_435
timestamp 1649977179
transform 1 0 41124 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_629
timestamp 1649977179
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_641
timestamp 1649977179
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_653
timestamp 1649977179
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_665
timestamp 1649977179
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_671
timestamp 1649977179
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_673
timestamp 1649977179
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_685
timestamp 1649977179
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_697
timestamp 1649977179
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_709
timestamp 1649977179
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_721
timestamp 1649977179
transform 1 0 67436 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_727
timestamp 1649977179
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_729
timestamp 1649977179
transform 1 0 68172 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_741
timestamp 1649977179
transform 1 0 69276 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_753
timestamp 1649977179
transform 1 0 70380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_765
timestamp 1649977179
transform 1 0 71484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_777
timestamp 1649977179
transform 1 0 72588 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_783
timestamp 1649977179
transform 1 0 73140 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_785
timestamp 1649977179
transform 1 0 73324 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_797
timestamp 1649977179
transform 1 0 74428 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_809
timestamp 1649977179
transform 1 0 75532 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_821
timestamp 1649977179
transform 1 0 76636 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_825
timestamp 1649977179
transform 1 0 77004 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_828
timestamp 1649977179
transform 1 0 77280 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_836
timestamp 1649977179
transform 1 0 78016 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_841
timestamp 1649977179
transform 1 0 78476 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_7
timestamp 1649977179
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_13
timestamp 1649977179
transform 1 0 2300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_25
timestamp 1649977179
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_443
timestamp 1649977179
transform 1 0 41860 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_455
timestamp 1649977179
transform 1 0 42964 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_467
timestamp 1649977179
transform 1 0 44068 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_625
timestamp 1649977179
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_637
timestamp 1649977179
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1649977179
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_645
timestamp 1649977179
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_657
timestamp 1649977179
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_669
timestamp 1649977179
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_681
timestamp 1649977179
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1649977179
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1649977179
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_701
timestamp 1649977179
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_713
timestamp 1649977179
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_725
timestamp 1649977179
transform 1 0 67804 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_737
timestamp 1649977179
transform 1 0 68908 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_749
timestamp 1649977179
transform 1 0 70012 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_755
timestamp 1649977179
transform 1 0 70564 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_757
timestamp 1649977179
transform 1 0 70748 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_769
timestamp 1649977179
transform 1 0 71852 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_781
timestamp 1649977179
transform 1 0 72956 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_793
timestamp 1649977179
transform 1 0 74060 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_805
timestamp 1649977179
transform 1 0 75164 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_811
timestamp 1649977179
transform 1 0 75716 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_813
timestamp 1649977179
transform 1 0 75900 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_825
timestamp 1649977179
transform 1 0 77004 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_830
timestamp 1649977179
transform 1 0 77464 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_838
timestamp 1649977179
transform 1 0 78200 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_7
timestamp 1649977179
transform 1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_13
timestamp 1649977179
transform 1 0 2300 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_25
timestamp 1649977179
transform 1 0 3404 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_37
timestamp 1649977179
transform 1 0 4508 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1649977179
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_435
timestamp 1649977179
transform 1 0 41124 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_443
timestamp 1649977179
transform 1 0 41860 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_453
timestamp 1649977179
transform 1 0 42780 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_465
timestamp 1649977179
transform 1 0 43884 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_477
timestamp 1649977179
transform 1 0 44988 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_489
timestamp 1649977179
transform 1 0 46092 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_501
timestamp 1649977179
transform 1 0 47196 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_629
timestamp 1649977179
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_641
timestamp 1649977179
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_653
timestamp 1649977179
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1649977179
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1649977179
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1649977179
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1649977179
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1649977179
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_709
timestamp 1649977179
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1649977179
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1649977179
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_729
timestamp 1649977179
transform 1 0 68172 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_741
timestamp 1649977179
transform 1 0 69276 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_753
timestamp 1649977179
transform 1 0 70380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_765
timestamp 1649977179
transform 1 0 71484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_777
timestamp 1649977179
transform 1 0 72588 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_783
timestamp 1649977179
transform 1 0 73140 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_785
timestamp 1649977179
transform 1 0 73324 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_797
timestamp 1649977179
transform 1 0 74428 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_809
timestamp 1649977179
transform 1 0 75532 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_821
timestamp 1649977179
transform 1 0 76636 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_825
timestamp 1649977179
transform 1 0 77004 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_828
timestamp 1649977179
transform 1 0 77280 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_836
timestamp 1649977179
transform 1 0 78016 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_841
timestamp 1649977179
transform 1 0 78476 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_441
timestamp 1649977179
transform 1 0 41676 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_451
timestamp 1649977179
transform 1 0 42596 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_625
timestamp 1649977179
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1649977179
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1649977179
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1649977179
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1649977179
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_669
timestamp 1649977179
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_681
timestamp 1649977179
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1649977179
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1649977179
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1649977179
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_713
timestamp 1649977179
transform 1 0 66700 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_725
timestamp 1649977179
transform 1 0 67804 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_737
timestamp 1649977179
transform 1 0 68908 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_749
timestamp 1649977179
transform 1 0 70012 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_755
timestamp 1649977179
transform 1 0 70564 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_757
timestamp 1649977179
transform 1 0 70748 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_769
timestamp 1649977179
transform 1 0 71852 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_781
timestamp 1649977179
transform 1 0 72956 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_793
timestamp 1649977179
transform 1 0 74060 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_805
timestamp 1649977179
transform 1 0 75164 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_811
timestamp 1649977179
transform 1 0 75716 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_813
timestamp 1649977179
transform 1 0 75900 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_825
timestamp 1649977179
transform 1 0 77004 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_837
timestamp 1649977179
transform 1 0 78108 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_841
timestamp 1649977179
transform 1 0 78476 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_7
timestamp 1649977179
transform 1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_13
timestamp 1649977179
transform 1 0 2300 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_25
timestamp 1649977179
transform 1 0 3404 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_37
timestamp 1649977179
transform 1 0 4508 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_49
timestamp 1649977179
transform 1 0 5612 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_453
timestamp 1649977179
transform 1 0 42780 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_467
timestamp 1649977179
transform 1 0 44068 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_479
timestamp 1649977179
transform 1 0 45172 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_491
timestamp 1649977179
transform 1 0 46276 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_629
timestamp 1649977179
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_641
timestamp 1649977179
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_653
timestamp 1649977179
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1649977179
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1649977179
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1649977179
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1649977179
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1649977179
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_709
timestamp 1649977179
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1649977179
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1649977179
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_729
timestamp 1649977179
transform 1 0 68172 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_741
timestamp 1649977179
transform 1 0 69276 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_753
timestamp 1649977179
transform 1 0 70380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_765
timestamp 1649977179
transform 1 0 71484 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_777
timestamp 1649977179
transform 1 0 72588 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_783
timestamp 1649977179
transform 1 0 73140 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_785
timestamp 1649977179
transform 1 0 73324 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_797
timestamp 1649977179
transform 1 0 74428 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_809
timestamp 1649977179
transform 1 0 75532 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_821
timestamp 1649977179
transform 1 0 76636 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_825
timestamp 1649977179
transform 1 0 77004 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_828
timestamp 1649977179
transform 1 0 77280 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_836
timestamp 1649977179
transform 1 0 78016 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_841
timestamp 1649977179
transform 1 0 78476 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_7
timestamp 1649977179
transform 1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_13
timestamp 1649977179
transform 1 0 2300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_25
timestamp 1649977179
transform 1 0 3404 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_448
timestamp 1649977179
transform 1 0 42320 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_456
timestamp 1649977179
transform 1 0 43056 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_466
timestamp 1649977179
transform 1 0 43976 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_472
timestamp 1649977179
transform 1 0 44528 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_625
timestamp 1649977179
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1649977179
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1649977179
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1649977179
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1649977179
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1649977179
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1649977179
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1649977179
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1649977179
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1649977179
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_713
timestamp 1649977179
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_725
timestamp 1649977179
transform 1 0 67804 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_737
timestamp 1649977179
transform 1 0 68908 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_749
timestamp 1649977179
transform 1 0 70012 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_755
timestamp 1649977179
transform 1 0 70564 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_757
timestamp 1649977179
transform 1 0 70748 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_769
timestamp 1649977179
transform 1 0 71852 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_781
timestamp 1649977179
transform 1 0 72956 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_793
timestamp 1649977179
transform 1 0 74060 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_805
timestamp 1649977179
transform 1 0 75164 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_811
timestamp 1649977179
transform 1 0 75716 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_813
timestamp 1649977179
transform 1 0 75900 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_825
timestamp 1649977179
transform 1 0 77004 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_830
timestamp 1649977179
transform 1 0 77464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_838
timestamp 1649977179
transform 1 0 78200 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_7
timestamp 1649977179
transform 1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_13
timestamp 1649977179
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_25
timestamp 1649977179
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_37
timestamp 1649977179
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1649977179
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_457
timestamp 1649977179
transform 1 0 43148 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_464
timestamp 1649977179
transform 1 0 43792 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_474
timestamp 1649977179
transform 1 0 44712 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_486
timestamp 1649977179
transform 1 0 45816 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_498
timestamp 1649977179
transform 1 0 46920 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_629
timestamp 1649977179
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_641
timestamp 1649977179
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_653
timestamp 1649977179
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1649977179
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1649977179
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1649977179
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_685
timestamp 1649977179
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_697
timestamp 1649977179
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_709
timestamp 1649977179
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_721
timestamp 1649977179
transform 1 0 67436 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_727
timestamp 1649977179
transform 1 0 67988 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_729
timestamp 1649977179
transform 1 0 68172 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_741
timestamp 1649977179
transform 1 0 69276 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_753
timestamp 1649977179
transform 1 0 70380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_765
timestamp 1649977179
transform 1 0 71484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_777
timestamp 1649977179
transform 1 0 72588 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_783
timestamp 1649977179
transform 1 0 73140 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_785
timestamp 1649977179
transform 1 0 73324 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_797
timestamp 1649977179
transform 1 0 74428 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_809
timestamp 1649977179
transform 1 0 75532 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_821
timestamp 1649977179
transform 1 0 76636 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_825
timestamp 1649977179
transform 1 0 77004 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_828
timestamp 1649977179
transform 1 0 77280 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_836
timestamp 1649977179
transform 1 0 78016 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_841
timestamp 1649977179
transform 1 0 78476 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_7
timestamp 1649977179
transform 1 0 1748 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_13
timestamp 1649977179
transform 1 0 2300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_25
timestamp 1649977179
transform 1 0 3404 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_463
timestamp 1649977179
transform 1 0 43700 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_466
timestamp 1649977179
transform 1 0 43976 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_472
timestamp 1649977179
transform 1 0 44528 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_625
timestamp 1649977179
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1649977179
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1649977179
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1649977179
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1649977179
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1649977179
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_681
timestamp 1649977179
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1649977179
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1649977179
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_701
timestamp 1649977179
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_713
timestamp 1649977179
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_725
timestamp 1649977179
transform 1 0 67804 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_737
timestamp 1649977179
transform 1 0 68908 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_749
timestamp 1649977179
transform 1 0 70012 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_755
timestamp 1649977179
transform 1 0 70564 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_757
timestamp 1649977179
transform 1 0 70748 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_769
timestamp 1649977179
transform 1 0 71852 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_781
timestamp 1649977179
transform 1 0 72956 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_793
timestamp 1649977179
transform 1 0 74060 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_805
timestamp 1649977179
transform 1 0 75164 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_811
timestamp 1649977179
transform 1 0 75716 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_813
timestamp 1649977179
transform 1 0 75900 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_825
timestamp 1649977179
transform 1 0 77004 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_830
timestamp 1649977179
transform 1 0 77464 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_838
timestamp 1649977179
transform 1 0 78200 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_464
timestamp 1649977179
transform 1 0 43792 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_472
timestamp 1649977179
transform 1 0 44528 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_482
timestamp 1649977179
transform 1 0 45448 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_488
timestamp 1649977179
transform 1 0 46000 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_494
timestamp 1649977179
transform 1 0 46552 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_502
timestamp 1649977179
transform 1 0 47288 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1649977179
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1649977179
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1649977179
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1649977179
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1649977179
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1649977179
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1649977179
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1649977179
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_709
timestamp 1649977179
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_721
timestamp 1649977179
transform 1 0 67436 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_727
timestamp 1649977179
transform 1 0 67988 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_729
timestamp 1649977179
transform 1 0 68172 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_741
timestamp 1649977179
transform 1 0 69276 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_753
timestamp 1649977179
transform 1 0 70380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_765
timestamp 1649977179
transform 1 0 71484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_777
timestamp 1649977179
transform 1 0 72588 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_783
timestamp 1649977179
transform 1 0 73140 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_785
timestamp 1649977179
transform 1 0 73324 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_797
timestamp 1649977179
transform 1 0 74428 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_809
timestamp 1649977179
transform 1 0 75532 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_821
timestamp 1649977179
transform 1 0 76636 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_833
timestamp 1649977179
transform 1 0 77740 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_839
timestamp 1649977179
transform 1 0 78292 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_841
timestamp 1649977179
transform 1 0 78476 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_7
timestamp 1649977179
transform 1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_13
timestamp 1649977179
transform 1 0 2300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_25
timestamp 1649977179
transform 1 0 3404 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_481
timestamp 1649977179
transform 1 0 45356 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_485
timestamp 1649977179
transform 1 0 45724 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_490
timestamp 1649977179
transform 1 0 46184 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_496
timestamp 1649977179
transform 1 0 46736 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_508
timestamp 1649977179
transform 1 0 47840 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_520
timestamp 1649977179
transform 1 0 48944 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1649977179
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1649977179
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1649977179
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1649977179
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1649977179
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1649977179
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1649977179
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1649977179
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1649977179
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_701
timestamp 1649977179
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_713
timestamp 1649977179
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_725
timestamp 1649977179
transform 1 0 67804 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_737
timestamp 1649977179
transform 1 0 68908 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_749
timestamp 1649977179
transform 1 0 70012 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_755
timestamp 1649977179
transform 1 0 70564 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_757
timestamp 1649977179
transform 1 0 70748 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_769
timestamp 1649977179
transform 1 0 71852 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_781
timestamp 1649977179
transform 1 0 72956 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_793
timestamp 1649977179
transform 1 0 74060 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_805
timestamp 1649977179
transform 1 0 75164 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_811
timestamp 1649977179
transform 1 0 75716 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_813
timestamp 1649977179
transform 1 0 75900 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_825
timestamp 1649977179
transform 1 0 77004 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_830
timestamp 1649977179
transform 1 0 77464 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_838
timestamp 1649977179
transform 1 0 78200 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_7
timestamp 1649977179
transform 1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_13
timestamp 1649977179
transform 1 0 2300 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_25
timestamp 1649977179
transform 1 0 3404 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_37
timestamp 1649977179
transform 1 0 4508 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_49
timestamp 1649977179
transform 1 0 5612 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_479
timestamp 1649977179
transform 1 0 45172 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_487
timestamp 1649977179
transform 1 0 45908 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_493
timestamp 1649977179
transform 1 0 46460 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_498
timestamp 1649977179
transform 1 0 46920 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_507
timestamp 1649977179
transform 1 0 47748 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_519
timestamp 1649977179
transform 1 0 48852 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_531
timestamp 1649977179
transform 1 0 49956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_543
timestamp 1649977179
transform 1 0 51060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_555
timestamp 1649977179
transform 1 0 52164 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1649977179
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1649977179
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1649977179
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1649977179
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1649977179
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1649977179
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1649977179
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1649977179
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_709
timestamp 1649977179
transform 1 0 66332 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_721
timestamp 1649977179
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_727
timestamp 1649977179
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_729
timestamp 1649977179
transform 1 0 68172 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_741
timestamp 1649977179
transform 1 0 69276 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_753
timestamp 1649977179
transform 1 0 70380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_765
timestamp 1649977179
transform 1 0 71484 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_777
timestamp 1649977179
transform 1 0 72588 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_783
timestamp 1649977179
transform 1 0 73140 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_785
timestamp 1649977179
transform 1 0 73324 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_797
timestamp 1649977179
transform 1 0 74428 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_809
timestamp 1649977179
transform 1 0 75532 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_821
timestamp 1649977179
transform 1 0 76636 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_825
timestamp 1649977179
transform 1 0 77004 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_828
timestamp 1649977179
transform 1 0 77280 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_836
timestamp 1649977179
transform 1 0 78016 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_841
timestamp 1649977179
transform 1 0 78476 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_7
timestamp 1649977179
transform 1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_13
timestamp 1649977179
transform 1 0 2300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_25
timestamp 1649977179
transform 1 0 3404 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_495
timestamp 1649977179
transform 1 0 46644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_506
timestamp 1649977179
transform 1 0 47656 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_512
timestamp 1649977179
transform 1 0 48208 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_524
timestamp 1649977179
transform 1 0 49312 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_625
timestamp 1649977179
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1649977179
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1649977179
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1649977179
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1649977179
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_669
timestamp 1649977179
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_681
timestamp 1649977179
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1649977179
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1649977179
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1649977179
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_713
timestamp 1649977179
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_725
timestamp 1649977179
transform 1 0 67804 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_737
timestamp 1649977179
transform 1 0 68908 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_749
timestamp 1649977179
transform 1 0 70012 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_755
timestamp 1649977179
transform 1 0 70564 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_757
timestamp 1649977179
transform 1 0 70748 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_769
timestamp 1649977179
transform 1 0 71852 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_781
timestamp 1649977179
transform 1 0 72956 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_793
timestamp 1649977179
transform 1 0 74060 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_805
timestamp 1649977179
transform 1 0 75164 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_811
timestamp 1649977179
transform 1 0 75716 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_813
timestamp 1649977179
transform 1 0 75900 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_825
timestamp 1649977179
transform 1 0 77004 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_830
timestamp 1649977179
transform 1 0 77464 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_838
timestamp 1649977179
transform 1 0 78200 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_7
timestamp 1649977179
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_13
timestamp 1649977179
transform 1 0 2300 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_25
timestamp 1649977179
transform 1 0 3404 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_37
timestamp 1649977179
transform 1 0 4508 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_49
timestamp 1649977179
transform 1 0 5612 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_493
timestamp 1649977179
transform 1 0 46460 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_507
timestamp 1649977179
transform 1 0 47748 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_519
timestamp 1649977179
transform 1 0 48852 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_531
timestamp 1649977179
transform 1 0 49956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_543
timestamp 1649977179
transform 1 0 51060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_555
timestamp 1649977179
transform 1 0 52164 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_629
timestamp 1649977179
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_641
timestamp 1649977179
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_653
timestamp 1649977179
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1649977179
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1649977179
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_673
timestamp 1649977179
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_685
timestamp 1649977179
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_697
timestamp 1649977179
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_709
timestamp 1649977179
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1649977179
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1649977179
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_729
timestamp 1649977179
transform 1 0 68172 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_741
timestamp 1649977179
transform 1 0 69276 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_753
timestamp 1649977179
transform 1 0 70380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_765
timestamp 1649977179
transform 1 0 71484 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_777
timestamp 1649977179
transform 1 0 72588 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_783
timestamp 1649977179
transform 1 0 73140 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_785
timestamp 1649977179
transform 1 0 73324 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_797
timestamp 1649977179
transform 1 0 74428 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_809
timestamp 1649977179
transform 1 0 75532 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_821
timestamp 1649977179
transform 1 0 76636 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_825
timestamp 1649977179
transform 1 0 77004 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_828
timestamp 1649977179
transform 1 0 77280 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_836
timestamp 1649977179
transform 1 0 78016 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_841
timestamp 1649977179
transform 1 0 78476 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_497
timestamp 1649977179
transform 1 0 46828 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_503
timestamp 1649977179
transform 1 0 47380 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_509
timestamp 1649977179
transform 1 0 47932 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_514
timestamp 1649977179
transform 1 0 48392 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_520
timestamp 1649977179
transform 1 0 48944 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_625
timestamp 1649977179
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1649977179
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1649977179
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_645
timestamp 1649977179
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_657
timestamp 1649977179
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_669
timestamp 1649977179
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_681
timestamp 1649977179
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1649977179
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1649977179
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_701
timestamp 1649977179
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_713
timestamp 1649977179
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_725
timestamp 1649977179
transform 1 0 67804 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_737
timestamp 1649977179
transform 1 0 68908 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_749
timestamp 1649977179
transform 1 0 70012 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_755
timestamp 1649977179
transform 1 0 70564 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_757
timestamp 1649977179
transform 1 0 70748 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_769
timestamp 1649977179
transform 1 0 71852 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_781
timestamp 1649977179
transform 1 0 72956 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_793
timestamp 1649977179
transform 1 0 74060 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_805
timestamp 1649977179
transform 1 0 75164 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_811
timestamp 1649977179
transform 1 0 75716 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_813
timestamp 1649977179
transform 1 0 75900 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_825
timestamp 1649977179
transform 1 0 77004 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_837
timestamp 1649977179
transform 1 0 78108 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_841
timestamp 1649977179
transform 1 0 78476 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_7
timestamp 1649977179
transform 1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_13
timestamp 1649977179
transform 1 0 2300 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_25
timestamp 1649977179
transform 1 0 3404 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_37
timestamp 1649977179
transform 1 0 4508 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_49
timestamp 1649977179
transform 1 0 5612 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_510
timestamp 1649977179
transform 1 0 48024 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_522
timestamp 1649977179
transform 1 0 49128 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_528
timestamp 1649977179
transform 1 0 49680 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_540
timestamp 1649977179
transform 1 0 50784 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_552
timestamp 1649977179
transform 1 0 51888 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_629
timestamp 1649977179
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_641
timestamp 1649977179
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_653
timestamp 1649977179
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1649977179
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1649977179
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_673
timestamp 1649977179
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_685
timestamp 1649977179
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_697
timestamp 1649977179
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_709
timestamp 1649977179
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_721
timestamp 1649977179
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1649977179
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_729
timestamp 1649977179
transform 1 0 68172 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_741
timestamp 1649977179
transform 1 0 69276 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_753
timestamp 1649977179
transform 1 0 70380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_765
timestamp 1649977179
transform 1 0 71484 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_777
timestamp 1649977179
transform 1 0 72588 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_783
timestamp 1649977179
transform 1 0 73140 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_785
timestamp 1649977179
transform 1 0 73324 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_797
timestamp 1649977179
transform 1 0 74428 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_809
timestamp 1649977179
transform 1 0 75532 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_821
timestamp 1649977179
transform 1 0 76636 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_825
timestamp 1649977179
transform 1 0 77004 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_828
timestamp 1649977179
transform 1 0 77280 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_836
timestamp 1649977179
transform 1 0 78016 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_841
timestamp 1649977179
transform 1 0 78476 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_7
timestamp 1649977179
transform 1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_13
timestamp 1649977179
transform 1 0 2300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_25
timestamp 1649977179
transform 1 0 3404 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_509
timestamp 1649977179
transform 1 0 47932 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_512
timestamp 1649977179
transform 1 0 48208 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_524
timestamp 1649977179
transform 1 0 49312 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_625
timestamp 1649977179
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1649977179
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1649977179
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_645
timestamp 1649977179
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_657
timestamp 1649977179
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_669
timestamp 1649977179
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_681
timestamp 1649977179
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1649977179
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1649977179
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_701
timestamp 1649977179
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_713
timestamp 1649977179
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_725
timestamp 1649977179
transform 1 0 67804 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_737
timestamp 1649977179
transform 1 0 68908 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_749
timestamp 1649977179
transform 1 0 70012 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_755
timestamp 1649977179
transform 1 0 70564 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_757
timestamp 1649977179
transform 1 0 70748 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_769
timestamp 1649977179
transform 1 0 71852 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_781
timestamp 1649977179
transform 1 0 72956 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_793
timestamp 1649977179
transform 1 0 74060 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_805
timestamp 1649977179
transform 1 0 75164 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_811
timestamp 1649977179
transform 1 0 75716 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_813
timestamp 1649977179
transform 1 0 75900 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_825
timestamp 1649977179
transform 1 0 77004 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_830
timestamp 1649977179
transform 1 0 77464 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_838
timestamp 1649977179
transform 1 0 78200 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_7
timestamp 1649977179
transform 1 0 1748 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_13
timestamp 1649977179
transform 1 0 2300 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_25
timestamp 1649977179
transform 1 0 3404 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_37
timestamp 1649977179
transform 1 0 4508 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_49
timestamp 1649977179
transform 1 0 5612 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_525
timestamp 1649977179
transform 1 0 49404 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_85_547
timestamp 1649977179
transform 1 0 51428 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_629
timestamp 1649977179
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_641
timestamp 1649977179
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_653
timestamp 1649977179
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1649977179
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1649977179
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_673
timestamp 1649977179
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_685
timestamp 1649977179
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_697
timestamp 1649977179
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_709
timestamp 1649977179
transform 1 0 66332 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_721
timestamp 1649977179
transform 1 0 67436 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_727
timestamp 1649977179
transform 1 0 67988 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_729
timestamp 1649977179
transform 1 0 68172 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_741
timestamp 1649977179
transform 1 0 69276 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_753
timestamp 1649977179
transform 1 0 70380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_765
timestamp 1649977179
transform 1 0 71484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_777
timestamp 1649977179
transform 1 0 72588 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_783
timestamp 1649977179
transform 1 0 73140 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_785
timestamp 1649977179
transform 1 0 73324 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_797
timestamp 1649977179
transform 1 0 74428 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_809
timestamp 1649977179
transform 1 0 75532 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_817
timestamp 1649977179
transform 1 0 76268 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_822
timestamp 1649977179
transform 1 0 76728 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_836
timestamp 1649977179
transform 1 0 78016 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_841
timestamp 1649977179
transform 1 0 78476 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_7
timestamp 1649977179
transform 1 0 1748 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_19
timestamp 1649977179
transform 1 0 2852 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_528
timestamp 1649977179
transform 1 0 49680 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_541
timestamp 1649977179
transform 1 0 50876 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_547
timestamp 1649977179
transform 1 0 51428 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_559
timestamp 1649977179
transform 1 0 52532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_571
timestamp 1649977179
transform 1 0 53636 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_583
timestamp 1649977179
transform 1 0 54740 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_625
timestamp 1649977179
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1649977179
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1649977179
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_645
timestamp 1649977179
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_657
timestamp 1649977179
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_669
timestamp 1649977179
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_681
timestamp 1649977179
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1649977179
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1649977179
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_701
timestamp 1649977179
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_713
timestamp 1649977179
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_725
timestamp 1649977179
transform 1 0 67804 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_737
timestamp 1649977179
transform 1 0 68908 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_749
timestamp 1649977179
transform 1 0 70012 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_755
timestamp 1649977179
transform 1 0 70564 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_757
timestamp 1649977179
transform 1 0 70748 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_769
timestamp 1649977179
transform 1 0 71852 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_781
timestamp 1649977179
transform 1 0 72956 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_793
timestamp 1649977179
transform 1 0 74060 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_805
timestamp 1649977179
transform 1 0 75164 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_811
timestamp 1649977179
transform 1 0 75716 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_813
timestamp 1649977179
transform 1 0 75900 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_825
timestamp 1649977179
transform 1 0 77004 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_838
timestamp 1649977179
transform 1 0 78200 0 1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_5
timestamp 1649977179
transform 1 0 1564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_17
timestamp 1649977179
transform 1 0 2668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_29
timestamp 1649977179
transform 1 0 3772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_41
timestamp 1649977179
transform 1 0 4876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1649977179
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_531
timestamp 1649977179
transform 1 0 49956 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_543
timestamp 1649977179
transform 1 0 51060 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_549
timestamp 1649977179
transform 1 0 51612 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_557
timestamp 1649977179
transform 1 0 52348 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_563
timestamp 1649977179
transform 1 0 52900 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_575
timestamp 1649977179
transform 1 0 54004 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_587
timestamp 1649977179
transform 1 0 55108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_599
timestamp 1649977179
transform 1 0 56212 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_611
timestamp 1649977179
transform 1 0 57316 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_629
timestamp 1649977179
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_641
timestamp 1649977179
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_653
timestamp 1649977179
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1649977179
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1649977179
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_673
timestamp 1649977179
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_685
timestamp 1649977179
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_697
timestamp 1649977179
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_709
timestamp 1649977179
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_721
timestamp 1649977179
transform 1 0 67436 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_727
timestamp 1649977179
transform 1 0 67988 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_729
timestamp 1649977179
transform 1 0 68172 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_741
timestamp 1649977179
transform 1 0 69276 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_753
timestamp 1649977179
transform 1 0 70380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_765
timestamp 1649977179
transform 1 0 71484 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_777
timestamp 1649977179
transform 1 0 72588 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_783
timestamp 1649977179
transform 1 0 73140 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_785
timestamp 1649977179
transform 1 0 73324 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_797
timestamp 1649977179
transform 1 0 74428 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_809
timestamp 1649977179
transform 1 0 75532 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_821
timestamp 1649977179
transform 1 0 76636 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_827
timestamp 1649977179
transform 1 0 77188 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_830
timestamp 1649977179
transform 1 0 77464 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_836
timestamp 1649977179
transform 1 0 78016 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_841
timestamp 1649977179
transform 1 0 78476 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_7
timestamp 1649977179
transform 1 0 1748 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_13
timestamp 1649977179
transform 1 0 2300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_88_25
timestamp 1649977179
transform 1 0 3404 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_536
timestamp 1649977179
transform 1 0 50416 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_548
timestamp 1649977179
transform 1 0 51520 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_554
timestamp 1649977179
transform 1 0 52072 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_88_570
timestamp 1649977179
transform 1 0 53544 0 1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_576
timestamp 1649977179
transform 1 0 54096 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_625
timestamp 1649977179
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1649977179
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1649977179
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_645
timestamp 1649977179
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_657
timestamp 1649977179
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_669
timestamp 1649977179
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_681
timestamp 1649977179
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1649977179
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1649977179
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_701
timestamp 1649977179
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_713
timestamp 1649977179
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_725
timestamp 1649977179
transform 1 0 67804 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_737
timestamp 1649977179
transform 1 0 68908 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_749
timestamp 1649977179
transform 1 0 70012 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_755
timestamp 1649977179
transform 1 0 70564 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_757
timestamp 1649977179
transform 1 0 70748 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_769
timestamp 1649977179
transform 1 0 71852 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_781
timestamp 1649977179
transform 1 0 72956 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_793
timestamp 1649977179
transform 1 0 74060 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_805
timestamp 1649977179
transform 1 0 75164 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_811
timestamp 1649977179
transform 1 0 75716 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_813
timestamp 1649977179
transform 1 0 75900 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_88_825
timestamp 1649977179
transform 1 0 77004 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_838
timestamp 1649977179
transform 1 0 78200 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_7
timestamp 1649977179
transform 1 0 1748 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_13
timestamp 1649977179
transform 1 0 2300 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_25
timestamp 1649977179
transform 1 0 3404 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_37
timestamp 1649977179
transform 1 0 4508 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_49
timestamp 1649977179
transform 1 0 5612 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_565
timestamp 1649977179
transform 1 0 53084 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_576
timestamp 1649977179
transform 1 0 54096 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_588
timestamp 1649977179
transform 1 0 55200 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_600
timestamp 1649977179
transform 1 0 56304 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_612
timestamp 1649977179
transform 1 0 57408 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_629
timestamp 1649977179
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_641
timestamp 1649977179
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_653
timestamp 1649977179
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1649977179
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1649977179
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_673
timestamp 1649977179
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_685
timestamp 1649977179
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_697
timestamp 1649977179
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_709
timestamp 1649977179
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_721
timestamp 1649977179
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_727
timestamp 1649977179
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_729
timestamp 1649977179
transform 1 0 68172 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_741
timestamp 1649977179
transform 1 0 69276 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_753
timestamp 1649977179
transform 1 0 70380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_765
timestamp 1649977179
transform 1 0 71484 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_777
timestamp 1649977179
transform 1 0 72588 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_783
timestamp 1649977179
transform 1 0 73140 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_785
timestamp 1649977179
transform 1 0 73324 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_797
timestamp 1649977179
transform 1 0 74428 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_809
timestamp 1649977179
transform 1 0 75532 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_817
timestamp 1649977179
transform 1 0 76268 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_822
timestamp 1649977179
transform 1 0 76728 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_836
timestamp 1649977179
transform 1 0 78016 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_841
timestamp 1649977179
transform 1 0 78476 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_7
timestamp 1649977179
transform 1 0 1748 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_13
timestamp 1649977179
transform 1 0 2300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_25
timestamp 1649977179
transform 1 0 3404 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_547
timestamp 1649977179
transform 1 0 51428 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_559
timestamp 1649977179
transform 1 0 52532 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_573
timestamp 1649977179
transform 1 0 53820 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_579
timestamp 1649977179
transform 1 0 54372 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_625
timestamp 1649977179
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1649977179
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1649977179
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_645
timestamp 1649977179
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_657
timestamp 1649977179
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_669
timestamp 1649977179
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_681
timestamp 1649977179
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1649977179
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1649977179
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_701
timestamp 1649977179
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_713
timestamp 1649977179
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_725
timestamp 1649977179
transform 1 0 67804 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_737
timestamp 1649977179
transform 1 0 68908 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_749
timestamp 1649977179
transform 1 0 70012 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_755
timestamp 1649977179
transform 1 0 70564 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_757
timestamp 1649977179
transform 1 0 70748 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_769
timestamp 1649977179
transform 1 0 71852 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_781
timestamp 1649977179
transform 1 0 72956 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_793
timestamp 1649977179
transform 1 0 74060 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_805
timestamp 1649977179
transform 1 0 75164 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_811
timestamp 1649977179
transform 1 0 75716 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_813
timestamp 1649977179
transform 1 0 75900 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_821
timestamp 1649977179
transform 1 0 76636 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_824
timestamp 1649977179
transform 1 0 76912 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_838
timestamp 1649977179
transform 1 0 78200 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_7
timestamp 1649977179
transform 1 0 1748 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_19
timestamp 1649977179
transform 1 0 2852 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_31
timestamp 1649977179
transform 1 0 3956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_43
timestamp 1649977179
transform 1 0 5060 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_544
timestamp 1649977179
transform 1 0 51152 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_556
timestamp 1649977179
transform 1 0 52256 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_575
timestamp 1649977179
transform 1 0 54004 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_587
timestamp 1649977179
transform 1 0 55108 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_593
timestamp 1649977179
transform 1 0 55660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_605
timestamp 1649977179
transform 1 0 56764 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_613
timestamp 1649977179
transform 1 0 57500 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_629
timestamp 1649977179
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_641
timestamp 1649977179
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_653
timestamp 1649977179
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1649977179
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1649977179
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_673
timestamp 1649977179
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_685
timestamp 1649977179
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_697
timestamp 1649977179
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_709
timestamp 1649977179
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1649977179
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1649977179
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_729
timestamp 1649977179
transform 1 0 68172 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_741
timestamp 1649977179
transform 1 0 69276 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_753
timestamp 1649977179
transform 1 0 70380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_765
timestamp 1649977179
transform 1 0 71484 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_777
timestamp 1649977179
transform 1 0 72588 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_783
timestamp 1649977179
transform 1 0 73140 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_785
timestamp 1649977179
transform 1 0 73324 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_797
timestamp 1649977179
transform 1 0 74428 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_809
timestamp 1649977179
transform 1 0 75532 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_821
timestamp 1649977179
transform 1 0 76636 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_825
timestamp 1649977179
transform 1 0 77004 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_836
timestamp 1649977179
transform 1 0 78016 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_841
timestamp 1649977179
transform 1 0 78476 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_5
timestamp 1649977179
transform 1 0 1564 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_17
timestamp 1649977179
transform 1 0 2668 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_25
timestamp 1649977179
transform 1 0 3404 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_553
timestamp 1649977179
transform 1 0 51980 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_558
timestamp 1649977179
transform 1 0 52440 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_564
timestamp 1649977179
transform 1 0 52992 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_578
timestamp 1649977179
transform 1 0 54280 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_584
timestamp 1649977179
transform 1 0 54832 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_625
timestamp 1649977179
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1649977179
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1649977179
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_645
timestamp 1649977179
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_657
timestamp 1649977179
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_669
timestamp 1649977179
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_681
timestamp 1649977179
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1649977179
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1649977179
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_701
timestamp 1649977179
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_713
timestamp 1649977179
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_725
timestamp 1649977179
transform 1 0 67804 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_737
timestamp 1649977179
transform 1 0 68908 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_749
timestamp 1649977179
transform 1 0 70012 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_755
timestamp 1649977179
transform 1 0 70564 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_757
timestamp 1649977179
transform 1 0 70748 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_769
timestamp 1649977179
transform 1 0 71852 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_781
timestamp 1649977179
transform 1 0 72956 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_793
timestamp 1649977179
transform 1 0 74060 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_805
timestamp 1649977179
transform 1 0 75164 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_811
timestamp 1649977179
transform 1 0 75716 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_813
timestamp 1649977179
transform 1 0 75900 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_825
timestamp 1649977179
transform 1 0 77004 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_829
timestamp 1649977179
transform 1 0 77372 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_832
timestamp 1649977179
transform 1 0 77648 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_838
timestamp 1649977179
transform 1 0 78200 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_7
timestamp 1649977179
transform 1 0 1748 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_13
timestamp 1649977179
transform 1 0 2300 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_25
timestamp 1649977179
transform 1 0 3404 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_37
timestamp 1649977179
transform 1 0 4508 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_49
timestamp 1649977179
transform 1 0 5612 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_572
timestamp 1649977179
transform 1 0 53728 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_584
timestamp 1649977179
transform 1 0 54832 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_590
timestamp 1649977179
transform 1 0 55384 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_602
timestamp 1649977179
transform 1 0 56488 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_614
timestamp 1649977179
transform 1 0 57592 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_629
timestamp 1649977179
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_641
timestamp 1649977179
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_653
timestamp 1649977179
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1649977179
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1649977179
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_673
timestamp 1649977179
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_685
timestamp 1649977179
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_697
timestamp 1649977179
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_709
timestamp 1649977179
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1649977179
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1649977179
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_729
timestamp 1649977179
transform 1 0 68172 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_741
timestamp 1649977179
transform 1 0 69276 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_753
timestamp 1649977179
transform 1 0 70380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_765
timestamp 1649977179
transform 1 0 71484 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_777
timestamp 1649977179
transform 1 0 72588 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_783
timestamp 1649977179
transform 1 0 73140 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_785
timestamp 1649977179
transform 1 0 73324 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_797
timestamp 1649977179
transform 1 0 74428 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_809
timestamp 1649977179
transform 1 0 75532 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_821
timestamp 1649977179
transform 1 0 76636 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_825
timestamp 1649977179
transform 1 0 77004 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_836
timestamp 1649977179
transform 1 0 78016 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_841
timestamp 1649977179
transform 1 0 78476 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_7
timestamp 1649977179
transform 1 0 1748 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_13
timestamp 1649977179
transform 1 0 2300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_25
timestamp 1649977179
transform 1 0 3404 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_574
timestamp 1649977179
transform 1 0 53912 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_580
timestamp 1649977179
transform 1 0 54464 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_625
timestamp 1649977179
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1649977179
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1649977179
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_645
timestamp 1649977179
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_657
timestamp 1649977179
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_669
timestamp 1649977179
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_681
timestamp 1649977179
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1649977179
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1649977179
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_701
timestamp 1649977179
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_713
timestamp 1649977179
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_725
timestamp 1649977179
transform 1 0 67804 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_737
timestamp 1649977179
transform 1 0 68908 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_749
timestamp 1649977179
transform 1 0 70012 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_755
timestamp 1649977179
transform 1 0 70564 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_757
timestamp 1649977179
transform 1 0 70748 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_769
timestamp 1649977179
transform 1 0 71852 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_781
timestamp 1649977179
transform 1 0 72956 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_793
timestamp 1649977179
transform 1 0 74060 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_805
timestamp 1649977179
transform 1 0 75164 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_811
timestamp 1649977179
transform 1 0 75716 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_813
timestamp 1649977179
transform 1 0 75900 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_821
timestamp 1649977179
transform 1 0 76636 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_824
timestamp 1649977179
transform 1 0 76912 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_838
timestamp 1649977179
transform 1 0 78200 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_7
timestamp 1649977179
transform 1 0 1748 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_95_13
timestamp 1649977179
transform 1 0 2300 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_25
timestamp 1649977179
transform 1 0 3404 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_37
timestamp 1649977179
transform 1 0 4508 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_49
timestamp 1649977179
transform 1 0 5612 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_593
timestamp 1649977179
transform 1 0 55660 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_605
timestamp 1649977179
transform 1 0 56764 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_611
timestamp 1649977179
transform 1 0 57316 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_629
timestamp 1649977179
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_641
timestamp 1649977179
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_653
timestamp 1649977179
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1649977179
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1649977179
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_673
timestamp 1649977179
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_685
timestamp 1649977179
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_697
timestamp 1649977179
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_709
timestamp 1649977179
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_721
timestamp 1649977179
transform 1 0 67436 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_727
timestamp 1649977179
transform 1 0 67988 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_729
timestamp 1649977179
transform 1 0 68172 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_741
timestamp 1649977179
transform 1 0 69276 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_753
timestamp 1649977179
transform 1 0 70380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_765
timestamp 1649977179
transform 1 0 71484 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_777
timestamp 1649977179
transform 1 0 72588 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_783
timestamp 1649977179
transform 1 0 73140 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_785
timestamp 1649977179
transform 1 0 73324 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_797
timestamp 1649977179
transform 1 0 74428 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_809
timestamp 1649977179
transform 1 0 75532 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_821
timestamp 1649977179
transform 1 0 76636 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_825
timestamp 1649977179
transform 1 0 77004 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_836
timestamp 1649977179
transform 1 0 78016 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_841
timestamp 1649977179
transform 1 0 78476 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_7
timestamp 1649977179
transform 1 0 1748 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_19
timestamp 1649977179
transform 1 0 2852 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_96_597
timestamp 1649977179
transform 1 0 56028 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_610
timestamp 1649977179
transform 1 0 57224 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_624
timestamp 1649977179
transform 1 0 58512 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_630
timestamp 1649977179
transform 1 0 59064 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_642
timestamp 1649977179
transform 1 0 60168 0 1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_645
timestamp 1649977179
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_657
timestamp 1649977179
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_669
timestamp 1649977179
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_681
timestamp 1649977179
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1649977179
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1649977179
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_701
timestamp 1649977179
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_713
timestamp 1649977179
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_725
timestamp 1649977179
transform 1 0 67804 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_737
timestamp 1649977179
transform 1 0 68908 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_749
timestamp 1649977179
transform 1 0 70012 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_755
timestamp 1649977179
transform 1 0 70564 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_757
timestamp 1649977179
transform 1 0 70748 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_769
timestamp 1649977179
transform 1 0 71852 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_781
timestamp 1649977179
transform 1 0 72956 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_793
timestamp 1649977179
transform 1 0 74060 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_805
timestamp 1649977179
transform 1 0 75164 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_811
timestamp 1649977179
transform 1 0 75716 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_813
timestamp 1649977179
transform 1 0 75900 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_825
timestamp 1649977179
transform 1 0 77004 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_831
timestamp 1649977179
transform 1 0 77556 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_838
timestamp 1649977179
transform 1 0 78200 0 1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_5
timestamp 1649977179
transform 1 0 1564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_17
timestamp 1649977179
transform 1 0 2668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_29
timestamp 1649977179
transform 1 0 3772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_41
timestamp 1649977179
transform 1 0 4876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_53
timestamp 1649977179
transform 1 0 5980 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1649977179
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1649977179
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1649977179
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1649977179
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_97_595
timestamp 1649977179
transform 1 0 55844 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_607
timestamp 1649977179
transform 1 0 56948 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_625
timestamp 1649977179
transform 1 0 58604 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_631
timestamp 1649977179
transform 1 0 59156 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_643
timestamp 1649977179
transform 1 0 60260 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_648
timestamp 1649977179
transform 1 0 60720 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_654
timestamp 1649977179
transform 1 0 61272 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_666
timestamp 1649977179
transform 1 0 62376 0 -1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_97_673
timestamp 1649977179
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_685
timestamp 1649977179
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_697
timestamp 1649977179
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_709
timestamp 1649977179
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_721
timestamp 1649977179
transform 1 0 67436 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_727
timestamp 1649977179
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_729
timestamp 1649977179
transform 1 0 68172 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_741
timestamp 1649977179
transform 1 0 69276 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_753
timestamp 1649977179
transform 1 0 70380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_765
timestamp 1649977179
transform 1 0 71484 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_777
timestamp 1649977179
transform 1 0 72588 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_783
timestamp 1649977179
transform 1 0 73140 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_785
timestamp 1649977179
transform 1 0 73324 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_797
timestamp 1649977179
transform 1 0 74428 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_809
timestamp 1649977179
transform 1 0 75532 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_821
timestamp 1649977179
transform 1 0 76636 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_833
timestamp 1649977179
transform 1 0 77740 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_836
timestamp 1649977179
transform 1 0 78016 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_841
timestamp 1649977179
transform 1 0 78476 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_7
timestamp 1649977179
transform 1 0 1748 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_13
timestamp 1649977179
transform 1 0 2300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_25
timestamp 1649977179
transform 1 0 3404 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1649977179
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1649977179
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1649977179
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1649977179
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1649977179
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1649977179
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1649977179
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1649977179
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1649977179
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1649977179
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1649977179
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1649977179
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1649977179
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1649977179
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1649977179
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1649977179
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1649977179
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1649977179
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1649977179
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_595
timestamp 1649977179
transform 1 0 55844 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_598
timestamp 1649977179
transform 1 0 56120 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_610
timestamp 1649977179
transform 1 0 57224 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_622
timestamp 1649977179
transform 1 0 58328 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_628
timestamp 1649977179
transform 1 0 58880 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_640
timestamp 1649977179
transform 1 0 59984 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_98_645
timestamp 1649977179
transform 1 0 60444 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_658
timestamp 1649977179
transform 1 0 61640 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_670
timestamp 1649977179
transform 1 0 62744 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_682
timestamp 1649977179
transform 1 0 63848 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_694
timestamp 1649977179
transform 1 0 64952 0 1 55488
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_98_701
timestamp 1649977179
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_713
timestamp 1649977179
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_725
timestamp 1649977179
transform 1 0 67804 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_737
timestamp 1649977179
transform 1 0 68908 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_749
timestamp 1649977179
transform 1 0 70012 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_755
timestamp 1649977179
transform 1 0 70564 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_757
timestamp 1649977179
transform 1 0 70748 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_769
timestamp 1649977179
transform 1 0 71852 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_781
timestamp 1649977179
transform 1 0 72956 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_793
timestamp 1649977179
transform 1 0 74060 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_805
timestamp 1649977179
transform 1 0 75164 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_811
timestamp 1649977179
transform 1 0 75716 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_813
timestamp 1649977179
transform 1 0 75900 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_98_825
timestamp 1649977179
transform 1 0 77004 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_831
timestamp 1649977179
transform 1 0 77556 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_838
timestamp 1649977179
transform 1 0 78200 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_7
timestamp 1649977179
transform 1 0 1748 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_13
timestamp 1649977179
transform 1 0 2300 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_25
timestamp 1649977179
transform 1 0 3404 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_37
timestamp 1649977179
transform 1 0 4508 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_49
timestamp 1649977179
transform 1 0 5612 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1649977179
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1649977179
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1649977179
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1649977179
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1649977179
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1649977179
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1649977179
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1649977179
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1649977179
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1649977179
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1649977179
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1649977179
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1649977179
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1649977179
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1649977179
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1649977179
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1649977179
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1649977179
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1649977179
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1649977179
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1649977179
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1649977179
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1649977179
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1649977179
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1649977179
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1649977179
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1649977179
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1649977179
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1649977179
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_605
timestamp 1649977179
transform 1 0 56764 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_619
timestamp 1649977179
transform 1 0 58052 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_625
timestamp 1649977179
transform 1 0 58604 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_635
timestamp 1649977179
transform 1 0 59524 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_649
timestamp 1649977179
transform 1 0 60812 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_663
timestamp 1649977179
transform 1 0 62100 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1649977179
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_673
timestamp 1649977179
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_685
timestamp 1649977179
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_697
timestamp 1649977179
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_709
timestamp 1649977179
transform 1 0 66332 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_721
timestamp 1649977179
transform 1 0 67436 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_727
timestamp 1649977179
transform 1 0 67988 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_729
timestamp 1649977179
transform 1 0 68172 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_741
timestamp 1649977179
transform 1 0 69276 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_753
timestamp 1649977179
transform 1 0 70380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_765
timestamp 1649977179
transform 1 0 71484 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_777
timestamp 1649977179
transform 1 0 72588 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_783
timestamp 1649977179
transform 1 0 73140 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_785
timestamp 1649977179
transform 1 0 73324 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_797
timestamp 1649977179
transform 1 0 74428 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_809
timestamp 1649977179
transform 1 0 75532 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_821
timestamp 1649977179
transform 1 0 76636 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_829
timestamp 1649977179
transform 1 0 77372 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_836
timestamp 1649977179
transform 1 0 78016 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_841
timestamp 1649977179
transform 1 0 78476 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_7
timestamp 1649977179
transform 1 0 1748 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_13
timestamp 1649977179
transform 1 0 2300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_25
timestamp 1649977179
transform 1 0 3404 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1649977179
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1649977179
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1649977179
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1649977179
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1649977179
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1649977179
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1649977179
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1649977179
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1649977179
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1649977179
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1649977179
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1649977179
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1649977179
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1649977179
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1649977179
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1649977179
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1649977179
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1649977179
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_625
timestamp 1649977179
transform 1 0 58604 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_628
timestamp 1649977179
transform 1 0 58880 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_640
timestamp 1649977179
transform 1 0 59984 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_655
timestamp 1649977179
transform 1 0 61364 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_669
timestamp 1649977179
transform 1 0 62652 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_675
timestamp 1649977179
transform 1 0 63204 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_687
timestamp 1649977179
transform 1 0 64308 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1649977179
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_701
timestamp 1649977179
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_713
timestamp 1649977179
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_725
timestamp 1649977179
transform 1 0 67804 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_737
timestamp 1649977179
transform 1 0 68908 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_749
timestamp 1649977179
transform 1 0 70012 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_755
timestamp 1649977179
transform 1 0 70564 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_757
timestamp 1649977179
transform 1 0 70748 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_769
timestamp 1649977179
transform 1 0 71852 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_781
timestamp 1649977179
transform 1 0 72956 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_793
timestamp 1649977179
transform 1 0 74060 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_805
timestamp 1649977179
transform 1 0 75164 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_811
timestamp 1649977179
transform 1 0 75716 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_813
timestamp 1649977179
transform 1 0 75900 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_825
timestamp 1649977179
transform 1 0 77004 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_831
timestamp 1649977179
transform 1 0 77556 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_838
timestamp 1649977179
transform 1 0 78200 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_7
timestamp 1649977179
transform 1 0 1748 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_19
timestamp 1649977179
transform 1 0 2852 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_31
timestamp 1649977179
transform 1 0 3956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_43
timestamp 1649977179
transform 1 0 5060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_55
timestamp 1649977179
transform 1 0 6164 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_69
timestamp 1649977179
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_81
timestamp 1649977179
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_93
timestamp 1649977179
transform 1 0 9660 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_105
timestamp 1649977179
transform 1 0 10764 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_111
timestamp 1649977179
transform 1 0 11316 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_113
timestamp 1649977179
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_125
timestamp 1649977179
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_137
timestamp 1649977179
transform 1 0 13708 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_149
timestamp 1649977179
transform 1 0 14812 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_161
timestamp 1649977179
transform 1 0 15916 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_167
timestamp 1649977179
transform 1 0 16468 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_169
timestamp 1649977179
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1649977179
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_193
timestamp 1649977179
transform 1 0 18860 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_205
timestamp 1649977179
transform 1 0 19964 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_217
timestamp 1649977179
transform 1 0 21068 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1649977179
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_237
timestamp 1649977179
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_249
timestamp 1649977179
transform 1 0 24012 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_261
timestamp 1649977179
transform 1 0 25116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1649977179
transform 1 0 26220 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1649977179
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_281
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_293
timestamp 1649977179
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_305
timestamp 1649977179
transform 1 0 29164 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_317
timestamp 1649977179
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_329
timestamp 1649977179
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1649977179
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_337
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_349
timestamp 1649977179
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_361
timestamp 1649977179
transform 1 0 34316 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_373
timestamp 1649977179
transform 1 0 35420 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_385
timestamp 1649977179
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_391
timestamp 1649977179
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_405
timestamp 1649977179
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_417
timestamp 1649977179
transform 1 0 39468 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_429
timestamp 1649977179
transform 1 0 40572 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_441
timestamp 1649977179
transform 1 0 41676 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_447
timestamp 1649977179
transform 1 0 42228 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_461
timestamp 1649977179
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_473
timestamp 1649977179
transform 1 0 44620 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_485
timestamp 1649977179
transform 1 0 45724 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_497
timestamp 1649977179
transform 1 0 46828 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1649977179
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_505
timestamp 1649977179
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_517
timestamp 1649977179
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_529
timestamp 1649977179
transform 1 0 49772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_541
timestamp 1649977179
transform 1 0 50876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_553
timestamp 1649977179
transform 1 0 51980 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1649977179
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_561
timestamp 1649977179
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1649977179
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_585
timestamp 1649977179
transform 1 0 54924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_597
timestamp 1649977179
transform 1 0 56028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_609
timestamp 1649977179
transform 1 0 57132 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1649977179
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_617
timestamp 1649977179
transform 1 0 57868 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_623
timestamp 1649977179
transform 1 0 58420 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_629
timestamp 1649977179
transform 1 0 58972 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_641
timestamp 1649977179
transform 1 0 60076 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_659
timestamp 1649977179
transform 1 0 61732 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_665
timestamp 1649977179
transform 1 0 62284 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_671
timestamp 1649977179
transform 1 0 62836 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_681
timestamp 1649977179
transform 1 0 63756 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_687
timestamp 1649977179
transform 1 0 64308 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_699
timestamp 1649977179
transform 1 0 65412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_711
timestamp 1649977179
transform 1 0 66516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_723
timestamp 1649977179
transform 1 0 67620 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_727
timestamp 1649977179
transform 1 0 67988 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_729
timestamp 1649977179
transform 1 0 68172 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_741
timestamp 1649977179
transform 1 0 69276 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_753
timestamp 1649977179
transform 1 0 70380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_765
timestamp 1649977179
transform 1 0 71484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_777
timestamp 1649977179
transform 1 0 72588 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_783
timestamp 1649977179
transform 1 0 73140 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_785
timestamp 1649977179
transform 1 0 73324 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_797
timestamp 1649977179
transform 1 0 74428 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_809
timestamp 1649977179
transform 1 0 75532 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_821
timestamp 1649977179
transform 1 0 76636 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_836
timestamp 1649977179
transform 1 0 78016 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_841
timestamp 1649977179
transform 1 0 78476 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_5
timestamp 1649977179
transform 1 0 1564 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_17
timestamp 1649977179
transform 1 0 2668 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_102_25
timestamp 1649977179
transform 1 0 3404 0 1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_102_29
timestamp 1649977179
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_41
timestamp 1649977179
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_53
timestamp 1649977179
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_65
timestamp 1649977179
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1649977179
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1649977179
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_85
timestamp 1649977179
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_97
timestamp 1649977179
transform 1 0 10028 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_109
timestamp 1649977179
transform 1 0 11132 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_121
timestamp 1649977179
transform 1 0 12236 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_133
timestamp 1649977179
transform 1 0 13340 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_139
timestamp 1649977179
transform 1 0 13892 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_141
timestamp 1649977179
transform 1 0 14076 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_153
timestamp 1649977179
transform 1 0 15180 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_165
timestamp 1649977179
transform 1 0 16284 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_177
timestamp 1649977179
transform 1 0 17388 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_189
timestamp 1649977179
transform 1 0 18492 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_195
timestamp 1649977179
transform 1 0 19044 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_197
timestamp 1649977179
transform 1 0 19228 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_209
timestamp 1649977179
transform 1 0 20332 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_221
timestamp 1649977179
transform 1 0 21436 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_233
timestamp 1649977179
transform 1 0 22540 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_245
timestamp 1649977179
transform 1 0 23644 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_251
timestamp 1649977179
transform 1 0 24196 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_253
timestamp 1649977179
transform 1 0 24380 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_265
timestamp 1649977179
transform 1 0 25484 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_277
timestamp 1649977179
transform 1 0 26588 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_289
timestamp 1649977179
transform 1 0 27692 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_301
timestamp 1649977179
transform 1 0 28796 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_307
timestamp 1649977179
transform 1 0 29348 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_309
timestamp 1649977179
transform 1 0 29532 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_321
timestamp 1649977179
transform 1 0 30636 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_333
timestamp 1649977179
transform 1 0 31740 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_345
timestamp 1649977179
transform 1 0 32844 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_357
timestamp 1649977179
transform 1 0 33948 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_363
timestamp 1649977179
transform 1 0 34500 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_365
timestamp 1649977179
transform 1 0 34684 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_377
timestamp 1649977179
transform 1 0 35788 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_389
timestamp 1649977179
transform 1 0 36892 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_401
timestamp 1649977179
transform 1 0 37996 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_413
timestamp 1649977179
transform 1 0 39100 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_419
timestamp 1649977179
transform 1 0 39652 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_421
timestamp 1649977179
transform 1 0 39836 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_433
timestamp 1649977179
transform 1 0 40940 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_445
timestamp 1649977179
transform 1 0 42044 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_457
timestamp 1649977179
transform 1 0 43148 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_469
timestamp 1649977179
transform 1 0 44252 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_475
timestamp 1649977179
transform 1 0 44804 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_477
timestamp 1649977179
transform 1 0 44988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_489
timestamp 1649977179
transform 1 0 46092 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_501
timestamp 1649977179
transform 1 0 47196 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_513
timestamp 1649977179
transform 1 0 48300 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_525
timestamp 1649977179
transform 1 0 49404 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_531
timestamp 1649977179
transform 1 0 49956 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_533
timestamp 1649977179
transform 1 0 50140 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_545
timestamp 1649977179
transform 1 0 51244 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_557
timestamp 1649977179
transform 1 0 52348 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_569
timestamp 1649977179
transform 1 0 53452 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_581
timestamp 1649977179
transform 1 0 54556 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_587
timestamp 1649977179
transform 1 0 55108 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_589
timestamp 1649977179
transform 1 0 55292 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_601
timestamp 1649977179
transform 1 0 56396 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_613
timestamp 1649977179
transform 1 0 57500 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_625
timestamp 1649977179
transform 1 0 58604 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_102_628
timestamp 1649977179
transform 1 0 58880 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_640
timestamp 1649977179
transform 1 0 59984 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_102_653
timestamp 1649977179
transform 1 0 61180 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_102_667
timestamp 1649977179
transform 1 0 62468 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_679
timestamp 1649977179
transform 1 0 63572 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_102_685
timestamp 1649977179
transform 1 0 64124 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_102_691
timestamp 1649977179
transform 1 0 64676 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_699
timestamp 1649977179
transform 1 0 65412 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_703
timestamp 1649977179
transform 1 0 65780 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_715
timestamp 1649977179
transform 1 0 66884 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_727
timestamp 1649977179
transform 1 0 67988 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_739
timestamp 1649977179
transform 1 0 69092 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_751
timestamp 1649977179
transform 1 0 70196 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_755
timestamp 1649977179
transform 1 0 70564 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_757
timestamp 1649977179
transform 1 0 70748 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_769
timestamp 1649977179
transform 1 0 71852 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_781
timestamp 1649977179
transform 1 0 72956 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_793
timestamp 1649977179
transform 1 0 74060 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_805
timestamp 1649977179
transform 1 0 75164 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_811
timestamp 1649977179
transform 1 0 75716 0 1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_813
timestamp 1649977179
transform 1 0 75900 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_102_825
timestamp 1649977179
transform 1 0 77004 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_102_833
timestamp 1649977179
transform 1 0 77740 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_102_838
timestamp 1649977179
transform 1 0 78200 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_7
timestamp 1649977179
transform 1 0 1748 0 -1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_103_13
timestamp 1649977179
transform 1 0 2300 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_25
timestamp 1649977179
transform 1 0 3404 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_37
timestamp 1649977179
transform 1 0 4508 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_49
timestamp 1649977179
transform 1 0 5612 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1649977179
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_57
timestamp 1649977179
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_69
timestamp 1649977179
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_81
timestamp 1649977179
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_93
timestamp 1649977179
transform 1 0 9660 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_105
timestamp 1649977179
transform 1 0 10764 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_111
timestamp 1649977179
transform 1 0 11316 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_113
timestamp 1649977179
transform 1 0 11500 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_125
timestamp 1649977179
transform 1 0 12604 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_137
timestamp 1649977179
transform 1 0 13708 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_149
timestamp 1649977179
transform 1 0 14812 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_161
timestamp 1649977179
transform 1 0 15916 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_167
timestamp 1649977179
transform 1 0 16468 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_169
timestamp 1649977179
transform 1 0 16652 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_181
timestamp 1649977179
transform 1 0 17756 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_193
timestamp 1649977179
transform 1 0 18860 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_205
timestamp 1649977179
transform 1 0 19964 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_217
timestamp 1649977179
transform 1 0 21068 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_223
timestamp 1649977179
transform 1 0 21620 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_225
timestamp 1649977179
transform 1 0 21804 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_237
timestamp 1649977179
transform 1 0 22908 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_249
timestamp 1649977179
transform 1 0 24012 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_261
timestamp 1649977179
transform 1 0 25116 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_273
timestamp 1649977179
transform 1 0 26220 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_279
timestamp 1649977179
transform 1 0 26772 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_281
timestamp 1649977179
transform 1 0 26956 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_293
timestamp 1649977179
transform 1 0 28060 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_305
timestamp 1649977179
transform 1 0 29164 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_317
timestamp 1649977179
transform 1 0 30268 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_329
timestamp 1649977179
transform 1 0 31372 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_335
timestamp 1649977179
transform 1 0 31924 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_337
timestamp 1649977179
transform 1 0 32108 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_349
timestamp 1649977179
transform 1 0 33212 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_361
timestamp 1649977179
transform 1 0 34316 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_373
timestamp 1649977179
transform 1 0 35420 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_385
timestamp 1649977179
transform 1 0 36524 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_391
timestamp 1649977179
transform 1 0 37076 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_393
timestamp 1649977179
transform 1 0 37260 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_405
timestamp 1649977179
transform 1 0 38364 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_417
timestamp 1649977179
transform 1 0 39468 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_429
timestamp 1649977179
transform 1 0 40572 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_441
timestamp 1649977179
transform 1 0 41676 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_447
timestamp 1649977179
transform 1 0 42228 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_449
timestamp 1649977179
transform 1 0 42412 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_461
timestamp 1649977179
transform 1 0 43516 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_473
timestamp 1649977179
transform 1 0 44620 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_485
timestamp 1649977179
transform 1 0 45724 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_497
timestamp 1649977179
transform 1 0 46828 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_503
timestamp 1649977179
transform 1 0 47380 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_505
timestamp 1649977179
transform 1 0 47564 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_517
timestamp 1649977179
transform 1 0 48668 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_529
timestamp 1649977179
transform 1 0 49772 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_541
timestamp 1649977179
transform 1 0 50876 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_553
timestamp 1649977179
transform 1 0 51980 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_559
timestamp 1649977179
transform 1 0 52532 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_561
timestamp 1649977179
transform 1 0 52716 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_573
timestamp 1649977179
transform 1 0 53820 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_585
timestamp 1649977179
transform 1 0 54924 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_597
timestamp 1649977179
transform 1 0 56028 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_609
timestamp 1649977179
transform 1 0 57132 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_615
timestamp 1649977179
transform 1 0 57684 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_617
timestamp 1649977179
transform 1 0 57868 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_103_629
timestamp 1649977179
transform 1 0 58972 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_633
timestamp 1649977179
transform 1 0 59340 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_103_636
timestamp 1649977179
transform 1 0 59616 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_648
timestamp 1649977179
transform 1 0 60720 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_103_654
timestamp 1649977179
transform 1 0 61272 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_103_668
timestamp 1649977179
transform 1 0 62560 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_675
timestamp 1649977179
transform 1 0 63204 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_681
timestamp 1649977179
transform 1 0 63756 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_695
timestamp 1649977179
transform 1 0 65044 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_701
timestamp 1649977179
transform 1 0 65596 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_707
timestamp 1649977179
transform 1 0 66148 0 -1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_103_713
timestamp 1649977179
transform 1 0 66700 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_725
timestamp 1649977179
transform 1 0 67804 0 -1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_103_729
timestamp 1649977179
transform 1 0 68172 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_741
timestamp 1649977179
transform 1 0 69276 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_753
timestamp 1649977179
transform 1 0 70380 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_765
timestamp 1649977179
transform 1 0 71484 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_777
timestamp 1649977179
transform 1 0 72588 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_783
timestamp 1649977179
transform 1 0 73140 0 -1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_785
timestamp 1649977179
transform 1 0 73324 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_797
timestamp 1649977179
transform 1 0 74428 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_809
timestamp 1649977179
transform 1 0 75532 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_821
timestamp 1649977179
transform 1 0 76636 0 -1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_103_829
timestamp 1649977179
transform 1 0 77372 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_103_836
timestamp 1649977179
transform 1 0 78016 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_841
timestamp 1649977179
transform 1 0 78476 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_7
timestamp 1649977179
transform 1 0 1748 0 1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_104_13
timestamp 1649977179
transform 1 0 2300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_104_25
timestamp 1649977179
transform 1 0 3404 0 1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_104_29
timestamp 1649977179
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_41
timestamp 1649977179
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_53
timestamp 1649977179
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_65
timestamp 1649977179
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1649977179
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1649977179
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_85
timestamp 1649977179
transform 1 0 8924 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_97
timestamp 1649977179
transform 1 0 10028 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_109
timestamp 1649977179
transform 1 0 11132 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_121
timestamp 1649977179
transform 1 0 12236 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_133
timestamp 1649977179
transform 1 0 13340 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_139
timestamp 1649977179
transform 1 0 13892 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_141
timestamp 1649977179
transform 1 0 14076 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_153
timestamp 1649977179
transform 1 0 15180 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_165
timestamp 1649977179
transform 1 0 16284 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_177
timestamp 1649977179
transform 1 0 17388 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_189
timestamp 1649977179
transform 1 0 18492 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_195
timestamp 1649977179
transform 1 0 19044 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_197
timestamp 1649977179
transform 1 0 19228 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_209
timestamp 1649977179
transform 1 0 20332 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_221
timestamp 1649977179
transform 1 0 21436 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_233
timestamp 1649977179
transform 1 0 22540 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_245
timestamp 1649977179
transform 1 0 23644 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_251
timestamp 1649977179
transform 1 0 24196 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_253
timestamp 1649977179
transform 1 0 24380 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_265
timestamp 1649977179
transform 1 0 25484 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_277
timestamp 1649977179
transform 1 0 26588 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_289
timestamp 1649977179
transform 1 0 27692 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_301
timestamp 1649977179
transform 1 0 28796 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_307
timestamp 1649977179
transform 1 0 29348 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_309
timestamp 1649977179
transform 1 0 29532 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_321
timestamp 1649977179
transform 1 0 30636 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_333
timestamp 1649977179
transform 1 0 31740 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_345
timestamp 1649977179
transform 1 0 32844 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_357
timestamp 1649977179
transform 1 0 33948 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_363
timestamp 1649977179
transform 1 0 34500 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_365
timestamp 1649977179
transform 1 0 34684 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_377
timestamp 1649977179
transform 1 0 35788 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_389
timestamp 1649977179
transform 1 0 36892 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_401
timestamp 1649977179
transform 1 0 37996 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_413
timestamp 1649977179
transform 1 0 39100 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_419
timestamp 1649977179
transform 1 0 39652 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_421
timestamp 1649977179
transform 1 0 39836 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_433
timestamp 1649977179
transform 1 0 40940 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_445
timestamp 1649977179
transform 1 0 42044 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_457
timestamp 1649977179
transform 1 0 43148 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_469
timestamp 1649977179
transform 1 0 44252 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_475
timestamp 1649977179
transform 1 0 44804 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_477
timestamp 1649977179
transform 1 0 44988 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_489
timestamp 1649977179
transform 1 0 46092 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_501
timestamp 1649977179
transform 1 0 47196 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_513
timestamp 1649977179
transform 1 0 48300 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_525
timestamp 1649977179
transform 1 0 49404 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_531
timestamp 1649977179
transform 1 0 49956 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_533
timestamp 1649977179
transform 1 0 50140 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_545
timestamp 1649977179
transform 1 0 51244 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_557
timestamp 1649977179
transform 1 0 52348 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_569
timestamp 1649977179
transform 1 0 53452 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_581
timestamp 1649977179
transform 1 0 54556 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_587
timestamp 1649977179
transform 1 0 55108 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_589
timestamp 1649977179
transform 1 0 55292 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_601
timestamp 1649977179
transform 1 0 56396 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_613
timestamp 1649977179
transform 1 0 57500 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_625
timestamp 1649977179
transform 1 0 58604 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_637
timestamp 1649977179
transform 1 0 59708 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_640
timestamp 1649977179
transform 1 0 59984 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_104_645
timestamp 1649977179
transform 1 0 60444 0 1 58752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_104_649
timestamp 1649977179
transform 1 0 60812 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_655
timestamp 1649977179
transform 1 0 61364 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_659
timestamp 1649977179
transform 1 0 61732 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_104_668
timestamp 1649977179
transform 1 0 62560 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_104_677
timestamp 1649977179
transform 1 0 63388 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_104_691
timestamp 1649977179
transform 1 0 64676 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_699
timestamp 1649977179
transform 1 0 65412 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_104_704
timestamp 1649977179
transform 1 0 65872 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_710
timestamp 1649977179
transform 1 0 66424 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_716
timestamp 1649977179
transform 1 0 66976 0 1 58752
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_104_722
timestamp 1649977179
transform 1 0 67528 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_734
timestamp 1649977179
transform 1 0 68632 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_746
timestamp 1649977179
transform 1 0 69736 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_104_754
timestamp 1649977179
transform 1 0 70472 0 1 58752
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_757
timestamp 1649977179
transform 1 0 70748 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_769
timestamp 1649977179
transform 1 0 71852 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_781
timestamp 1649977179
transform 1 0 72956 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_793
timestamp 1649977179
transform 1 0 74060 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_805
timestamp 1649977179
transform 1 0 75164 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_811
timestamp 1649977179
transform 1 0 75716 0 1 58752
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_813
timestamp 1649977179
transform 1 0 75900 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_104_825
timestamp 1649977179
transform 1 0 77004 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_831
timestamp 1649977179
transform 1 0 77556 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_104_838
timestamp 1649977179
transform 1 0 78200 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_7
timestamp 1649977179
transform 1 0 1748 0 -1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_105_13
timestamp 1649977179
transform 1 0 2300 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_25
timestamp 1649977179
transform 1 0 3404 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_37
timestamp 1649977179
transform 1 0 4508 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_49
timestamp 1649977179
transform 1 0 5612 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1649977179
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_57
timestamp 1649977179
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_69
timestamp 1649977179
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_81
timestamp 1649977179
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_93
timestamp 1649977179
transform 1 0 9660 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_105
timestamp 1649977179
transform 1 0 10764 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_111
timestamp 1649977179
transform 1 0 11316 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_113
timestamp 1649977179
transform 1 0 11500 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_125
timestamp 1649977179
transform 1 0 12604 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_137
timestamp 1649977179
transform 1 0 13708 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_149
timestamp 1649977179
transform 1 0 14812 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_161
timestamp 1649977179
transform 1 0 15916 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_167
timestamp 1649977179
transform 1 0 16468 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_169
timestamp 1649977179
transform 1 0 16652 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_181
timestamp 1649977179
transform 1 0 17756 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_193
timestamp 1649977179
transform 1 0 18860 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_205
timestamp 1649977179
transform 1 0 19964 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_217
timestamp 1649977179
transform 1 0 21068 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_223
timestamp 1649977179
transform 1 0 21620 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_225
timestamp 1649977179
transform 1 0 21804 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_237
timestamp 1649977179
transform 1 0 22908 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_249
timestamp 1649977179
transform 1 0 24012 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_261
timestamp 1649977179
transform 1 0 25116 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_273
timestamp 1649977179
transform 1 0 26220 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_279
timestamp 1649977179
transform 1 0 26772 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_281
timestamp 1649977179
transform 1 0 26956 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_293
timestamp 1649977179
transform 1 0 28060 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_305
timestamp 1649977179
transform 1 0 29164 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_317
timestamp 1649977179
transform 1 0 30268 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_329
timestamp 1649977179
transform 1 0 31372 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_335
timestamp 1649977179
transform 1 0 31924 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_337
timestamp 1649977179
transform 1 0 32108 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_349
timestamp 1649977179
transform 1 0 33212 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_361
timestamp 1649977179
transform 1 0 34316 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_373
timestamp 1649977179
transform 1 0 35420 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_385
timestamp 1649977179
transform 1 0 36524 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_391
timestamp 1649977179
transform 1 0 37076 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_393
timestamp 1649977179
transform 1 0 37260 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_405
timestamp 1649977179
transform 1 0 38364 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_417
timestamp 1649977179
transform 1 0 39468 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_429
timestamp 1649977179
transform 1 0 40572 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_441
timestamp 1649977179
transform 1 0 41676 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_447
timestamp 1649977179
transform 1 0 42228 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_449
timestamp 1649977179
transform 1 0 42412 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_461
timestamp 1649977179
transform 1 0 43516 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_473
timestamp 1649977179
transform 1 0 44620 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_485
timestamp 1649977179
transform 1 0 45724 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_497
timestamp 1649977179
transform 1 0 46828 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_503
timestamp 1649977179
transform 1 0 47380 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_505
timestamp 1649977179
transform 1 0 47564 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_517
timestamp 1649977179
transform 1 0 48668 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_529
timestamp 1649977179
transform 1 0 49772 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_541
timestamp 1649977179
transform 1 0 50876 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_553
timestamp 1649977179
transform 1 0 51980 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_559
timestamp 1649977179
transform 1 0 52532 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_561
timestamp 1649977179
transform 1 0 52716 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_573
timestamp 1649977179
transform 1 0 53820 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_585
timestamp 1649977179
transform 1 0 54924 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_597
timestamp 1649977179
transform 1 0 56028 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_609
timestamp 1649977179
transform 1 0 57132 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_615
timestamp 1649977179
transform 1 0 57684 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_617
timestamp 1649977179
transform 1 0 57868 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_629
timestamp 1649977179
transform 1 0 58972 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_641
timestamp 1649977179
transform 1 0 60076 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_653
timestamp 1649977179
transform 1 0 61180 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_657
timestamp 1649977179
transform 1 0 61548 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_105_660
timestamp 1649977179
transform 1 0 61824 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_105_668
timestamp 1649977179
transform 1 0 62560 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_105_673
timestamp 1649977179
transform 1 0 63020 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_684
timestamp 1649977179
transform 1 0 64032 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_696
timestamp 1649977179
transform 1 0 65136 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_708
timestamp 1649977179
transform 1 0 66240 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_714
timestamp 1649977179
transform 1 0 66792 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_105_720
timestamp 1649977179
transform 1 0 67344 0 -1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_105_729
timestamp 1649977179
transform 1 0 68172 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_741
timestamp 1649977179
transform 1 0 69276 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_753
timestamp 1649977179
transform 1 0 70380 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_765
timestamp 1649977179
transform 1 0 71484 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_777
timestamp 1649977179
transform 1 0 72588 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_105_783
timestamp 1649977179
transform 1 0 73140 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_785
timestamp 1649977179
transform 1 0 73324 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_797
timestamp 1649977179
transform 1 0 74428 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_809
timestamp 1649977179
transform 1 0 75532 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_105_821
timestamp 1649977179
transform 1 0 76636 0 -1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_105_829
timestamp 1649977179
transform 1 0 77372 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_836
timestamp 1649977179
transform 1 0 78016 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_841
timestamp 1649977179
transform 1 0 78476 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_7
timestamp 1649977179
transform 1 0 1748 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_19
timestamp 1649977179
transform 1 0 2852 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1649977179
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1649977179
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1649977179
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_53
timestamp 1649977179
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_65
timestamp 1649977179
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1649977179
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1649977179
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_85
timestamp 1649977179
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_97
timestamp 1649977179
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_109
timestamp 1649977179
transform 1 0 11132 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_121
timestamp 1649977179
transform 1 0 12236 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_133
timestamp 1649977179
transform 1 0 13340 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_139
timestamp 1649977179
transform 1 0 13892 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_141
timestamp 1649977179
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_153
timestamp 1649977179
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_165
timestamp 1649977179
transform 1 0 16284 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_177
timestamp 1649977179
transform 1 0 17388 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_189
timestamp 1649977179
transform 1 0 18492 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_195
timestamp 1649977179
transform 1 0 19044 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_197
timestamp 1649977179
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_209
timestamp 1649977179
transform 1 0 20332 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_221
timestamp 1649977179
transform 1 0 21436 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_233
timestamp 1649977179
transform 1 0 22540 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_245
timestamp 1649977179
transform 1 0 23644 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_251
timestamp 1649977179
transform 1 0 24196 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_253
timestamp 1649977179
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_265
timestamp 1649977179
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_277
timestamp 1649977179
transform 1 0 26588 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_289
timestamp 1649977179
transform 1 0 27692 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_301
timestamp 1649977179
transform 1 0 28796 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_307
timestamp 1649977179
transform 1 0 29348 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_309
timestamp 1649977179
transform 1 0 29532 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_321
timestamp 1649977179
transform 1 0 30636 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_333
timestamp 1649977179
transform 1 0 31740 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_345
timestamp 1649977179
transform 1 0 32844 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_357
timestamp 1649977179
transform 1 0 33948 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_363
timestamp 1649977179
transform 1 0 34500 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_365
timestamp 1649977179
transform 1 0 34684 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_377
timestamp 1649977179
transform 1 0 35788 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_389
timestamp 1649977179
transform 1 0 36892 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_401
timestamp 1649977179
transform 1 0 37996 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_413
timestamp 1649977179
transform 1 0 39100 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_419
timestamp 1649977179
transform 1 0 39652 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_421
timestamp 1649977179
transform 1 0 39836 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_433
timestamp 1649977179
transform 1 0 40940 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_445
timestamp 1649977179
transform 1 0 42044 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_457
timestamp 1649977179
transform 1 0 43148 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_469
timestamp 1649977179
transform 1 0 44252 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_475
timestamp 1649977179
transform 1 0 44804 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_477
timestamp 1649977179
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_489
timestamp 1649977179
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_501
timestamp 1649977179
transform 1 0 47196 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_513
timestamp 1649977179
transform 1 0 48300 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_525
timestamp 1649977179
transform 1 0 49404 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1649977179
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_533
timestamp 1649977179
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_545
timestamp 1649977179
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_557
timestamp 1649977179
transform 1 0 52348 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_569
timestamp 1649977179
transform 1 0 53452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_581
timestamp 1649977179
transform 1 0 54556 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_587
timestamp 1649977179
transform 1 0 55108 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_589
timestamp 1649977179
transform 1 0 55292 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_601
timestamp 1649977179
transform 1 0 56396 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_613
timestamp 1649977179
transform 1 0 57500 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_625
timestamp 1649977179
transform 1 0 58604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_637
timestamp 1649977179
transform 1 0 59708 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_643
timestamp 1649977179
transform 1 0 60260 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_645
timestamp 1649977179
transform 1 0 60444 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_657
timestamp 1649977179
transform 1 0 61548 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_661
timestamp 1649977179
transform 1 0 61916 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_664
timestamp 1649977179
transform 1 0 62192 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_670
timestamp 1649977179
transform 1 0 62744 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_678
timestamp 1649977179
transform 1 0 63480 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_684
timestamp 1649977179
transform 1 0 64032 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_696
timestamp 1649977179
transform 1 0 65136 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_709
timestamp 1649977179
transform 1 0 66332 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_718
timestamp 1649977179
transform 1 0 67160 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_724
timestamp 1649977179
transform 1 0 67712 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_730
timestamp 1649977179
transform 1 0 68264 0 1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_106_736
timestamp 1649977179
transform 1 0 68816 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_748
timestamp 1649977179
transform 1 0 69920 0 1 59840
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_106_757
timestamp 1649977179
transform 1 0 70748 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_769
timestamp 1649977179
transform 1 0 71852 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_781
timestamp 1649977179
transform 1 0 72956 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_793
timestamp 1649977179
transform 1 0 74060 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_805
timestamp 1649977179
transform 1 0 75164 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_811
timestamp 1649977179
transform 1 0 75716 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_813
timestamp 1649977179
transform 1 0 75900 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_825
timestamp 1649977179
transform 1 0 77004 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_831
timestamp 1649977179
transform 1 0 77556 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_106_838
timestamp 1649977179
transform 1 0 78200 0 1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_5
timestamp 1649977179
transform 1 0 1564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_17
timestamp 1649977179
transform 1 0 2668 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_29
timestamp 1649977179
transform 1 0 3772 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_41
timestamp 1649977179
transform 1 0 4876 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_53
timestamp 1649977179
transform 1 0 5980 0 -1 60928
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1649977179
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_69
timestamp 1649977179
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_81
timestamp 1649977179
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_93
timestamp 1649977179
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_105
timestamp 1649977179
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_111
timestamp 1649977179
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_113
timestamp 1649977179
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_125
timestamp 1649977179
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_137
timestamp 1649977179
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_149
timestamp 1649977179
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_161
timestamp 1649977179
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_167
timestamp 1649977179
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_169
timestamp 1649977179
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_181
timestamp 1649977179
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_193
timestamp 1649977179
transform 1 0 18860 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_205
timestamp 1649977179
transform 1 0 19964 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_217
timestamp 1649977179
transform 1 0 21068 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_223
timestamp 1649977179
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_225
timestamp 1649977179
transform 1 0 21804 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_237
timestamp 1649977179
transform 1 0 22908 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_249
timestamp 1649977179
transform 1 0 24012 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_261
timestamp 1649977179
transform 1 0 25116 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_273
timestamp 1649977179
transform 1 0 26220 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_279
timestamp 1649977179
transform 1 0 26772 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_281
timestamp 1649977179
transform 1 0 26956 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_293
timestamp 1649977179
transform 1 0 28060 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_305
timestamp 1649977179
transform 1 0 29164 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_317
timestamp 1649977179
transform 1 0 30268 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_329
timestamp 1649977179
transform 1 0 31372 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_335
timestamp 1649977179
transform 1 0 31924 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_337
timestamp 1649977179
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_349
timestamp 1649977179
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_361
timestamp 1649977179
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_373
timestamp 1649977179
transform 1 0 35420 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_385
timestamp 1649977179
transform 1 0 36524 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_391
timestamp 1649977179
transform 1 0 37076 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_393
timestamp 1649977179
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_405
timestamp 1649977179
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_417
timestamp 1649977179
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_429
timestamp 1649977179
transform 1 0 40572 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_441
timestamp 1649977179
transform 1 0 41676 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_447
timestamp 1649977179
transform 1 0 42228 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_449
timestamp 1649977179
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_461
timestamp 1649977179
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_473
timestamp 1649977179
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_485
timestamp 1649977179
transform 1 0 45724 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_497
timestamp 1649977179
transform 1 0 46828 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_503
timestamp 1649977179
transform 1 0 47380 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_505
timestamp 1649977179
transform 1 0 47564 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_517
timestamp 1649977179
transform 1 0 48668 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_529
timestamp 1649977179
transform 1 0 49772 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_541
timestamp 1649977179
transform 1 0 50876 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_553
timestamp 1649977179
transform 1 0 51980 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_559
timestamp 1649977179
transform 1 0 52532 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_561
timestamp 1649977179
transform 1 0 52716 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_573
timestamp 1649977179
transform 1 0 53820 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_585
timestamp 1649977179
transform 1 0 54924 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_597
timestamp 1649977179
transform 1 0 56028 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_609
timestamp 1649977179
transform 1 0 57132 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_615
timestamp 1649977179
transform 1 0 57684 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_617
timestamp 1649977179
transform 1 0 57868 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_629
timestamp 1649977179
transform 1 0 58972 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_641
timestamp 1649977179
transform 1 0 60076 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_653
timestamp 1649977179
transform 1 0 61180 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_107_665
timestamp 1649977179
transform 1 0 62284 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_107_668
timestamp 1649977179
transform 1 0 62560 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_675
timestamp 1649977179
transform 1 0 63204 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_684
timestamp 1649977179
transform 1 0 64032 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_696
timestamp 1649977179
transform 1 0 65136 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_107_705
timestamp 1649977179
transform 1 0 65964 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_107_719
timestamp 1649977179
transform 1 0 67252 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_107_727
timestamp 1649977179
transform 1 0 67988 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_729
timestamp 1649977179
transform 1 0 68172 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_741
timestamp 1649977179
transform 1 0 69276 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_753
timestamp 1649977179
transform 1 0 70380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_765
timestamp 1649977179
transform 1 0 71484 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_777
timestamp 1649977179
transform 1 0 72588 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_783
timestamp 1649977179
transform 1 0 73140 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_785
timestamp 1649977179
transform 1 0 73324 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_797
timestamp 1649977179
transform 1 0 74428 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_809
timestamp 1649977179
transform 1 0 75532 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_821
timestamp 1649977179
transform 1 0 76636 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_833
timestamp 1649977179
transform 1 0 77740 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_839
timestamp 1649977179
transform 1 0 78292 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_107_841
timestamp 1649977179
transform 1 0 78476 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_7
timestamp 1649977179
transform 1 0 1748 0 1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_108_13
timestamp 1649977179
transform 1 0 2300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_108_25
timestamp 1649977179
transform 1 0 3404 0 1 60928
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1649977179
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1649977179
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1649977179
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_65
timestamp 1649977179
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1649977179
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1649977179
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_85
timestamp 1649977179
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_97
timestamp 1649977179
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_109
timestamp 1649977179
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_121
timestamp 1649977179
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_133
timestamp 1649977179
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_139
timestamp 1649977179
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_141
timestamp 1649977179
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_153
timestamp 1649977179
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_165
timestamp 1649977179
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_177
timestamp 1649977179
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_189
timestamp 1649977179
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_195
timestamp 1649977179
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_197
timestamp 1649977179
transform 1 0 19228 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_209
timestamp 1649977179
transform 1 0 20332 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_221
timestamp 1649977179
transform 1 0 21436 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_233
timestamp 1649977179
transform 1 0 22540 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_245
timestamp 1649977179
transform 1 0 23644 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_251
timestamp 1649977179
transform 1 0 24196 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_253
timestamp 1649977179
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_265
timestamp 1649977179
transform 1 0 25484 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_277
timestamp 1649977179
transform 1 0 26588 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_289
timestamp 1649977179
transform 1 0 27692 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_301
timestamp 1649977179
transform 1 0 28796 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_307
timestamp 1649977179
transform 1 0 29348 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_309
timestamp 1649977179
transform 1 0 29532 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_321
timestamp 1649977179
transform 1 0 30636 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_333
timestamp 1649977179
transform 1 0 31740 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_345
timestamp 1649977179
transform 1 0 32844 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_357
timestamp 1649977179
transform 1 0 33948 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_363
timestamp 1649977179
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_365
timestamp 1649977179
transform 1 0 34684 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_377
timestamp 1649977179
transform 1 0 35788 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_389
timestamp 1649977179
transform 1 0 36892 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_401
timestamp 1649977179
transform 1 0 37996 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_413
timestamp 1649977179
transform 1 0 39100 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1649977179
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_421
timestamp 1649977179
transform 1 0 39836 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_433
timestamp 1649977179
transform 1 0 40940 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_445
timestamp 1649977179
transform 1 0 42044 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_457
timestamp 1649977179
transform 1 0 43148 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_469
timestamp 1649977179
transform 1 0 44252 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_475
timestamp 1649977179
transform 1 0 44804 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_477
timestamp 1649977179
transform 1 0 44988 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_489
timestamp 1649977179
transform 1 0 46092 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_501
timestamp 1649977179
transform 1 0 47196 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_513
timestamp 1649977179
transform 1 0 48300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_525
timestamp 1649977179
transform 1 0 49404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1649977179
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_533
timestamp 1649977179
transform 1 0 50140 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_545
timestamp 1649977179
transform 1 0 51244 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_557
timestamp 1649977179
transform 1 0 52348 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_569
timestamp 1649977179
transform 1 0 53452 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_581
timestamp 1649977179
transform 1 0 54556 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_587
timestamp 1649977179
transform 1 0 55108 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_589
timestamp 1649977179
transform 1 0 55292 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_601
timestamp 1649977179
transform 1 0 56396 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_613
timestamp 1649977179
transform 1 0 57500 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_625
timestamp 1649977179
transform 1 0 58604 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_637
timestamp 1649977179
transform 1 0 59708 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_643
timestamp 1649977179
transform 1 0 60260 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_645
timestamp 1649977179
transform 1 0 60444 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_657
timestamp 1649977179
transform 1 0 61548 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_669
timestamp 1649977179
transform 1 0 62652 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_673
timestamp 1649977179
transform 1 0 63020 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_676
timestamp 1649977179
transform 1 0 63296 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_684
timestamp 1649977179
transform 1 0 64032 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_696
timestamp 1649977179
transform 1 0 65136 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_709
timestamp 1649977179
transform 1 0 66332 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_716
timestamp 1649977179
transform 1 0 66976 0 1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_108_722
timestamp 1649977179
transform 1 0 67528 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_734
timestamp 1649977179
transform 1 0 68632 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_746
timestamp 1649977179
transform 1 0 69736 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_754
timestamp 1649977179
transform 1 0 70472 0 1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_108_757
timestamp 1649977179
transform 1 0 70748 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_769
timestamp 1649977179
transform 1 0 71852 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_781
timestamp 1649977179
transform 1 0 72956 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_793
timestamp 1649977179
transform 1 0 74060 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_805
timestamp 1649977179
transform 1 0 75164 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_811
timestamp 1649977179
transform 1 0 75716 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_813
timestamp 1649977179
transform 1 0 75900 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_108_825
timestamp 1649977179
transform 1 0 77004 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_831
timestamp 1649977179
transform 1 0 77556 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_108_838
timestamp 1649977179
transform 1 0 78200 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_7
timestamp 1649977179
transform 1 0 1748 0 -1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_109_13
timestamp 1649977179
transform 1 0 2300 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_25
timestamp 1649977179
transform 1 0 3404 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_37
timestamp 1649977179
transform 1 0 4508 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_49
timestamp 1649977179
transform 1 0 5612 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1649977179
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1649977179
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_69
timestamp 1649977179
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_81
timestamp 1649977179
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_93
timestamp 1649977179
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_105
timestamp 1649977179
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_111
timestamp 1649977179
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_113
timestamp 1649977179
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_125
timestamp 1649977179
transform 1 0 12604 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_137
timestamp 1649977179
transform 1 0 13708 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_149
timestamp 1649977179
transform 1 0 14812 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_161
timestamp 1649977179
transform 1 0 15916 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_167
timestamp 1649977179
transform 1 0 16468 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_169
timestamp 1649977179
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_181
timestamp 1649977179
transform 1 0 17756 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_193
timestamp 1649977179
transform 1 0 18860 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_205
timestamp 1649977179
transform 1 0 19964 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_217
timestamp 1649977179
transform 1 0 21068 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_223
timestamp 1649977179
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_225
timestamp 1649977179
transform 1 0 21804 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_237
timestamp 1649977179
transform 1 0 22908 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_249
timestamp 1649977179
transform 1 0 24012 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_261
timestamp 1649977179
transform 1 0 25116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_273
timestamp 1649977179
transform 1 0 26220 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_279
timestamp 1649977179
transform 1 0 26772 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_281
timestamp 1649977179
transform 1 0 26956 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_293
timestamp 1649977179
transform 1 0 28060 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_305
timestamp 1649977179
transform 1 0 29164 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_317
timestamp 1649977179
transform 1 0 30268 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_329
timestamp 1649977179
transform 1 0 31372 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_335
timestamp 1649977179
transform 1 0 31924 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_337
timestamp 1649977179
transform 1 0 32108 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_349
timestamp 1649977179
transform 1 0 33212 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_361
timestamp 1649977179
transform 1 0 34316 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_373
timestamp 1649977179
transform 1 0 35420 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_385
timestamp 1649977179
transform 1 0 36524 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_391
timestamp 1649977179
transform 1 0 37076 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_393
timestamp 1649977179
transform 1 0 37260 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_405
timestamp 1649977179
transform 1 0 38364 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_417
timestamp 1649977179
transform 1 0 39468 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_429
timestamp 1649977179
transform 1 0 40572 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_441
timestamp 1649977179
transform 1 0 41676 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_447
timestamp 1649977179
transform 1 0 42228 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_449
timestamp 1649977179
transform 1 0 42412 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_461
timestamp 1649977179
transform 1 0 43516 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_473
timestamp 1649977179
transform 1 0 44620 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_485
timestamp 1649977179
transform 1 0 45724 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_497
timestamp 1649977179
transform 1 0 46828 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_503
timestamp 1649977179
transform 1 0 47380 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_505
timestamp 1649977179
transform 1 0 47564 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_517
timestamp 1649977179
transform 1 0 48668 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_529
timestamp 1649977179
transform 1 0 49772 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_541
timestamp 1649977179
transform 1 0 50876 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_553
timestamp 1649977179
transform 1 0 51980 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_559
timestamp 1649977179
transform 1 0 52532 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_561
timestamp 1649977179
transform 1 0 52716 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_573
timestamp 1649977179
transform 1 0 53820 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_585
timestamp 1649977179
transform 1 0 54924 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_597
timestamp 1649977179
transform 1 0 56028 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_609
timestamp 1649977179
transform 1 0 57132 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_615
timestamp 1649977179
transform 1 0 57684 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_617
timestamp 1649977179
transform 1 0 57868 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_629
timestamp 1649977179
transform 1 0 58972 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_641
timestamp 1649977179
transform 1 0 60076 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_653
timestamp 1649977179
transform 1 0 61180 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_665
timestamp 1649977179
transform 1 0 62284 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_671
timestamp 1649977179
transform 1 0 62836 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_673
timestamp 1649977179
transform 1 0 63020 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_109_685
timestamp 1649977179
transform 1 0 64124 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_691
timestamp 1649977179
transform 1 0 64676 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_697
timestamp 1649977179
transform 1 0 65228 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_703
timestamp 1649977179
transform 1 0 65780 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_709
timestamp 1649977179
transform 1 0 66332 0 -1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_109_715
timestamp 1649977179
transform 1 0 66884 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_727
timestamp 1649977179
transform 1 0 67988 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_729
timestamp 1649977179
transform 1 0 68172 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_741
timestamp 1649977179
transform 1 0 69276 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_753
timestamp 1649977179
transform 1 0 70380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_765
timestamp 1649977179
transform 1 0 71484 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_777
timestamp 1649977179
transform 1 0 72588 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_783
timestamp 1649977179
transform 1 0 73140 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_785
timestamp 1649977179
transform 1 0 73324 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_797
timestamp 1649977179
transform 1 0 74428 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_809
timestamp 1649977179
transform 1 0 75532 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_821
timestamp 1649977179
transform 1 0 76636 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_109_829
timestamp 1649977179
transform 1 0 77372 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_109_836
timestamp 1649977179
transform 1 0 78016 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_841
timestamp 1649977179
transform 1 0 78476 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_7
timestamp 1649977179
transform 1 0 1748 0 1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_110_13
timestamp 1649977179
transform 1 0 2300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_110_25
timestamp 1649977179
transform 1 0 3404 0 1 62016
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1649977179
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_41
timestamp 1649977179
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_53
timestamp 1649977179
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_65
timestamp 1649977179
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1649977179
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1649977179
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_85
timestamp 1649977179
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_97
timestamp 1649977179
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_109
timestamp 1649977179
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_121
timestamp 1649977179
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_133
timestamp 1649977179
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_139
timestamp 1649977179
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_141
timestamp 1649977179
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_153
timestamp 1649977179
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_165
timestamp 1649977179
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_177
timestamp 1649977179
transform 1 0 17388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_189
timestamp 1649977179
transform 1 0 18492 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_195
timestamp 1649977179
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_197
timestamp 1649977179
transform 1 0 19228 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_209
timestamp 1649977179
transform 1 0 20332 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_221
timestamp 1649977179
transform 1 0 21436 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_233
timestamp 1649977179
transform 1 0 22540 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_245
timestamp 1649977179
transform 1 0 23644 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_251
timestamp 1649977179
transform 1 0 24196 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_253
timestamp 1649977179
transform 1 0 24380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_265
timestamp 1649977179
transform 1 0 25484 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_277
timestamp 1649977179
transform 1 0 26588 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_289
timestamp 1649977179
transform 1 0 27692 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_301
timestamp 1649977179
transform 1 0 28796 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_307
timestamp 1649977179
transform 1 0 29348 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_309
timestamp 1649977179
transform 1 0 29532 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_321
timestamp 1649977179
transform 1 0 30636 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_333
timestamp 1649977179
transform 1 0 31740 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_345
timestamp 1649977179
transform 1 0 32844 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_357
timestamp 1649977179
transform 1 0 33948 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_363
timestamp 1649977179
transform 1 0 34500 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_365
timestamp 1649977179
transform 1 0 34684 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_377
timestamp 1649977179
transform 1 0 35788 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_389
timestamp 1649977179
transform 1 0 36892 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_401
timestamp 1649977179
transform 1 0 37996 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_413
timestamp 1649977179
transform 1 0 39100 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_419
timestamp 1649977179
transform 1 0 39652 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_421
timestamp 1649977179
transform 1 0 39836 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_433
timestamp 1649977179
transform 1 0 40940 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_445
timestamp 1649977179
transform 1 0 42044 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_457
timestamp 1649977179
transform 1 0 43148 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_469
timestamp 1649977179
transform 1 0 44252 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_475
timestamp 1649977179
transform 1 0 44804 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_477
timestamp 1649977179
transform 1 0 44988 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_489
timestamp 1649977179
transform 1 0 46092 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_501
timestamp 1649977179
transform 1 0 47196 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_513
timestamp 1649977179
transform 1 0 48300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_525
timestamp 1649977179
transform 1 0 49404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_531
timestamp 1649977179
transform 1 0 49956 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_533
timestamp 1649977179
transform 1 0 50140 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_545
timestamp 1649977179
transform 1 0 51244 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_557
timestamp 1649977179
transform 1 0 52348 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_569
timestamp 1649977179
transform 1 0 53452 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_581
timestamp 1649977179
transform 1 0 54556 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_587
timestamp 1649977179
transform 1 0 55108 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_589
timestamp 1649977179
transform 1 0 55292 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_601
timestamp 1649977179
transform 1 0 56396 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_613
timestamp 1649977179
transform 1 0 57500 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_625
timestamp 1649977179
transform 1 0 58604 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_637
timestamp 1649977179
transform 1 0 59708 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_643
timestamp 1649977179
transform 1 0 60260 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_645
timestamp 1649977179
transform 1 0 60444 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_657
timestamp 1649977179
transform 1 0 61548 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_669
timestamp 1649977179
transform 1 0 62652 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_681
timestamp 1649977179
transform 1 0 63756 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_685
timestamp 1649977179
transform 1 0 64124 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_688
timestamp 1649977179
transform 1 0 64400 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_703
timestamp 1649977179
transform 1 0 65780 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_715
timestamp 1649977179
transform 1 0 66884 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_727
timestamp 1649977179
transform 1 0 67988 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_739
timestamp 1649977179
transform 1 0 69092 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_751
timestamp 1649977179
transform 1 0 70196 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_755
timestamp 1649977179
transform 1 0 70564 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_757
timestamp 1649977179
transform 1 0 70748 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_769
timestamp 1649977179
transform 1 0 71852 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_781
timestamp 1649977179
transform 1 0 72956 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_793
timestamp 1649977179
transform 1 0 74060 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_805
timestamp 1649977179
transform 1 0 75164 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_811
timestamp 1649977179
transform 1 0 75716 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_813
timestamp 1649977179
transform 1 0 75900 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_825
timestamp 1649977179
transform 1 0 77004 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_831
timestamp 1649977179
transform 1 0 77556 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_110_838
timestamp 1649977179
transform 1 0 78200 0 1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_111_7
timestamp 1649977179
transform 1 0 1748 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_19
timestamp 1649977179
transform 1 0 2852 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_31
timestamp 1649977179
transform 1 0 3956 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_43
timestamp 1649977179
transform 1 0 5060 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1649977179
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_57
timestamp 1649977179
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_69
timestamp 1649977179
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_81
timestamp 1649977179
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_93
timestamp 1649977179
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_105
timestamp 1649977179
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_111
timestamp 1649977179
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_113
timestamp 1649977179
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_125
timestamp 1649977179
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_137
timestamp 1649977179
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_149
timestamp 1649977179
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_161
timestamp 1649977179
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_167
timestamp 1649977179
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_169
timestamp 1649977179
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_181
timestamp 1649977179
transform 1 0 17756 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_193
timestamp 1649977179
transform 1 0 18860 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_205
timestamp 1649977179
transform 1 0 19964 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_217
timestamp 1649977179
transform 1 0 21068 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_223
timestamp 1649977179
transform 1 0 21620 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_225
timestamp 1649977179
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_237
timestamp 1649977179
transform 1 0 22908 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_249
timestamp 1649977179
transform 1 0 24012 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_261
timestamp 1649977179
transform 1 0 25116 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_273
timestamp 1649977179
transform 1 0 26220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_279
timestamp 1649977179
transform 1 0 26772 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_281
timestamp 1649977179
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_293
timestamp 1649977179
transform 1 0 28060 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_305
timestamp 1649977179
transform 1 0 29164 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_317
timestamp 1649977179
transform 1 0 30268 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_329
timestamp 1649977179
transform 1 0 31372 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_335
timestamp 1649977179
transform 1 0 31924 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_337
timestamp 1649977179
transform 1 0 32108 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_349
timestamp 1649977179
transform 1 0 33212 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_361
timestamp 1649977179
transform 1 0 34316 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_373
timestamp 1649977179
transform 1 0 35420 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_385
timestamp 1649977179
transform 1 0 36524 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_391
timestamp 1649977179
transform 1 0 37076 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_393
timestamp 1649977179
transform 1 0 37260 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_405
timestamp 1649977179
transform 1 0 38364 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_417
timestamp 1649977179
transform 1 0 39468 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_429
timestamp 1649977179
transform 1 0 40572 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_441
timestamp 1649977179
transform 1 0 41676 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_447
timestamp 1649977179
transform 1 0 42228 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_449
timestamp 1649977179
transform 1 0 42412 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_461
timestamp 1649977179
transform 1 0 43516 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_473
timestamp 1649977179
transform 1 0 44620 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_485
timestamp 1649977179
transform 1 0 45724 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_497
timestamp 1649977179
transform 1 0 46828 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_503
timestamp 1649977179
transform 1 0 47380 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_505
timestamp 1649977179
transform 1 0 47564 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_517
timestamp 1649977179
transform 1 0 48668 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_529
timestamp 1649977179
transform 1 0 49772 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_541
timestamp 1649977179
transform 1 0 50876 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_553
timestamp 1649977179
transform 1 0 51980 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_559
timestamp 1649977179
transform 1 0 52532 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_561
timestamp 1649977179
transform 1 0 52716 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_573
timestamp 1649977179
transform 1 0 53820 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_585
timestamp 1649977179
transform 1 0 54924 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_597
timestamp 1649977179
transform 1 0 56028 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_609
timestamp 1649977179
transform 1 0 57132 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_615
timestamp 1649977179
transform 1 0 57684 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_617
timestamp 1649977179
transform 1 0 57868 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_629
timestamp 1649977179
transform 1 0 58972 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_641
timestamp 1649977179
transform 1 0 60076 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_653
timestamp 1649977179
transform 1 0 61180 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_665
timestamp 1649977179
transform 1 0 62284 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_671
timestamp 1649977179
transform 1 0 62836 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_673
timestamp 1649977179
transform 1 0 63020 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_685
timestamp 1649977179
transform 1 0 64124 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_697
timestamp 1649977179
transform 1 0 65228 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_709
timestamp 1649977179
transform 1 0 66332 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_721
timestamp 1649977179
transform 1 0 67436 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_727
timestamp 1649977179
transform 1 0 67988 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_729
timestamp 1649977179
transform 1 0 68172 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_741
timestamp 1649977179
transform 1 0 69276 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_753
timestamp 1649977179
transform 1 0 70380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_765
timestamp 1649977179
transform 1 0 71484 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_777
timestamp 1649977179
transform 1 0 72588 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_783
timestamp 1649977179
transform 1 0 73140 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_785
timestamp 1649977179
transform 1 0 73324 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_797
timestamp 1649977179
transform 1 0 74428 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_809
timestamp 1649977179
transform 1 0 75532 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_821
timestamp 1649977179
transform 1 0 76636 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_836
timestamp 1649977179
transform 1 0 78016 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_841
timestamp 1649977179
transform 1 0 78476 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_5
timestamp 1649977179
transform 1 0 1564 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_17
timestamp 1649977179
transform 1 0 2668 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_112_25
timestamp 1649977179
transform 1 0 3404 0 1 63104
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1649977179
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1649977179
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_53
timestamp 1649977179
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_65
timestamp 1649977179
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1649977179
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1649977179
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_85
timestamp 1649977179
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_97
timestamp 1649977179
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_109
timestamp 1649977179
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_121
timestamp 1649977179
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_133
timestamp 1649977179
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_139
timestamp 1649977179
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_141
timestamp 1649977179
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_153
timestamp 1649977179
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_165
timestamp 1649977179
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_177
timestamp 1649977179
transform 1 0 17388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_189
timestamp 1649977179
transform 1 0 18492 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_195
timestamp 1649977179
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_197
timestamp 1649977179
transform 1 0 19228 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_209
timestamp 1649977179
transform 1 0 20332 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_221
timestamp 1649977179
transform 1 0 21436 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_233
timestamp 1649977179
transform 1 0 22540 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_245
timestamp 1649977179
transform 1 0 23644 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_251
timestamp 1649977179
transform 1 0 24196 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_253
timestamp 1649977179
transform 1 0 24380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_265
timestamp 1649977179
transform 1 0 25484 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_277
timestamp 1649977179
transform 1 0 26588 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_289
timestamp 1649977179
transform 1 0 27692 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_301
timestamp 1649977179
transform 1 0 28796 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_307
timestamp 1649977179
transform 1 0 29348 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_309
timestamp 1649977179
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_321
timestamp 1649977179
transform 1 0 30636 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_333
timestamp 1649977179
transform 1 0 31740 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_345
timestamp 1649977179
transform 1 0 32844 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_357
timestamp 1649977179
transform 1 0 33948 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_363
timestamp 1649977179
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_365
timestamp 1649977179
transform 1 0 34684 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_377
timestamp 1649977179
transform 1 0 35788 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_389
timestamp 1649977179
transform 1 0 36892 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_401
timestamp 1649977179
transform 1 0 37996 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_413
timestamp 1649977179
transform 1 0 39100 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_419
timestamp 1649977179
transform 1 0 39652 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_421
timestamp 1649977179
transform 1 0 39836 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_433
timestamp 1649977179
transform 1 0 40940 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_445
timestamp 1649977179
transform 1 0 42044 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_457
timestamp 1649977179
transform 1 0 43148 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_469
timestamp 1649977179
transform 1 0 44252 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_475
timestamp 1649977179
transform 1 0 44804 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_477
timestamp 1649977179
transform 1 0 44988 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_489
timestamp 1649977179
transform 1 0 46092 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_501
timestamp 1649977179
transform 1 0 47196 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_513
timestamp 1649977179
transform 1 0 48300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_525
timestamp 1649977179
transform 1 0 49404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_531
timestamp 1649977179
transform 1 0 49956 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_533
timestamp 1649977179
transform 1 0 50140 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_545
timestamp 1649977179
transform 1 0 51244 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_557
timestamp 1649977179
transform 1 0 52348 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_569
timestamp 1649977179
transform 1 0 53452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_581
timestamp 1649977179
transform 1 0 54556 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_587
timestamp 1649977179
transform 1 0 55108 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_589
timestamp 1649977179
transform 1 0 55292 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_601
timestamp 1649977179
transform 1 0 56396 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_613
timestamp 1649977179
transform 1 0 57500 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_625
timestamp 1649977179
transform 1 0 58604 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_637
timestamp 1649977179
transform 1 0 59708 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_643
timestamp 1649977179
transform 1 0 60260 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_645
timestamp 1649977179
transform 1 0 60444 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_657
timestamp 1649977179
transform 1 0 61548 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_669
timestamp 1649977179
transform 1 0 62652 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_681
timestamp 1649977179
transform 1 0 63756 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_693
timestamp 1649977179
transform 1 0 64860 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_699
timestamp 1649977179
transform 1 0 65412 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_701
timestamp 1649977179
transform 1 0 65596 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_713
timestamp 1649977179
transform 1 0 66700 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_725
timestamp 1649977179
transform 1 0 67804 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_737
timestamp 1649977179
transform 1 0 68908 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_749
timestamp 1649977179
transform 1 0 70012 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_755
timestamp 1649977179
transform 1 0 70564 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_757
timestamp 1649977179
transform 1 0 70748 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_769
timestamp 1649977179
transform 1 0 71852 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_781
timestamp 1649977179
transform 1 0 72956 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_793
timestamp 1649977179
transform 1 0 74060 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_805
timestamp 1649977179
transform 1 0 75164 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_811
timestamp 1649977179
transform 1 0 75716 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_813
timestamp 1649977179
transform 1 0 75900 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_825
timestamp 1649977179
transform 1 0 77004 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_112_833
timestamp 1649977179
transform 1 0 77740 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_112_838
timestamp 1649977179
transform 1 0 78200 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_7
timestamp 1649977179
transform 1 0 1748 0 -1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_113_13
timestamp 1649977179
transform 1 0 2300 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_25
timestamp 1649977179
transform 1 0 3404 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_37
timestamp 1649977179
transform 1 0 4508 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_49
timestamp 1649977179
transform 1 0 5612 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1649977179
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1649977179
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_69
timestamp 1649977179
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_81
timestamp 1649977179
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_93
timestamp 1649977179
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_105
timestamp 1649977179
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_111
timestamp 1649977179
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_113
timestamp 1649977179
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_125
timestamp 1649977179
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_137
timestamp 1649977179
transform 1 0 13708 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_149
timestamp 1649977179
transform 1 0 14812 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_161
timestamp 1649977179
transform 1 0 15916 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_167
timestamp 1649977179
transform 1 0 16468 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_169
timestamp 1649977179
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_181
timestamp 1649977179
transform 1 0 17756 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_193
timestamp 1649977179
transform 1 0 18860 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_205
timestamp 1649977179
transform 1 0 19964 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_217
timestamp 1649977179
transform 1 0 21068 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_223
timestamp 1649977179
transform 1 0 21620 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_225
timestamp 1649977179
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_237
timestamp 1649977179
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_249
timestamp 1649977179
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_261
timestamp 1649977179
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_273
timestamp 1649977179
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_279
timestamp 1649977179
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_281
timestamp 1649977179
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_293
timestamp 1649977179
transform 1 0 28060 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_305
timestamp 1649977179
transform 1 0 29164 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_317
timestamp 1649977179
transform 1 0 30268 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_329
timestamp 1649977179
transform 1 0 31372 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_335
timestamp 1649977179
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_337
timestamp 1649977179
transform 1 0 32108 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_349
timestamp 1649977179
transform 1 0 33212 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_361
timestamp 1649977179
transform 1 0 34316 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_373
timestamp 1649977179
transform 1 0 35420 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_385
timestamp 1649977179
transform 1 0 36524 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_391
timestamp 1649977179
transform 1 0 37076 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_393
timestamp 1649977179
transform 1 0 37260 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_405
timestamp 1649977179
transform 1 0 38364 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_417
timestamp 1649977179
transform 1 0 39468 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_429
timestamp 1649977179
transform 1 0 40572 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_441
timestamp 1649977179
transform 1 0 41676 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_447
timestamp 1649977179
transform 1 0 42228 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_449
timestamp 1649977179
transform 1 0 42412 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_461
timestamp 1649977179
transform 1 0 43516 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_473
timestamp 1649977179
transform 1 0 44620 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_485
timestamp 1649977179
transform 1 0 45724 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_497
timestamp 1649977179
transform 1 0 46828 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_503
timestamp 1649977179
transform 1 0 47380 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_505
timestamp 1649977179
transform 1 0 47564 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_517
timestamp 1649977179
transform 1 0 48668 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_529
timestamp 1649977179
transform 1 0 49772 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_541
timestamp 1649977179
transform 1 0 50876 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_553
timestamp 1649977179
transform 1 0 51980 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_559
timestamp 1649977179
transform 1 0 52532 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_561
timestamp 1649977179
transform 1 0 52716 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_573
timestamp 1649977179
transform 1 0 53820 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_585
timestamp 1649977179
transform 1 0 54924 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_597
timestamp 1649977179
transform 1 0 56028 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_609
timestamp 1649977179
transform 1 0 57132 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_615
timestamp 1649977179
transform 1 0 57684 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_617
timestamp 1649977179
transform 1 0 57868 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_629
timestamp 1649977179
transform 1 0 58972 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_641
timestamp 1649977179
transform 1 0 60076 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_653
timestamp 1649977179
transform 1 0 61180 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_665
timestamp 1649977179
transform 1 0 62284 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_671
timestamp 1649977179
transform 1 0 62836 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_673
timestamp 1649977179
transform 1 0 63020 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_685
timestamp 1649977179
transform 1 0 64124 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_697
timestamp 1649977179
transform 1 0 65228 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_709
timestamp 1649977179
transform 1 0 66332 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_721
timestamp 1649977179
transform 1 0 67436 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_727
timestamp 1649977179
transform 1 0 67988 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_729
timestamp 1649977179
transform 1 0 68172 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_741
timestamp 1649977179
transform 1 0 69276 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_753
timestamp 1649977179
transform 1 0 70380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_765
timestamp 1649977179
transform 1 0 71484 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_777
timestamp 1649977179
transform 1 0 72588 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_783
timestamp 1649977179
transform 1 0 73140 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_785
timestamp 1649977179
transform 1 0 73324 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_797
timestamp 1649977179
transform 1 0 74428 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_809
timestamp 1649977179
transform 1 0 75532 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_821
timestamp 1649977179
transform 1 0 76636 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_113_829
timestamp 1649977179
transform 1 0 77372 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_836
timestamp 1649977179
transform 1 0 78016 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_841
timestamp 1649977179
transform 1 0 78476 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_114_7
timestamp 1649977179
transform 1 0 1748 0 1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_114_13
timestamp 1649977179
transform 1 0 2300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_114_25
timestamp 1649977179
transform 1 0 3404 0 1 64192
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1649977179
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1649977179
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_53
timestamp 1649977179
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_65
timestamp 1649977179
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1649977179
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1649977179
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_85
timestamp 1649977179
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_97
timestamp 1649977179
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_109
timestamp 1649977179
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_121
timestamp 1649977179
transform 1 0 12236 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_133
timestamp 1649977179
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_139
timestamp 1649977179
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_141
timestamp 1649977179
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_153
timestamp 1649977179
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_165
timestamp 1649977179
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_177
timestamp 1649977179
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_189
timestamp 1649977179
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_195
timestamp 1649977179
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_197
timestamp 1649977179
transform 1 0 19228 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_209
timestamp 1649977179
transform 1 0 20332 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_221
timestamp 1649977179
transform 1 0 21436 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_233
timestamp 1649977179
transform 1 0 22540 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_245
timestamp 1649977179
transform 1 0 23644 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_251
timestamp 1649977179
transform 1 0 24196 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_253
timestamp 1649977179
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_265
timestamp 1649977179
transform 1 0 25484 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_277
timestamp 1649977179
transform 1 0 26588 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_289
timestamp 1649977179
transform 1 0 27692 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_301
timestamp 1649977179
transform 1 0 28796 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_307
timestamp 1649977179
transform 1 0 29348 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_309
timestamp 1649977179
transform 1 0 29532 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_321
timestamp 1649977179
transform 1 0 30636 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_333
timestamp 1649977179
transform 1 0 31740 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_345
timestamp 1649977179
transform 1 0 32844 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_357
timestamp 1649977179
transform 1 0 33948 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_363
timestamp 1649977179
transform 1 0 34500 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_365
timestamp 1649977179
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_377
timestamp 1649977179
transform 1 0 35788 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_389
timestamp 1649977179
transform 1 0 36892 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_401
timestamp 1649977179
transform 1 0 37996 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_413
timestamp 1649977179
transform 1 0 39100 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_419
timestamp 1649977179
transform 1 0 39652 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_421
timestamp 1649977179
transform 1 0 39836 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_433
timestamp 1649977179
transform 1 0 40940 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_445
timestamp 1649977179
transform 1 0 42044 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_457
timestamp 1649977179
transform 1 0 43148 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_469
timestamp 1649977179
transform 1 0 44252 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_475
timestamp 1649977179
transform 1 0 44804 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_477
timestamp 1649977179
transform 1 0 44988 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_489
timestamp 1649977179
transform 1 0 46092 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_501
timestamp 1649977179
transform 1 0 47196 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_513
timestamp 1649977179
transform 1 0 48300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_525
timestamp 1649977179
transform 1 0 49404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_531
timestamp 1649977179
transform 1 0 49956 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_533
timestamp 1649977179
transform 1 0 50140 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_545
timestamp 1649977179
transform 1 0 51244 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_557
timestamp 1649977179
transform 1 0 52348 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_569
timestamp 1649977179
transform 1 0 53452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_581
timestamp 1649977179
transform 1 0 54556 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_587
timestamp 1649977179
transform 1 0 55108 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_589
timestamp 1649977179
transform 1 0 55292 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_601
timestamp 1649977179
transform 1 0 56396 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_613
timestamp 1649977179
transform 1 0 57500 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_625
timestamp 1649977179
transform 1 0 58604 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_637
timestamp 1649977179
transform 1 0 59708 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_643
timestamp 1649977179
transform 1 0 60260 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_645
timestamp 1649977179
transform 1 0 60444 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_657
timestamp 1649977179
transform 1 0 61548 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_669
timestamp 1649977179
transform 1 0 62652 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_681
timestamp 1649977179
transform 1 0 63756 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_693
timestamp 1649977179
transform 1 0 64860 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_699
timestamp 1649977179
transform 1 0 65412 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_701
timestamp 1649977179
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_713
timestamp 1649977179
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_725
timestamp 1649977179
transform 1 0 67804 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_737
timestamp 1649977179
transform 1 0 68908 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_749
timestamp 1649977179
transform 1 0 70012 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_755
timestamp 1649977179
transform 1 0 70564 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_757
timestamp 1649977179
transform 1 0 70748 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_769
timestamp 1649977179
transform 1 0 71852 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_781
timestamp 1649977179
transform 1 0 72956 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_793
timestamp 1649977179
transform 1 0 74060 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_805
timestamp 1649977179
transform 1 0 75164 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_811
timestamp 1649977179
transform 1 0 75716 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_813
timestamp 1649977179
transform 1 0 75900 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_114_825
timestamp 1649977179
transform 1 0 77004 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_831
timestamp 1649977179
transform 1 0 77556 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_838
timestamp 1649977179
transform 1 0 78200 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_7
timestamp 1649977179
transform 1 0 1748 0 -1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_115_13
timestamp 1649977179
transform 1 0 2300 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_25
timestamp 1649977179
transform 1 0 3404 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_37
timestamp 1649977179
transform 1 0 4508 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_49
timestamp 1649977179
transform 1 0 5612 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1649977179
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_57
timestamp 1649977179
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_69
timestamp 1649977179
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_81
timestamp 1649977179
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_93
timestamp 1649977179
transform 1 0 9660 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_105
timestamp 1649977179
transform 1 0 10764 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_111
timestamp 1649977179
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_113
timestamp 1649977179
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_125
timestamp 1649977179
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_137
timestamp 1649977179
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_149
timestamp 1649977179
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_161
timestamp 1649977179
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_167
timestamp 1649977179
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_169
timestamp 1649977179
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_181
timestamp 1649977179
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_193
timestamp 1649977179
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_205
timestamp 1649977179
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_217
timestamp 1649977179
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_223
timestamp 1649977179
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_225
timestamp 1649977179
transform 1 0 21804 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_237
timestamp 1649977179
transform 1 0 22908 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_249
timestamp 1649977179
transform 1 0 24012 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_261
timestamp 1649977179
transform 1 0 25116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_273
timestamp 1649977179
transform 1 0 26220 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_279
timestamp 1649977179
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_281
timestamp 1649977179
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_293
timestamp 1649977179
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_305
timestamp 1649977179
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_317
timestamp 1649977179
transform 1 0 30268 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_329
timestamp 1649977179
transform 1 0 31372 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_335
timestamp 1649977179
transform 1 0 31924 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_337
timestamp 1649977179
transform 1 0 32108 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_349
timestamp 1649977179
transform 1 0 33212 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_361
timestamp 1649977179
transform 1 0 34316 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_373
timestamp 1649977179
transform 1 0 35420 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_385
timestamp 1649977179
transform 1 0 36524 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_391
timestamp 1649977179
transform 1 0 37076 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_393
timestamp 1649977179
transform 1 0 37260 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_405
timestamp 1649977179
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_417
timestamp 1649977179
transform 1 0 39468 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_429
timestamp 1649977179
transform 1 0 40572 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_441
timestamp 1649977179
transform 1 0 41676 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_447
timestamp 1649977179
transform 1 0 42228 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_449
timestamp 1649977179
transform 1 0 42412 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_461
timestamp 1649977179
transform 1 0 43516 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_473
timestamp 1649977179
transform 1 0 44620 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_485
timestamp 1649977179
transform 1 0 45724 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_497
timestamp 1649977179
transform 1 0 46828 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_503
timestamp 1649977179
transform 1 0 47380 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_505
timestamp 1649977179
transform 1 0 47564 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_517
timestamp 1649977179
transform 1 0 48668 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_529
timestamp 1649977179
transform 1 0 49772 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_541
timestamp 1649977179
transform 1 0 50876 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_553
timestamp 1649977179
transform 1 0 51980 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_559
timestamp 1649977179
transform 1 0 52532 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_561
timestamp 1649977179
transform 1 0 52716 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_573
timestamp 1649977179
transform 1 0 53820 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_585
timestamp 1649977179
transform 1 0 54924 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_597
timestamp 1649977179
transform 1 0 56028 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_609
timestamp 1649977179
transform 1 0 57132 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_615
timestamp 1649977179
transform 1 0 57684 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_617
timestamp 1649977179
transform 1 0 57868 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_629
timestamp 1649977179
transform 1 0 58972 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_641
timestamp 1649977179
transform 1 0 60076 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_653
timestamp 1649977179
transform 1 0 61180 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_665
timestamp 1649977179
transform 1 0 62284 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_671
timestamp 1649977179
transform 1 0 62836 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_673
timestamp 1649977179
transform 1 0 63020 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_685
timestamp 1649977179
transform 1 0 64124 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_697
timestamp 1649977179
transform 1 0 65228 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_709
timestamp 1649977179
transform 1 0 66332 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_721
timestamp 1649977179
transform 1 0 67436 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_727
timestamp 1649977179
transform 1 0 67988 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_729
timestamp 1649977179
transform 1 0 68172 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_741
timestamp 1649977179
transform 1 0 69276 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_753
timestamp 1649977179
transform 1 0 70380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_765
timestamp 1649977179
transform 1 0 71484 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_777
timestamp 1649977179
transform 1 0 72588 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_783
timestamp 1649977179
transform 1 0 73140 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_785
timestamp 1649977179
transform 1 0 73324 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_797
timestamp 1649977179
transform 1 0 74428 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_809
timestamp 1649977179
transform 1 0 75532 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_821
timestamp 1649977179
transform 1 0 76636 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_115_829
timestamp 1649977179
transform 1 0 77372 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_115_836
timestamp 1649977179
transform 1 0 78016 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_841
timestamp 1649977179
transform 1 0 78476 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_7
timestamp 1649977179
transform 1 0 1748 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_19
timestamp 1649977179
transform 1 0 2852 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1649977179
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1649977179
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_41
timestamp 1649977179
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_53
timestamp 1649977179
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_65
timestamp 1649977179
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1649977179
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1649977179
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_85
timestamp 1649977179
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_97
timestamp 1649977179
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_109
timestamp 1649977179
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_121
timestamp 1649977179
transform 1 0 12236 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_133
timestamp 1649977179
transform 1 0 13340 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_139
timestamp 1649977179
transform 1 0 13892 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_141
timestamp 1649977179
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_153
timestamp 1649977179
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_165
timestamp 1649977179
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_177
timestamp 1649977179
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_189
timestamp 1649977179
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_195
timestamp 1649977179
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_197
timestamp 1649977179
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_209
timestamp 1649977179
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_221
timestamp 1649977179
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_233
timestamp 1649977179
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_245
timestamp 1649977179
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_251
timestamp 1649977179
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_253
timestamp 1649977179
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_265
timestamp 1649977179
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_277
timestamp 1649977179
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_289
timestamp 1649977179
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_301
timestamp 1649977179
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_307
timestamp 1649977179
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_309
timestamp 1649977179
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_321
timestamp 1649977179
transform 1 0 30636 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_333
timestamp 1649977179
transform 1 0 31740 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_345
timestamp 1649977179
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_357
timestamp 1649977179
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_363
timestamp 1649977179
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_365
timestamp 1649977179
transform 1 0 34684 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_377
timestamp 1649977179
transform 1 0 35788 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_389
timestamp 1649977179
transform 1 0 36892 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_401
timestamp 1649977179
transform 1 0 37996 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_413
timestamp 1649977179
transform 1 0 39100 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_419
timestamp 1649977179
transform 1 0 39652 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_421
timestamp 1649977179
transform 1 0 39836 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_433
timestamp 1649977179
transform 1 0 40940 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_445
timestamp 1649977179
transform 1 0 42044 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_457
timestamp 1649977179
transform 1 0 43148 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_469
timestamp 1649977179
transform 1 0 44252 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_475
timestamp 1649977179
transform 1 0 44804 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_477
timestamp 1649977179
transform 1 0 44988 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_489
timestamp 1649977179
transform 1 0 46092 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_501
timestamp 1649977179
transform 1 0 47196 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_513
timestamp 1649977179
transform 1 0 48300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_525
timestamp 1649977179
transform 1 0 49404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_531
timestamp 1649977179
transform 1 0 49956 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_533
timestamp 1649977179
transform 1 0 50140 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_545
timestamp 1649977179
transform 1 0 51244 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_557
timestamp 1649977179
transform 1 0 52348 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_569
timestamp 1649977179
transform 1 0 53452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_581
timestamp 1649977179
transform 1 0 54556 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_587
timestamp 1649977179
transform 1 0 55108 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_589
timestamp 1649977179
transform 1 0 55292 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_601
timestamp 1649977179
transform 1 0 56396 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_613
timestamp 1649977179
transform 1 0 57500 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_625
timestamp 1649977179
transform 1 0 58604 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_637
timestamp 1649977179
transform 1 0 59708 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_643
timestamp 1649977179
transform 1 0 60260 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_645
timestamp 1649977179
transform 1 0 60444 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_657
timestamp 1649977179
transform 1 0 61548 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_669
timestamp 1649977179
transform 1 0 62652 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_681
timestamp 1649977179
transform 1 0 63756 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_693
timestamp 1649977179
transform 1 0 64860 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_699
timestamp 1649977179
transform 1 0 65412 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_701
timestamp 1649977179
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_713
timestamp 1649977179
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_725
timestamp 1649977179
transform 1 0 67804 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_737
timestamp 1649977179
transform 1 0 68908 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_749
timestamp 1649977179
transform 1 0 70012 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_755
timestamp 1649977179
transform 1 0 70564 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_757
timestamp 1649977179
transform 1 0 70748 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_769
timestamp 1649977179
transform 1 0 71852 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_781
timestamp 1649977179
transform 1 0 72956 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_793
timestamp 1649977179
transform 1 0 74060 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_805
timestamp 1649977179
transform 1 0 75164 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_811
timestamp 1649977179
transform 1 0 75716 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_813
timestamp 1649977179
transform 1 0 75900 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_116_825
timestamp 1649977179
transform 1 0 77004 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_831
timestamp 1649977179
transform 1 0 77556 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_838
timestamp 1649977179
transform 1 0 78200 0 1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_117_5
timestamp 1649977179
transform 1 0 1564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_17
timestamp 1649977179
transform 1 0 2668 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_29
timestamp 1649977179
transform 1 0 3772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_41
timestamp 1649977179
transform 1 0 4876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_53
timestamp 1649977179
transform 1 0 5980 0 -1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1649977179
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_69
timestamp 1649977179
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_81
timestamp 1649977179
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_93
timestamp 1649977179
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_105
timestamp 1649977179
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_111
timestamp 1649977179
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_113
timestamp 1649977179
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_125
timestamp 1649977179
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_137
timestamp 1649977179
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_149
timestamp 1649977179
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_161
timestamp 1649977179
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_167
timestamp 1649977179
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_169
timestamp 1649977179
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_181
timestamp 1649977179
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_193
timestamp 1649977179
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_205
timestamp 1649977179
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_217
timestamp 1649977179
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_223
timestamp 1649977179
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_225
timestamp 1649977179
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_237
timestamp 1649977179
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_249
timestamp 1649977179
transform 1 0 24012 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_261
timestamp 1649977179
transform 1 0 25116 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_273
timestamp 1649977179
transform 1 0 26220 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_279
timestamp 1649977179
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_281
timestamp 1649977179
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_293
timestamp 1649977179
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_305
timestamp 1649977179
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_317
timestamp 1649977179
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_329
timestamp 1649977179
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_335
timestamp 1649977179
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_337
timestamp 1649977179
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_349
timestamp 1649977179
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_361
timestamp 1649977179
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_373
timestamp 1649977179
transform 1 0 35420 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_385
timestamp 1649977179
transform 1 0 36524 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_391
timestamp 1649977179
transform 1 0 37076 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_393
timestamp 1649977179
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_405
timestamp 1649977179
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_417
timestamp 1649977179
transform 1 0 39468 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_429
timestamp 1649977179
transform 1 0 40572 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_441
timestamp 1649977179
transform 1 0 41676 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_447
timestamp 1649977179
transform 1 0 42228 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_449
timestamp 1649977179
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_461
timestamp 1649977179
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_473
timestamp 1649977179
transform 1 0 44620 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_485
timestamp 1649977179
transform 1 0 45724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_497
timestamp 1649977179
transform 1 0 46828 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_503
timestamp 1649977179
transform 1 0 47380 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_505
timestamp 1649977179
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_517
timestamp 1649977179
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_529
timestamp 1649977179
transform 1 0 49772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_541
timestamp 1649977179
transform 1 0 50876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_553
timestamp 1649977179
transform 1 0 51980 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_559
timestamp 1649977179
transform 1 0 52532 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_561
timestamp 1649977179
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_573
timestamp 1649977179
transform 1 0 53820 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_585
timestamp 1649977179
transform 1 0 54924 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_597
timestamp 1649977179
transform 1 0 56028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_609
timestamp 1649977179
transform 1 0 57132 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_615
timestamp 1649977179
transform 1 0 57684 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_617
timestamp 1649977179
transform 1 0 57868 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_629
timestamp 1649977179
transform 1 0 58972 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_641
timestamp 1649977179
transform 1 0 60076 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_653
timestamp 1649977179
transform 1 0 61180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_665
timestamp 1649977179
transform 1 0 62284 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_671
timestamp 1649977179
transform 1 0 62836 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_673
timestamp 1649977179
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_685
timestamp 1649977179
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_697
timestamp 1649977179
transform 1 0 65228 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_709
timestamp 1649977179
transform 1 0 66332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_721
timestamp 1649977179
transform 1 0 67436 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_727
timestamp 1649977179
transform 1 0 67988 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_729
timestamp 1649977179
transform 1 0 68172 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_741
timestamp 1649977179
transform 1 0 69276 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_753
timestamp 1649977179
transform 1 0 70380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_765
timestamp 1649977179
transform 1 0 71484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_777
timestamp 1649977179
transform 1 0 72588 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_783
timestamp 1649977179
transform 1 0 73140 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_785
timestamp 1649977179
transform 1 0 73324 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_797
timestamp 1649977179
transform 1 0 74428 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_809
timestamp 1649977179
transform 1 0 75532 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_821
timestamp 1649977179
transform 1 0 76636 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_833
timestamp 1649977179
transform 1 0 77740 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_839
timestamp 1649977179
transform 1 0 78292 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_117_841
timestamp 1649977179
transform 1 0 78476 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_7
timestamp 1649977179
transform 1 0 1748 0 1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_118_13
timestamp 1649977179
transform 1 0 2300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_118_25
timestamp 1649977179
transform 1 0 3404 0 1 66368
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1649977179
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1649977179
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1649977179
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_65
timestamp 1649977179
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1649977179
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1649977179
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_85
timestamp 1649977179
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_97
timestamp 1649977179
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_109
timestamp 1649977179
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_121
timestamp 1649977179
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1649977179
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1649977179
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_141
timestamp 1649977179
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_153
timestamp 1649977179
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_165
timestamp 1649977179
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_177
timestamp 1649977179
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1649977179
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1649977179
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_197
timestamp 1649977179
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_209
timestamp 1649977179
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_221
timestamp 1649977179
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_233
timestamp 1649977179
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1649977179
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1649977179
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_253
timestamp 1649977179
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_265
timestamp 1649977179
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_277
timestamp 1649977179
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_289
timestamp 1649977179
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1649977179
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1649977179
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_309
timestamp 1649977179
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_321
timestamp 1649977179
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_333
timestamp 1649977179
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_345
timestamp 1649977179
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1649977179
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1649977179
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_365
timestamp 1649977179
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_377
timestamp 1649977179
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_389
timestamp 1649977179
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_401
timestamp 1649977179
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1649977179
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1649977179
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_421
timestamp 1649977179
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_433
timestamp 1649977179
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_445
timestamp 1649977179
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_457
timestamp 1649977179
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1649977179
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1649977179
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_477
timestamp 1649977179
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_489
timestamp 1649977179
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_501
timestamp 1649977179
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_513
timestamp 1649977179
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1649977179
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1649977179
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_533
timestamp 1649977179
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_545
timestamp 1649977179
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_557
timestamp 1649977179
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_569
timestamp 1649977179
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1649977179
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1649977179
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_589
timestamp 1649977179
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_601
timestamp 1649977179
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_613
timestamp 1649977179
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_625
timestamp 1649977179
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1649977179
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1649977179
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_645
timestamp 1649977179
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_657
timestamp 1649977179
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_669
timestamp 1649977179
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_681
timestamp 1649977179
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1649977179
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1649977179
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_701
timestamp 1649977179
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_713
timestamp 1649977179
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_725
timestamp 1649977179
transform 1 0 67804 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_737
timestamp 1649977179
transform 1 0 68908 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_749
timestamp 1649977179
transform 1 0 70012 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_755
timestamp 1649977179
transform 1 0 70564 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_757
timestamp 1649977179
transform 1 0 70748 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_769
timestamp 1649977179
transform 1 0 71852 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_781
timestamp 1649977179
transform 1 0 72956 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_793
timestamp 1649977179
transform 1 0 74060 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_805
timestamp 1649977179
transform 1 0 75164 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_811
timestamp 1649977179
transform 1 0 75716 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_813
timestamp 1649977179
transform 1 0 75900 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_118_825
timestamp 1649977179
transform 1 0 77004 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_831
timestamp 1649977179
transform 1 0 77556 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_838
timestamp 1649977179
transform 1 0 78200 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_7
timestamp 1649977179
transform 1 0 1748 0 -1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_119_13
timestamp 1649977179
transform 1 0 2300 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_25
timestamp 1649977179
transform 1 0 3404 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_37
timestamp 1649977179
transform 1 0 4508 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_49
timestamp 1649977179
transform 1 0 5612 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1649977179
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1649977179
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_69
timestamp 1649977179
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_81
timestamp 1649977179
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_93
timestamp 1649977179
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1649977179
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1649977179
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_113
timestamp 1649977179
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_125
timestamp 1649977179
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_137
timestamp 1649977179
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_149
timestamp 1649977179
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1649977179
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1649977179
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_169
timestamp 1649977179
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_181
timestamp 1649977179
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_193
timestamp 1649977179
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_205
timestamp 1649977179
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1649977179
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1649977179
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_225
timestamp 1649977179
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_237
timestamp 1649977179
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_249
timestamp 1649977179
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_261
timestamp 1649977179
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1649977179
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1649977179
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_281
timestamp 1649977179
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_293
timestamp 1649977179
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_305
timestamp 1649977179
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_317
timestamp 1649977179
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1649977179
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1649977179
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_337
timestamp 1649977179
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_349
timestamp 1649977179
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_361
timestamp 1649977179
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_373
timestamp 1649977179
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1649977179
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1649977179
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_393
timestamp 1649977179
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_405
timestamp 1649977179
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_417
timestamp 1649977179
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_429
timestamp 1649977179
transform 1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1649977179
transform 1 0 41676 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1649977179
transform 1 0 42228 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_449
timestamp 1649977179
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_461
timestamp 1649977179
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_473
timestamp 1649977179
transform 1 0 44620 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_485
timestamp 1649977179
transform 1 0 45724 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_497
timestamp 1649977179
transform 1 0 46828 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1649977179
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_505
timestamp 1649977179
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_517
timestamp 1649977179
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_529
timestamp 1649977179
transform 1 0 49772 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_541
timestamp 1649977179
transform 1 0 50876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_553
timestamp 1649977179
transform 1 0 51980 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1649977179
transform 1 0 52532 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_561
timestamp 1649977179
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_573
timestamp 1649977179
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_585
timestamp 1649977179
transform 1 0 54924 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_597
timestamp 1649977179
transform 1 0 56028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1649977179
transform 1 0 57132 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1649977179
transform 1 0 57684 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_617
timestamp 1649977179
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_629
timestamp 1649977179
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_641
timestamp 1649977179
transform 1 0 60076 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_653
timestamp 1649977179
transform 1 0 61180 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_665
timestamp 1649977179
transform 1 0 62284 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_671
timestamp 1649977179
transform 1 0 62836 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_673
timestamp 1649977179
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_685
timestamp 1649977179
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_697
timestamp 1649977179
transform 1 0 65228 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_709
timestamp 1649977179
transform 1 0 66332 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_721
timestamp 1649977179
transform 1 0 67436 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_727
timestamp 1649977179
transform 1 0 67988 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_729
timestamp 1649977179
transform 1 0 68172 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_741
timestamp 1649977179
transform 1 0 69276 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_753
timestamp 1649977179
transform 1 0 70380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_765
timestamp 1649977179
transform 1 0 71484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_777
timestamp 1649977179
transform 1 0 72588 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_783
timestamp 1649977179
transform 1 0 73140 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_785
timestamp 1649977179
transform 1 0 73324 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_797
timestamp 1649977179
transform 1 0 74428 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_809
timestamp 1649977179
transform 1 0 75532 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_821
timestamp 1649977179
transform 1 0 76636 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_119_829
timestamp 1649977179
transform 1 0 77372 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_836
timestamp 1649977179
transform 1 0 78016 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_841
timestamp 1649977179
transform 1 0 78476 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_7
timestamp 1649977179
transform 1 0 1748 0 1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_120_13
timestamp 1649977179
transform 1 0 2300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_25
timestamp 1649977179
transform 1 0 3404 0 1 67456
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1649977179
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1649977179
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_53
timestamp 1649977179
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_65
timestamp 1649977179
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1649977179
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1649977179
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_85
timestamp 1649977179
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_97
timestamp 1649977179
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_109
timestamp 1649977179
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_121
timestamp 1649977179
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1649977179
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1649977179
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_141
timestamp 1649977179
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_153
timestamp 1649977179
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_165
timestamp 1649977179
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_177
timestamp 1649977179
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1649977179
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1649977179
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_197
timestamp 1649977179
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_209
timestamp 1649977179
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_221
timestamp 1649977179
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_233
timestamp 1649977179
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1649977179
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1649977179
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_253
timestamp 1649977179
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_265
timestamp 1649977179
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_277
timestamp 1649977179
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_289
timestamp 1649977179
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1649977179
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1649977179
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_309
timestamp 1649977179
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_321
timestamp 1649977179
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_333
timestamp 1649977179
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_345
timestamp 1649977179
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1649977179
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1649977179
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_365
timestamp 1649977179
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_377
timestamp 1649977179
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_389
timestamp 1649977179
transform 1 0 36892 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_401
timestamp 1649977179
transform 1 0 37996 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_413
timestamp 1649977179
transform 1 0 39100 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_419
timestamp 1649977179
transform 1 0 39652 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_421
timestamp 1649977179
transform 1 0 39836 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_433
timestamp 1649977179
transform 1 0 40940 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_445
timestamp 1649977179
transform 1 0 42044 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_457
timestamp 1649977179
transform 1 0 43148 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_469
timestamp 1649977179
transform 1 0 44252 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_475
timestamp 1649977179
transform 1 0 44804 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_477
timestamp 1649977179
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_489
timestamp 1649977179
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_501
timestamp 1649977179
transform 1 0 47196 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_513
timestamp 1649977179
transform 1 0 48300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1649977179
transform 1 0 49404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1649977179
transform 1 0 49956 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_533
timestamp 1649977179
transform 1 0 50140 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_545
timestamp 1649977179
transform 1 0 51244 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_557
timestamp 1649977179
transform 1 0 52348 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_569
timestamp 1649977179
transform 1 0 53452 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_581
timestamp 1649977179
transform 1 0 54556 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_587
timestamp 1649977179
transform 1 0 55108 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_589
timestamp 1649977179
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_601
timestamp 1649977179
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_613
timestamp 1649977179
transform 1 0 57500 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_625
timestamp 1649977179
transform 1 0 58604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1649977179
transform 1 0 59708 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1649977179
transform 1 0 60260 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_645
timestamp 1649977179
transform 1 0 60444 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_657
timestamp 1649977179
transform 1 0 61548 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_669
timestamp 1649977179
transform 1 0 62652 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_681
timestamp 1649977179
transform 1 0 63756 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_693
timestamp 1649977179
transform 1 0 64860 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1649977179
transform 1 0 65412 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_701
timestamp 1649977179
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_713
timestamp 1649977179
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_725
timestamp 1649977179
transform 1 0 67804 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_737
timestamp 1649977179
transform 1 0 68908 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_749
timestamp 1649977179
transform 1 0 70012 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_755
timestamp 1649977179
transform 1 0 70564 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_757
timestamp 1649977179
transform 1 0 70748 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_769
timestamp 1649977179
transform 1 0 71852 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_781
timestamp 1649977179
transform 1 0 72956 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_793
timestamp 1649977179
transform 1 0 74060 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_805
timestamp 1649977179
transform 1 0 75164 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_811
timestamp 1649977179
transform 1 0 75716 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_813
timestamp 1649977179
transform 1 0 75900 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_120_825
timestamp 1649977179
transform 1 0 77004 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_120_831
timestamp 1649977179
transform 1 0 77556 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_120_838
timestamp 1649977179
transform 1 0 78200 0 1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_121_7
timestamp 1649977179
transform 1 0 1748 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_19
timestamp 1649977179
transform 1 0 2852 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_31
timestamp 1649977179
transform 1 0 3956 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_43
timestamp 1649977179
transform 1 0 5060 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1649977179
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1649977179
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_69
timestamp 1649977179
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_81
timestamp 1649977179
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_93
timestamp 1649977179
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1649977179
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1649977179
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_113
timestamp 1649977179
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_125
timestamp 1649977179
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_137
timestamp 1649977179
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_149
timestamp 1649977179
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1649977179
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1649977179
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_169
timestamp 1649977179
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_181
timestamp 1649977179
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_193
timestamp 1649977179
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_205
timestamp 1649977179
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1649977179
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1649977179
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_225
timestamp 1649977179
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_237
timestamp 1649977179
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_249
timestamp 1649977179
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_261
timestamp 1649977179
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1649977179
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1649977179
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_281
timestamp 1649977179
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_293
timestamp 1649977179
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_305
timestamp 1649977179
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_317
timestamp 1649977179
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_329
timestamp 1649977179
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_335
timestamp 1649977179
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_337
timestamp 1649977179
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_349
timestamp 1649977179
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_361
timestamp 1649977179
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_373
timestamp 1649977179
transform 1 0 35420 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_385
timestamp 1649977179
transform 1 0 36524 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1649977179
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_393
timestamp 1649977179
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_405
timestamp 1649977179
transform 1 0 38364 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_417
timestamp 1649977179
transform 1 0 39468 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_429
timestamp 1649977179
transform 1 0 40572 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_441
timestamp 1649977179
transform 1 0 41676 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_447
timestamp 1649977179
transform 1 0 42228 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_449
timestamp 1649977179
transform 1 0 42412 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_461
timestamp 1649977179
transform 1 0 43516 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_473
timestamp 1649977179
transform 1 0 44620 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_485
timestamp 1649977179
transform 1 0 45724 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_497
timestamp 1649977179
transform 1 0 46828 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_503
timestamp 1649977179
transform 1 0 47380 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_505
timestamp 1649977179
transform 1 0 47564 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_517
timestamp 1649977179
transform 1 0 48668 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_529
timestamp 1649977179
transform 1 0 49772 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_541
timestamp 1649977179
transform 1 0 50876 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_553
timestamp 1649977179
transform 1 0 51980 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_559
timestamp 1649977179
transform 1 0 52532 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_561
timestamp 1649977179
transform 1 0 52716 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_573
timestamp 1649977179
transform 1 0 53820 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_585
timestamp 1649977179
transform 1 0 54924 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_597
timestamp 1649977179
transform 1 0 56028 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_609
timestamp 1649977179
transform 1 0 57132 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_615
timestamp 1649977179
transform 1 0 57684 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_617
timestamp 1649977179
transform 1 0 57868 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_629
timestamp 1649977179
transform 1 0 58972 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_641
timestamp 1649977179
transform 1 0 60076 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_653
timestamp 1649977179
transform 1 0 61180 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_665
timestamp 1649977179
transform 1 0 62284 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_671
timestamp 1649977179
transform 1 0 62836 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_673
timestamp 1649977179
transform 1 0 63020 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_685
timestamp 1649977179
transform 1 0 64124 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_697
timestamp 1649977179
transform 1 0 65228 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_709
timestamp 1649977179
transform 1 0 66332 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1649977179
transform 1 0 67436 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1649977179
transform 1 0 67988 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_729
timestamp 1649977179
transform 1 0 68172 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_741
timestamp 1649977179
transform 1 0 69276 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_753
timestamp 1649977179
transform 1 0 70380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_765
timestamp 1649977179
transform 1 0 71484 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_777
timestamp 1649977179
transform 1 0 72588 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_783
timestamp 1649977179
transform 1 0 73140 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_785
timestamp 1649977179
transform 1 0 73324 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_797
timestamp 1649977179
transform 1 0 74428 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_809
timestamp 1649977179
transform 1 0 75532 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_821
timestamp 1649977179
transform 1 0 76636 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_836
timestamp 1649977179
transform 1 0 78016 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_841
timestamp 1649977179
transform 1 0 78476 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_5
timestamp 1649977179
transform 1 0 1564 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_17
timestamp 1649977179
transform 1 0 2668 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_25
timestamp 1649977179
transform 1 0 3404 0 1 68544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1649977179
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1649977179
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1649977179
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_65
timestamp 1649977179
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1649977179
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1649977179
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_85
timestamp 1649977179
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_97
timestamp 1649977179
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_109
timestamp 1649977179
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_121
timestamp 1649977179
transform 1 0 12236 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_133
timestamp 1649977179
transform 1 0 13340 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_139
timestamp 1649977179
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_141
timestamp 1649977179
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_153
timestamp 1649977179
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_165
timestamp 1649977179
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_177
timestamp 1649977179
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_189
timestamp 1649977179
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1649977179
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_197
timestamp 1649977179
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_209
timestamp 1649977179
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_221
timestamp 1649977179
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_233
timestamp 1649977179
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1649977179
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1649977179
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_253
timestamp 1649977179
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_265
timestamp 1649977179
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_277
timestamp 1649977179
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_289
timestamp 1649977179
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_301
timestamp 1649977179
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1649977179
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_309
timestamp 1649977179
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_321
timestamp 1649977179
transform 1 0 30636 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_333
timestamp 1649977179
transform 1 0 31740 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_345
timestamp 1649977179
transform 1 0 32844 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_357
timestamp 1649977179
transform 1 0 33948 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_363
timestamp 1649977179
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_365
timestamp 1649977179
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_377
timestamp 1649977179
transform 1 0 35788 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_389
timestamp 1649977179
transform 1 0 36892 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_401
timestamp 1649977179
transform 1 0 37996 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_413
timestamp 1649977179
transform 1 0 39100 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_419
timestamp 1649977179
transform 1 0 39652 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_421
timestamp 1649977179
transform 1 0 39836 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_433
timestamp 1649977179
transform 1 0 40940 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_445
timestamp 1649977179
transform 1 0 42044 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_457
timestamp 1649977179
transform 1 0 43148 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_469
timestamp 1649977179
transform 1 0 44252 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_475
timestamp 1649977179
transform 1 0 44804 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_477
timestamp 1649977179
transform 1 0 44988 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_489
timestamp 1649977179
transform 1 0 46092 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_501
timestamp 1649977179
transform 1 0 47196 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_513
timestamp 1649977179
transform 1 0 48300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_525
timestamp 1649977179
transform 1 0 49404 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_531
timestamp 1649977179
transform 1 0 49956 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_533
timestamp 1649977179
transform 1 0 50140 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_545
timestamp 1649977179
transform 1 0 51244 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_557
timestamp 1649977179
transform 1 0 52348 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_569
timestamp 1649977179
transform 1 0 53452 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_581
timestamp 1649977179
transform 1 0 54556 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_587
timestamp 1649977179
transform 1 0 55108 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_589
timestamp 1649977179
transform 1 0 55292 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_601
timestamp 1649977179
transform 1 0 56396 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_613
timestamp 1649977179
transform 1 0 57500 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_625
timestamp 1649977179
transform 1 0 58604 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_637
timestamp 1649977179
transform 1 0 59708 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_643
timestamp 1649977179
transform 1 0 60260 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_645
timestamp 1649977179
transform 1 0 60444 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_657
timestamp 1649977179
transform 1 0 61548 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_669
timestamp 1649977179
transform 1 0 62652 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_681
timestamp 1649977179
transform 1 0 63756 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_693
timestamp 1649977179
transform 1 0 64860 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_699
timestamp 1649977179
transform 1 0 65412 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_701
timestamp 1649977179
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_713
timestamp 1649977179
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_725
timestamp 1649977179
transform 1 0 67804 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_737
timestamp 1649977179
transform 1 0 68908 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_122_745
timestamp 1649977179
transform 1 0 69644 0 1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_122_751
timestamp 1649977179
transform 1 0 70196 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_122_755
timestamp 1649977179
transform 1 0 70564 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_759
timestamp 1649977179
transform 1 0 70932 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_771
timestamp 1649977179
transform 1 0 72036 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_786
timestamp 1649977179
transform 1 0 73416 0 1 68544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_122_792
timestamp 1649977179
transform 1 0 73968 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_804
timestamp 1649977179
transform 1 0 75072 0 1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_122_813
timestamp 1649977179
transform 1 0 75900 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_825
timestamp 1649977179
transform 1 0 77004 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_122_833
timestamp 1649977179
transform 1 0 77740 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_838
timestamp 1649977179
transform 1 0 78200 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_7
timestamp 1649977179
transform 1 0 1748 0 -1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_123_13
timestamp 1649977179
transform 1 0 2300 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_25
timestamp 1649977179
transform 1 0 3404 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_37
timestamp 1649977179
transform 1 0 4508 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_49
timestamp 1649977179
transform 1 0 5612 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1649977179
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1649977179
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_69
timestamp 1649977179
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_81
timestamp 1649977179
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_93
timestamp 1649977179
transform 1 0 9660 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_105
timestamp 1649977179
transform 1 0 10764 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_111
timestamp 1649977179
transform 1 0 11316 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_113
timestamp 1649977179
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_125
timestamp 1649977179
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_137
timestamp 1649977179
transform 1 0 13708 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_149
timestamp 1649977179
transform 1 0 14812 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_161
timestamp 1649977179
transform 1 0 15916 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1649977179
transform 1 0 16468 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_169
timestamp 1649977179
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_181
timestamp 1649977179
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_193
timestamp 1649977179
transform 1 0 18860 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_205
timestamp 1649977179
transform 1 0 19964 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_217
timestamp 1649977179
transform 1 0 21068 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_223
timestamp 1649977179
transform 1 0 21620 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_225
timestamp 1649977179
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_237
timestamp 1649977179
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_249
timestamp 1649977179
transform 1 0 24012 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_261
timestamp 1649977179
transform 1 0 25116 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_273
timestamp 1649977179
transform 1 0 26220 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_279
timestamp 1649977179
transform 1 0 26772 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_281
timestamp 1649977179
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_293
timestamp 1649977179
transform 1 0 28060 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_305
timestamp 1649977179
transform 1 0 29164 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_317
timestamp 1649977179
transform 1 0 30268 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_329
timestamp 1649977179
transform 1 0 31372 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_335
timestamp 1649977179
transform 1 0 31924 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_337
timestamp 1649977179
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_349
timestamp 1649977179
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_361
timestamp 1649977179
transform 1 0 34316 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_373
timestamp 1649977179
transform 1 0 35420 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_385
timestamp 1649977179
transform 1 0 36524 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_391
timestamp 1649977179
transform 1 0 37076 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_393
timestamp 1649977179
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_405
timestamp 1649977179
transform 1 0 38364 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_417
timestamp 1649977179
transform 1 0 39468 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_429
timestamp 1649977179
transform 1 0 40572 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_441
timestamp 1649977179
transform 1 0 41676 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_447
timestamp 1649977179
transform 1 0 42228 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_449
timestamp 1649977179
transform 1 0 42412 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_461
timestamp 1649977179
transform 1 0 43516 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_473
timestamp 1649977179
transform 1 0 44620 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_485
timestamp 1649977179
transform 1 0 45724 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_497
timestamp 1649977179
transform 1 0 46828 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_503
timestamp 1649977179
transform 1 0 47380 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_505
timestamp 1649977179
transform 1 0 47564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_517
timestamp 1649977179
transform 1 0 48668 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_529
timestamp 1649977179
transform 1 0 49772 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_541
timestamp 1649977179
transform 1 0 50876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_553
timestamp 1649977179
transform 1 0 51980 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_559
timestamp 1649977179
transform 1 0 52532 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_561
timestamp 1649977179
transform 1 0 52716 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_573
timestamp 1649977179
transform 1 0 53820 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_585
timestamp 1649977179
transform 1 0 54924 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_597
timestamp 1649977179
transform 1 0 56028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_609
timestamp 1649977179
transform 1 0 57132 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_615
timestamp 1649977179
transform 1 0 57684 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_617
timestamp 1649977179
transform 1 0 57868 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_629
timestamp 1649977179
transform 1 0 58972 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_641
timestamp 1649977179
transform 1 0 60076 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_653
timestamp 1649977179
transform 1 0 61180 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_665
timestamp 1649977179
transform 1 0 62284 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_671
timestamp 1649977179
transform 1 0 62836 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_673
timestamp 1649977179
transform 1 0 63020 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_685
timestamp 1649977179
transform 1 0 64124 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_697
timestamp 1649977179
transform 1 0 65228 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_709
timestamp 1649977179
transform 1 0 66332 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_721
timestamp 1649977179
transform 1 0 67436 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_727
timestamp 1649977179
transform 1 0 67988 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_729
timestamp 1649977179
transform 1 0 68172 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_741
timestamp 1649977179
transform 1 0 69276 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_753
timestamp 1649977179
transform 1 0 70380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_765
timestamp 1649977179
transform 1 0 71484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_777
timestamp 1649977179
transform 1 0 72588 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_783
timestamp 1649977179
transform 1 0 73140 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_785
timestamp 1649977179
transform 1 0 73324 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_797
timestamp 1649977179
transform 1 0 74428 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_809
timestamp 1649977179
transform 1 0 75532 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_821
timestamp 1649977179
transform 1 0 76636 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_123_829
timestamp 1649977179
transform 1 0 77372 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_123_836
timestamp 1649977179
transform 1 0 78016 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_841
timestamp 1649977179
transform 1 0 78476 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_124_7
timestamp 1649977179
transform 1 0 1748 0 1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_124_13
timestamp 1649977179
transform 1 0 2300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_124_25
timestamp 1649977179
transform 1 0 3404 0 1 69632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_124_29
timestamp 1649977179
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_41
timestamp 1649977179
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_53
timestamp 1649977179
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_65
timestamp 1649977179
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1649977179
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1649977179
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_85
timestamp 1649977179
transform 1 0 8924 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_97
timestamp 1649977179
transform 1 0 10028 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_109
timestamp 1649977179
transform 1 0 11132 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_121
timestamp 1649977179
transform 1 0 12236 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_133
timestamp 1649977179
transform 1 0 13340 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_139
timestamp 1649977179
transform 1 0 13892 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_141
timestamp 1649977179
transform 1 0 14076 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_153
timestamp 1649977179
transform 1 0 15180 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_165
timestamp 1649977179
transform 1 0 16284 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_177
timestamp 1649977179
transform 1 0 17388 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_189
timestamp 1649977179
transform 1 0 18492 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_195
timestamp 1649977179
transform 1 0 19044 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_197
timestamp 1649977179
transform 1 0 19228 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_209
timestamp 1649977179
transform 1 0 20332 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_221
timestamp 1649977179
transform 1 0 21436 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_233
timestamp 1649977179
transform 1 0 22540 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_245
timestamp 1649977179
transform 1 0 23644 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_251
timestamp 1649977179
transform 1 0 24196 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_253
timestamp 1649977179
transform 1 0 24380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_265
timestamp 1649977179
transform 1 0 25484 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_277
timestamp 1649977179
transform 1 0 26588 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_289
timestamp 1649977179
transform 1 0 27692 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_301
timestamp 1649977179
transform 1 0 28796 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_307
timestamp 1649977179
transform 1 0 29348 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_309
timestamp 1649977179
transform 1 0 29532 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_321
timestamp 1649977179
transform 1 0 30636 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_333
timestamp 1649977179
transform 1 0 31740 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_345
timestamp 1649977179
transform 1 0 32844 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_357
timestamp 1649977179
transform 1 0 33948 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_363
timestamp 1649977179
transform 1 0 34500 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_365
timestamp 1649977179
transform 1 0 34684 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_377
timestamp 1649977179
transform 1 0 35788 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_389
timestamp 1649977179
transform 1 0 36892 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_401
timestamp 1649977179
transform 1 0 37996 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_413
timestamp 1649977179
transform 1 0 39100 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_419
timestamp 1649977179
transform 1 0 39652 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_421
timestamp 1649977179
transform 1 0 39836 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_433
timestamp 1649977179
transform 1 0 40940 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_445
timestamp 1649977179
transform 1 0 42044 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_457
timestamp 1649977179
transform 1 0 43148 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_469
timestamp 1649977179
transform 1 0 44252 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_475
timestamp 1649977179
transform 1 0 44804 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_477
timestamp 1649977179
transform 1 0 44988 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_489
timestamp 1649977179
transform 1 0 46092 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_501
timestamp 1649977179
transform 1 0 47196 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_513
timestamp 1649977179
transform 1 0 48300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_525
timestamp 1649977179
transform 1 0 49404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_531
timestamp 1649977179
transform 1 0 49956 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_533
timestamp 1649977179
transform 1 0 50140 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_545
timestamp 1649977179
transform 1 0 51244 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_557
timestamp 1649977179
transform 1 0 52348 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_569
timestamp 1649977179
transform 1 0 53452 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_581
timestamp 1649977179
transform 1 0 54556 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_587
timestamp 1649977179
transform 1 0 55108 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_589
timestamp 1649977179
transform 1 0 55292 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_601
timestamp 1649977179
transform 1 0 56396 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_613
timestamp 1649977179
transform 1 0 57500 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_625
timestamp 1649977179
transform 1 0 58604 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_637
timestamp 1649977179
transform 1 0 59708 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_643
timestamp 1649977179
transform 1 0 60260 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_645
timestamp 1649977179
transform 1 0 60444 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_657
timestamp 1649977179
transform 1 0 61548 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_669
timestamp 1649977179
transform 1 0 62652 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_681
timestamp 1649977179
transform 1 0 63756 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_693
timestamp 1649977179
transform 1 0 64860 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_699
timestamp 1649977179
transform 1 0 65412 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_701
timestamp 1649977179
transform 1 0 65596 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_713
timestamp 1649977179
transform 1 0 66700 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_725
timestamp 1649977179
transform 1 0 67804 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_737
timestamp 1649977179
transform 1 0 68908 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_749
timestamp 1649977179
transform 1 0 70012 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_755
timestamp 1649977179
transform 1 0 70564 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_124_761
timestamp 1649977179
transform 1 0 71116 0 1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_124_767
timestamp 1649977179
transform 1 0 71668 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_779
timestamp 1649977179
transform 1 0 72772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_794
timestamp 1649977179
transform 1 0 74152 0 1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_124_800
timestamp 1649977179
transform 1 0 74704 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_813
timestamp 1649977179
transform 1 0 75900 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_825
timestamp 1649977179
transform 1 0 77004 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_124_831
timestamp 1649977179
transform 1 0 77556 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_124_838
timestamp 1649977179
transform 1 0 78200 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_125_7
timestamp 1649977179
transform 1 0 1748 0 -1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_125_13
timestamp 1649977179
transform 1 0 2300 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_25
timestamp 1649977179
transform 1 0 3404 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_37
timestamp 1649977179
transform 1 0 4508 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_49
timestamp 1649977179
transform 1 0 5612 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1649977179
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_57
timestamp 1649977179
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_69
timestamp 1649977179
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_81
timestamp 1649977179
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_93
timestamp 1649977179
transform 1 0 9660 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_105
timestamp 1649977179
transform 1 0 10764 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_111
timestamp 1649977179
transform 1 0 11316 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_113
timestamp 1649977179
transform 1 0 11500 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_125
timestamp 1649977179
transform 1 0 12604 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_137
timestamp 1649977179
transform 1 0 13708 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_149
timestamp 1649977179
transform 1 0 14812 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_161
timestamp 1649977179
transform 1 0 15916 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_167
timestamp 1649977179
transform 1 0 16468 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_169
timestamp 1649977179
transform 1 0 16652 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_181
timestamp 1649977179
transform 1 0 17756 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_193
timestamp 1649977179
transform 1 0 18860 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_205
timestamp 1649977179
transform 1 0 19964 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_217
timestamp 1649977179
transform 1 0 21068 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_223
timestamp 1649977179
transform 1 0 21620 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_225
timestamp 1649977179
transform 1 0 21804 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_237
timestamp 1649977179
transform 1 0 22908 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_249
timestamp 1649977179
transform 1 0 24012 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_261
timestamp 1649977179
transform 1 0 25116 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_273
timestamp 1649977179
transform 1 0 26220 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_279
timestamp 1649977179
transform 1 0 26772 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_281
timestamp 1649977179
transform 1 0 26956 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_293
timestamp 1649977179
transform 1 0 28060 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_305
timestamp 1649977179
transform 1 0 29164 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_317
timestamp 1649977179
transform 1 0 30268 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_329
timestamp 1649977179
transform 1 0 31372 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_335
timestamp 1649977179
transform 1 0 31924 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_337
timestamp 1649977179
transform 1 0 32108 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_349
timestamp 1649977179
transform 1 0 33212 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_361
timestamp 1649977179
transform 1 0 34316 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_373
timestamp 1649977179
transform 1 0 35420 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_385
timestamp 1649977179
transform 1 0 36524 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_391
timestamp 1649977179
transform 1 0 37076 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_393
timestamp 1649977179
transform 1 0 37260 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_405
timestamp 1649977179
transform 1 0 38364 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_417
timestamp 1649977179
transform 1 0 39468 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_429
timestamp 1649977179
transform 1 0 40572 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_441
timestamp 1649977179
transform 1 0 41676 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_447
timestamp 1649977179
transform 1 0 42228 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_449
timestamp 1649977179
transform 1 0 42412 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_461
timestamp 1649977179
transform 1 0 43516 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_473
timestamp 1649977179
transform 1 0 44620 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_485
timestamp 1649977179
transform 1 0 45724 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_497
timestamp 1649977179
transform 1 0 46828 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_503
timestamp 1649977179
transform 1 0 47380 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_505
timestamp 1649977179
transform 1 0 47564 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_517
timestamp 1649977179
transform 1 0 48668 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_529
timestamp 1649977179
transform 1 0 49772 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_541
timestamp 1649977179
transform 1 0 50876 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_553
timestamp 1649977179
transform 1 0 51980 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_559
timestamp 1649977179
transform 1 0 52532 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_561
timestamp 1649977179
transform 1 0 52716 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_573
timestamp 1649977179
transform 1 0 53820 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_585
timestamp 1649977179
transform 1 0 54924 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_597
timestamp 1649977179
transform 1 0 56028 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_609
timestamp 1649977179
transform 1 0 57132 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_615
timestamp 1649977179
transform 1 0 57684 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_617
timestamp 1649977179
transform 1 0 57868 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_629
timestamp 1649977179
transform 1 0 58972 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_641
timestamp 1649977179
transform 1 0 60076 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_653
timestamp 1649977179
transform 1 0 61180 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_665
timestamp 1649977179
transform 1 0 62284 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_671
timestamp 1649977179
transform 1 0 62836 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_673
timestamp 1649977179
transform 1 0 63020 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_685
timestamp 1649977179
transform 1 0 64124 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_697
timestamp 1649977179
transform 1 0 65228 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_709
timestamp 1649977179
transform 1 0 66332 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_721
timestamp 1649977179
transform 1 0 67436 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_727
timestamp 1649977179
transform 1 0 67988 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_729
timestamp 1649977179
transform 1 0 68172 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_741
timestamp 1649977179
transform 1 0 69276 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_753
timestamp 1649977179
transform 1 0 70380 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_125_765
timestamp 1649977179
transform 1 0 71484 0 -1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_125_771
timestamp 1649977179
transform 1 0 72036 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_783
timestamp 1649977179
transform 1 0 73140 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_785
timestamp 1649977179
transform 1 0 73324 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_125_797
timestamp 1649977179
transform 1 0 74428 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_125_802
timestamp 1649977179
transform 1 0 74888 0 -1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_125_808
timestamp 1649977179
transform 1 0 75440 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_820
timestamp 1649977179
transform 1 0 76544 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_836
timestamp 1649977179
transform 1 0 78016 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_841
timestamp 1649977179
transform 1 0 78476 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_126_7
timestamp 1649977179
transform 1 0 1748 0 1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_126_13
timestamp 1649977179
transform 1 0 2300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_126_25
timestamp 1649977179
transform 1 0 3404 0 1 70720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1649977179
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_41
timestamp 1649977179
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_53
timestamp 1649977179
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_65
timestamp 1649977179
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1649977179
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1649977179
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_85
timestamp 1649977179
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_97
timestamp 1649977179
transform 1 0 10028 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_109
timestamp 1649977179
transform 1 0 11132 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_121
timestamp 1649977179
transform 1 0 12236 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_133
timestamp 1649977179
transform 1 0 13340 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_139
timestamp 1649977179
transform 1 0 13892 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_141
timestamp 1649977179
transform 1 0 14076 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_153
timestamp 1649977179
transform 1 0 15180 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_165
timestamp 1649977179
transform 1 0 16284 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_177
timestamp 1649977179
transform 1 0 17388 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_189
timestamp 1649977179
transform 1 0 18492 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_195
timestamp 1649977179
transform 1 0 19044 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_197
timestamp 1649977179
transform 1 0 19228 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_209
timestamp 1649977179
transform 1 0 20332 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_221
timestamp 1649977179
transform 1 0 21436 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_233
timestamp 1649977179
transform 1 0 22540 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_245
timestamp 1649977179
transform 1 0 23644 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_251
timestamp 1649977179
transform 1 0 24196 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_253
timestamp 1649977179
transform 1 0 24380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_265
timestamp 1649977179
transform 1 0 25484 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_277
timestamp 1649977179
transform 1 0 26588 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_289
timestamp 1649977179
transform 1 0 27692 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_301
timestamp 1649977179
transform 1 0 28796 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_307
timestamp 1649977179
transform 1 0 29348 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_309
timestamp 1649977179
transform 1 0 29532 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_321
timestamp 1649977179
transform 1 0 30636 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_333
timestamp 1649977179
transform 1 0 31740 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_345
timestamp 1649977179
transform 1 0 32844 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_357
timestamp 1649977179
transform 1 0 33948 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_363
timestamp 1649977179
transform 1 0 34500 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_365
timestamp 1649977179
transform 1 0 34684 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_377
timestamp 1649977179
transform 1 0 35788 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_389
timestamp 1649977179
transform 1 0 36892 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_401
timestamp 1649977179
transform 1 0 37996 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_413
timestamp 1649977179
transform 1 0 39100 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_419
timestamp 1649977179
transform 1 0 39652 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_421
timestamp 1649977179
transform 1 0 39836 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_433
timestamp 1649977179
transform 1 0 40940 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_445
timestamp 1649977179
transform 1 0 42044 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_457
timestamp 1649977179
transform 1 0 43148 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_469
timestamp 1649977179
transform 1 0 44252 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_475
timestamp 1649977179
transform 1 0 44804 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_477
timestamp 1649977179
transform 1 0 44988 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_489
timestamp 1649977179
transform 1 0 46092 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_501
timestamp 1649977179
transform 1 0 47196 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_513
timestamp 1649977179
transform 1 0 48300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_525
timestamp 1649977179
transform 1 0 49404 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_531
timestamp 1649977179
transform 1 0 49956 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_533
timestamp 1649977179
transform 1 0 50140 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_545
timestamp 1649977179
transform 1 0 51244 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_557
timestamp 1649977179
transform 1 0 52348 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_569
timestamp 1649977179
transform 1 0 53452 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_581
timestamp 1649977179
transform 1 0 54556 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_587
timestamp 1649977179
transform 1 0 55108 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_589
timestamp 1649977179
transform 1 0 55292 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_601
timestamp 1649977179
transform 1 0 56396 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_613
timestamp 1649977179
transform 1 0 57500 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_625
timestamp 1649977179
transform 1 0 58604 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_637
timestamp 1649977179
transform 1 0 59708 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_643
timestamp 1649977179
transform 1 0 60260 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_645
timestamp 1649977179
transform 1 0 60444 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_657
timestamp 1649977179
transform 1 0 61548 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_669
timestamp 1649977179
transform 1 0 62652 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_681
timestamp 1649977179
transform 1 0 63756 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_693
timestamp 1649977179
transform 1 0 64860 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_699
timestamp 1649977179
transform 1 0 65412 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_701
timestamp 1649977179
transform 1 0 65596 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_713
timestamp 1649977179
transform 1 0 66700 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_725
timestamp 1649977179
transform 1 0 67804 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_737
timestamp 1649977179
transform 1 0 68908 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_749
timestamp 1649977179
transform 1 0 70012 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_755
timestamp 1649977179
transform 1 0 70564 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_126_757
timestamp 1649977179
transform 1 0 70748 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_126_765
timestamp 1649977179
transform 1 0 71484 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_126_772
timestamp 1649977179
transform 1 0 72128 0 1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_126_778
timestamp 1649977179
transform 1 0 72680 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_790
timestamp 1649977179
transform 1 0 73784 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_802
timestamp 1649977179
transform 1 0 74888 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_126_810
timestamp 1649977179
transform 1 0 75624 0 1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_126_816
timestamp 1649977179
transform 1 0 76176 0 1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_126_822
timestamp 1649977179
transform 1 0 76728 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_838
timestamp 1649977179
transform 1 0 78200 0 1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1649977179
transform 1 0 1380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_15
timestamp 1649977179
transform 1 0 2484 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_27
timestamp 1649977179
transform 1 0 3588 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_39
timestamp 1649977179
transform 1 0 4692 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_51
timestamp 1649977179
transform 1 0 5796 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1649977179
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_57
timestamp 1649977179
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_69
timestamp 1649977179
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_81
timestamp 1649977179
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_93
timestamp 1649977179
transform 1 0 9660 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_105
timestamp 1649977179
transform 1 0 10764 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_111
timestamp 1649977179
transform 1 0 11316 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_113
timestamp 1649977179
transform 1 0 11500 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_125
timestamp 1649977179
transform 1 0 12604 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_137
timestamp 1649977179
transform 1 0 13708 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_149
timestamp 1649977179
transform 1 0 14812 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_161
timestamp 1649977179
transform 1 0 15916 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_167
timestamp 1649977179
transform 1 0 16468 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_169
timestamp 1649977179
transform 1 0 16652 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_181
timestamp 1649977179
transform 1 0 17756 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_193
timestamp 1649977179
transform 1 0 18860 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_205
timestamp 1649977179
transform 1 0 19964 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_217
timestamp 1649977179
transform 1 0 21068 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_223
timestamp 1649977179
transform 1 0 21620 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_225
timestamp 1649977179
transform 1 0 21804 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_237
timestamp 1649977179
transform 1 0 22908 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_249
timestamp 1649977179
transform 1 0 24012 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_261
timestamp 1649977179
transform 1 0 25116 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_273
timestamp 1649977179
transform 1 0 26220 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_279
timestamp 1649977179
transform 1 0 26772 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_281
timestamp 1649977179
transform 1 0 26956 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_293
timestamp 1649977179
transform 1 0 28060 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_305
timestamp 1649977179
transform 1 0 29164 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_317
timestamp 1649977179
transform 1 0 30268 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_329
timestamp 1649977179
transform 1 0 31372 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_335
timestamp 1649977179
transform 1 0 31924 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_337
timestamp 1649977179
transform 1 0 32108 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_349
timestamp 1649977179
transform 1 0 33212 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_361
timestamp 1649977179
transform 1 0 34316 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_373
timestamp 1649977179
transform 1 0 35420 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_385
timestamp 1649977179
transform 1 0 36524 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_391
timestamp 1649977179
transform 1 0 37076 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_393
timestamp 1649977179
transform 1 0 37260 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_405
timestamp 1649977179
transform 1 0 38364 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_417
timestamp 1649977179
transform 1 0 39468 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_429
timestamp 1649977179
transform 1 0 40572 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_441
timestamp 1649977179
transform 1 0 41676 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_447
timestamp 1649977179
transform 1 0 42228 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_449
timestamp 1649977179
transform 1 0 42412 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_461
timestamp 1649977179
transform 1 0 43516 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_473
timestamp 1649977179
transform 1 0 44620 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_485
timestamp 1649977179
transform 1 0 45724 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_497
timestamp 1649977179
transform 1 0 46828 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_503
timestamp 1649977179
transform 1 0 47380 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_505
timestamp 1649977179
transform 1 0 47564 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_517
timestamp 1649977179
transform 1 0 48668 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_529
timestamp 1649977179
transform 1 0 49772 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_541
timestamp 1649977179
transform 1 0 50876 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_553
timestamp 1649977179
transform 1 0 51980 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_559
timestamp 1649977179
transform 1 0 52532 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_561
timestamp 1649977179
transform 1 0 52716 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_573
timestamp 1649977179
transform 1 0 53820 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_585
timestamp 1649977179
transform 1 0 54924 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_597
timestamp 1649977179
transform 1 0 56028 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_609
timestamp 1649977179
transform 1 0 57132 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_615
timestamp 1649977179
transform 1 0 57684 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_617
timestamp 1649977179
transform 1 0 57868 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_629
timestamp 1649977179
transform 1 0 58972 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_641
timestamp 1649977179
transform 1 0 60076 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_653
timestamp 1649977179
transform 1 0 61180 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_665
timestamp 1649977179
transform 1 0 62284 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_671
timestamp 1649977179
transform 1 0 62836 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_673
timestamp 1649977179
transform 1 0 63020 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_685
timestamp 1649977179
transform 1 0 64124 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_697
timestamp 1649977179
transform 1 0 65228 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_709
timestamp 1649977179
transform 1 0 66332 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_721
timestamp 1649977179
transform 1 0 67436 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_727
timestamp 1649977179
transform 1 0 67988 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_729
timestamp 1649977179
transform 1 0 68172 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_741
timestamp 1649977179
transform 1 0 69276 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_753
timestamp 1649977179
transform 1 0 70380 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_765
timestamp 1649977179
transform 1 0 71484 0 -1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_127_773
timestamp 1649977179
transform 1 0 72220 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_127_778
timestamp 1649977179
transform 1 0 72680 0 -1 71808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_127_787
timestamp 1649977179
transform 1 0 73508 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_799
timestamp 1649977179
transform 1 0 74612 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_811
timestamp 1649977179
transform 1 0 75716 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_817
timestamp 1649977179
transform 1 0 76268 0 -1 71808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_127_823
timestamp 1649977179
transform 1 0 76820 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_835
timestamp 1649977179
transform 1 0 77924 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_839
timestamp 1649977179
transform 1 0 78292 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_127_841
timestamp 1649977179
transform 1 0 78476 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_128_7
timestamp 1649977179
transform 1 0 1748 0 1 71808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_128_13
timestamp 1649977179
transform 1 0 2300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_128_25
timestamp 1649977179
transform 1 0 3404 0 1 71808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1649977179
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_41
timestamp 1649977179
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_53
timestamp 1649977179
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_65
timestamp 1649977179
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1649977179
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1649977179
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_85
timestamp 1649977179
transform 1 0 8924 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_97
timestamp 1649977179
transform 1 0 10028 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_109
timestamp 1649977179
transform 1 0 11132 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_121
timestamp 1649977179
transform 1 0 12236 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_133
timestamp 1649977179
transform 1 0 13340 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_139
timestamp 1649977179
transform 1 0 13892 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_141
timestamp 1649977179
transform 1 0 14076 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_153
timestamp 1649977179
transform 1 0 15180 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_165
timestamp 1649977179
transform 1 0 16284 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_177
timestamp 1649977179
transform 1 0 17388 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_189
timestamp 1649977179
transform 1 0 18492 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_195
timestamp 1649977179
transform 1 0 19044 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_197
timestamp 1649977179
transform 1 0 19228 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_209
timestamp 1649977179
transform 1 0 20332 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_221
timestamp 1649977179
transform 1 0 21436 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_233
timestamp 1649977179
transform 1 0 22540 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_245
timestamp 1649977179
transform 1 0 23644 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_251
timestamp 1649977179
transform 1 0 24196 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_253
timestamp 1649977179
transform 1 0 24380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_265
timestamp 1649977179
transform 1 0 25484 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_277
timestamp 1649977179
transform 1 0 26588 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_289
timestamp 1649977179
transform 1 0 27692 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_301
timestamp 1649977179
transform 1 0 28796 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_307
timestamp 1649977179
transform 1 0 29348 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_309
timestamp 1649977179
transform 1 0 29532 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_321
timestamp 1649977179
transform 1 0 30636 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_333
timestamp 1649977179
transform 1 0 31740 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_345
timestamp 1649977179
transform 1 0 32844 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_357
timestamp 1649977179
transform 1 0 33948 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_363
timestamp 1649977179
transform 1 0 34500 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_365
timestamp 1649977179
transform 1 0 34684 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_377
timestamp 1649977179
transform 1 0 35788 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_389
timestamp 1649977179
transform 1 0 36892 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_401
timestamp 1649977179
transform 1 0 37996 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_413
timestamp 1649977179
transform 1 0 39100 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_419
timestamp 1649977179
transform 1 0 39652 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_421
timestamp 1649977179
transform 1 0 39836 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_433
timestamp 1649977179
transform 1 0 40940 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_445
timestamp 1649977179
transform 1 0 42044 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_457
timestamp 1649977179
transform 1 0 43148 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_469
timestamp 1649977179
transform 1 0 44252 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_475
timestamp 1649977179
transform 1 0 44804 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_477
timestamp 1649977179
transform 1 0 44988 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_489
timestamp 1649977179
transform 1 0 46092 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_501
timestamp 1649977179
transform 1 0 47196 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_513
timestamp 1649977179
transform 1 0 48300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_525
timestamp 1649977179
transform 1 0 49404 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_531
timestamp 1649977179
transform 1 0 49956 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_533
timestamp 1649977179
transform 1 0 50140 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_545
timestamp 1649977179
transform 1 0 51244 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_557
timestamp 1649977179
transform 1 0 52348 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_569
timestamp 1649977179
transform 1 0 53452 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_581
timestamp 1649977179
transform 1 0 54556 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_587
timestamp 1649977179
transform 1 0 55108 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_589
timestamp 1649977179
transform 1 0 55292 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_601
timestamp 1649977179
transform 1 0 56396 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_613
timestamp 1649977179
transform 1 0 57500 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_625
timestamp 1649977179
transform 1 0 58604 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_637
timestamp 1649977179
transform 1 0 59708 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_643
timestamp 1649977179
transform 1 0 60260 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_645
timestamp 1649977179
transform 1 0 60444 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_657
timestamp 1649977179
transform 1 0 61548 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_669
timestamp 1649977179
transform 1 0 62652 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_681
timestamp 1649977179
transform 1 0 63756 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_693
timestamp 1649977179
transform 1 0 64860 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_699
timestamp 1649977179
transform 1 0 65412 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_701
timestamp 1649977179
transform 1 0 65596 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_713
timestamp 1649977179
transform 1 0 66700 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_725
timestamp 1649977179
transform 1 0 67804 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_737
timestamp 1649977179
transform 1 0 68908 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_749
timestamp 1649977179
transform 1 0 70012 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_755
timestamp 1649977179
transform 1 0 70564 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_757
timestamp 1649977179
transform 1 0 70748 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_769
timestamp 1649977179
transform 1 0 71852 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_781
timestamp 1649977179
transform 1 0 72956 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_793
timestamp 1649977179
transform 1 0 74060 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_805
timestamp 1649977179
transform 1 0 75164 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_811
timestamp 1649977179
transform 1 0 75716 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_813
timestamp 1649977179
transform 1 0 75900 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_825
timestamp 1649977179
transform 1 0 77004 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_833
timestamp 1649977179
transform 1 0 77740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_128_838
timestamp 1649977179
transform 1 0 78200 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_129_7
timestamp 1649977179
transform 1 0 1748 0 -1 72896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_129_13
timestamp 1649977179
transform 1 0 2300 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_25
timestamp 1649977179
transform 1 0 3404 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_37
timestamp 1649977179
transform 1 0 4508 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_49
timestamp 1649977179
transform 1 0 5612 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1649977179
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_57
timestamp 1649977179
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_69
timestamp 1649977179
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_81
timestamp 1649977179
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_93
timestamp 1649977179
transform 1 0 9660 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_105
timestamp 1649977179
transform 1 0 10764 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_111
timestamp 1649977179
transform 1 0 11316 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_113
timestamp 1649977179
transform 1 0 11500 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_125
timestamp 1649977179
transform 1 0 12604 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_137
timestamp 1649977179
transform 1 0 13708 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_149
timestamp 1649977179
transform 1 0 14812 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_161
timestamp 1649977179
transform 1 0 15916 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_167
timestamp 1649977179
transform 1 0 16468 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_169
timestamp 1649977179
transform 1 0 16652 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_181
timestamp 1649977179
transform 1 0 17756 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_193
timestamp 1649977179
transform 1 0 18860 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_205
timestamp 1649977179
transform 1 0 19964 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_217
timestamp 1649977179
transform 1 0 21068 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_223
timestamp 1649977179
transform 1 0 21620 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_225
timestamp 1649977179
transform 1 0 21804 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_237
timestamp 1649977179
transform 1 0 22908 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_249
timestamp 1649977179
transform 1 0 24012 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_261
timestamp 1649977179
transform 1 0 25116 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_273
timestamp 1649977179
transform 1 0 26220 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_279
timestamp 1649977179
transform 1 0 26772 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_281
timestamp 1649977179
transform 1 0 26956 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_293
timestamp 1649977179
transform 1 0 28060 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_305
timestamp 1649977179
transform 1 0 29164 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_317
timestamp 1649977179
transform 1 0 30268 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_329
timestamp 1649977179
transform 1 0 31372 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_335
timestamp 1649977179
transform 1 0 31924 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_337
timestamp 1649977179
transform 1 0 32108 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_349
timestamp 1649977179
transform 1 0 33212 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_361
timestamp 1649977179
transform 1 0 34316 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_373
timestamp 1649977179
transform 1 0 35420 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_385
timestamp 1649977179
transform 1 0 36524 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_391
timestamp 1649977179
transform 1 0 37076 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_393
timestamp 1649977179
transform 1 0 37260 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_405
timestamp 1649977179
transform 1 0 38364 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_417
timestamp 1649977179
transform 1 0 39468 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_429
timestamp 1649977179
transform 1 0 40572 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_441
timestamp 1649977179
transform 1 0 41676 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_447
timestamp 1649977179
transform 1 0 42228 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_449
timestamp 1649977179
transform 1 0 42412 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_461
timestamp 1649977179
transform 1 0 43516 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_473
timestamp 1649977179
transform 1 0 44620 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_485
timestamp 1649977179
transform 1 0 45724 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_497
timestamp 1649977179
transform 1 0 46828 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_503
timestamp 1649977179
transform 1 0 47380 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_505
timestamp 1649977179
transform 1 0 47564 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_517
timestamp 1649977179
transform 1 0 48668 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_529
timestamp 1649977179
transform 1 0 49772 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_541
timestamp 1649977179
transform 1 0 50876 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_553
timestamp 1649977179
transform 1 0 51980 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_559
timestamp 1649977179
transform 1 0 52532 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_561
timestamp 1649977179
transform 1 0 52716 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_573
timestamp 1649977179
transform 1 0 53820 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_585
timestamp 1649977179
transform 1 0 54924 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_597
timestamp 1649977179
transform 1 0 56028 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_609
timestamp 1649977179
transform 1 0 57132 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_615
timestamp 1649977179
transform 1 0 57684 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_617
timestamp 1649977179
transform 1 0 57868 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_629
timestamp 1649977179
transform 1 0 58972 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_641
timestamp 1649977179
transform 1 0 60076 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_653
timestamp 1649977179
transform 1 0 61180 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_665
timestamp 1649977179
transform 1 0 62284 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_671
timestamp 1649977179
transform 1 0 62836 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_673
timestamp 1649977179
transform 1 0 63020 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_685
timestamp 1649977179
transform 1 0 64124 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_697
timestamp 1649977179
transform 1 0 65228 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_709
timestamp 1649977179
transform 1 0 66332 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_721
timestamp 1649977179
transform 1 0 67436 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_727
timestamp 1649977179
transform 1 0 67988 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_729
timestamp 1649977179
transform 1 0 68172 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_741
timestamp 1649977179
transform 1 0 69276 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_753
timestamp 1649977179
transform 1 0 70380 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_765
timestamp 1649977179
transform 1 0 71484 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_777
timestamp 1649977179
transform 1 0 72588 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_783
timestamp 1649977179
transform 1 0 73140 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_785
timestamp 1649977179
transform 1 0 73324 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_797
timestamp 1649977179
transform 1 0 74428 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_809
timestamp 1649977179
transform 1 0 75532 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_821
timestamp 1649977179
transform 1 0 76636 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_129_829
timestamp 1649977179
transform 1 0 77372 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_836
timestamp 1649977179
transform 1 0 78016 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_841
timestamp 1649977179
transform 1 0 78476 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_130_7
timestamp 1649977179
transform 1 0 1748 0 1 72896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_130_13
timestamp 1649977179
transform 1 0 2300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_130_25
timestamp 1649977179
transform 1 0 3404 0 1 72896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1649977179
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_41
timestamp 1649977179
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_53
timestamp 1649977179
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_65
timestamp 1649977179
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1649977179
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1649977179
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_85
timestamp 1649977179
transform 1 0 8924 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_97
timestamp 1649977179
transform 1 0 10028 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_109
timestamp 1649977179
transform 1 0 11132 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_121
timestamp 1649977179
transform 1 0 12236 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_133
timestamp 1649977179
transform 1 0 13340 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_139
timestamp 1649977179
transform 1 0 13892 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_141
timestamp 1649977179
transform 1 0 14076 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_153
timestamp 1649977179
transform 1 0 15180 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_165
timestamp 1649977179
transform 1 0 16284 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_177
timestamp 1649977179
transform 1 0 17388 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_189
timestamp 1649977179
transform 1 0 18492 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_195
timestamp 1649977179
transform 1 0 19044 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_197
timestamp 1649977179
transform 1 0 19228 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_209
timestamp 1649977179
transform 1 0 20332 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_221
timestamp 1649977179
transform 1 0 21436 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_233
timestamp 1649977179
transform 1 0 22540 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_245
timestamp 1649977179
transform 1 0 23644 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_251
timestamp 1649977179
transform 1 0 24196 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_253
timestamp 1649977179
transform 1 0 24380 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_265
timestamp 1649977179
transform 1 0 25484 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_277
timestamp 1649977179
transform 1 0 26588 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_289
timestamp 1649977179
transform 1 0 27692 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_301
timestamp 1649977179
transform 1 0 28796 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_307
timestamp 1649977179
transform 1 0 29348 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_309
timestamp 1649977179
transform 1 0 29532 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_321
timestamp 1649977179
transform 1 0 30636 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_333
timestamp 1649977179
transform 1 0 31740 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_345
timestamp 1649977179
transform 1 0 32844 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_357
timestamp 1649977179
transform 1 0 33948 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_363
timestamp 1649977179
transform 1 0 34500 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_365
timestamp 1649977179
transform 1 0 34684 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_377
timestamp 1649977179
transform 1 0 35788 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_389
timestamp 1649977179
transform 1 0 36892 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_401
timestamp 1649977179
transform 1 0 37996 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_413
timestamp 1649977179
transform 1 0 39100 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_419
timestamp 1649977179
transform 1 0 39652 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_421
timestamp 1649977179
transform 1 0 39836 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_433
timestamp 1649977179
transform 1 0 40940 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_445
timestamp 1649977179
transform 1 0 42044 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_457
timestamp 1649977179
transform 1 0 43148 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_469
timestamp 1649977179
transform 1 0 44252 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_475
timestamp 1649977179
transform 1 0 44804 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_477
timestamp 1649977179
transform 1 0 44988 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_489
timestamp 1649977179
transform 1 0 46092 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_501
timestamp 1649977179
transform 1 0 47196 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_513
timestamp 1649977179
transform 1 0 48300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_525
timestamp 1649977179
transform 1 0 49404 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_531
timestamp 1649977179
transform 1 0 49956 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_533
timestamp 1649977179
transform 1 0 50140 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_545
timestamp 1649977179
transform 1 0 51244 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_557
timestamp 1649977179
transform 1 0 52348 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_569
timestamp 1649977179
transform 1 0 53452 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_581
timestamp 1649977179
transform 1 0 54556 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_587
timestamp 1649977179
transform 1 0 55108 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_589
timestamp 1649977179
transform 1 0 55292 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_601
timestamp 1649977179
transform 1 0 56396 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_613
timestamp 1649977179
transform 1 0 57500 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_625
timestamp 1649977179
transform 1 0 58604 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_637
timestamp 1649977179
transform 1 0 59708 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_643
timestamp 1649977179
transform 1 0 60260 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_645
timestamp 1649977179
transform 1 0 60444 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_657
timestamp 1649977179
transform 1 0 61548 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_669
timestamp 1649977179
transform 1 0 62652 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_681
timestamp 1649977179
transform 1 0 63756 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_693
timestamp 1649977179
transform 1 0 64860 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_699
timestamp 1649977179
transform 1 0 65412 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_701
timestamp 1649977179
transform 1 0 65596 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_713
timestamp 1649977179
transform 1 0 66700 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_725
timestamp 1649977179
transform 1 0 67804 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_737
timestamp 1649977179
transform 1 0 68908 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_749
timestamp 1649977179
transform 1 0 70012 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_755
timestamp 1649977179
transform 1 0 70564 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_757
timestamp 1649977179
transform 1 0 70748 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_769
timestamp 1649977179
transform 1 0 71852 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_781
timestamp 1649977179
transform 1 0 72956 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_793
timestamp 1649977179
transform 1 0 74060 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_805
timestamp 1649977179
transform 1 0 75164 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_811
timestamp 1649977179
transform 1 0 75716 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_813
timestamp 1649977179
transform 1 0 75900 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_825
timestamp 1649977179
transform 1 0 77004 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_833
timestamp 1649977179
transform 1 0 77740 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_130_838
timestamp 1649977179
transform 1 0 78200 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_131_7
timestamp 1649977179
transform 1 0 1748 0 -1 73984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_131_13
timestamp 1649977179
transform 1 0 2300 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_25
timestamp 1649977179
transform 1 0 3404 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_37
timestamp 1649977179
transform 1 0 4508 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_49
timestamp 1649977179
transform 1 0 5612 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_55
timestamp 1649977179
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_57
timestamp 1649977179
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_69
timestamp 1649977179
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_81
timestamp 1649977179
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_93
timestamp 1649977179
transform 1 0 9660 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_105
timestamp 1649977179
transform 1 0 10764 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_111
timestamp 1649977179
transform 1 0 11316 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_113
timestamp 1649977179
transform 1 0 11500 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_125
timestamp 1649977179
transform 1 0 12604 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_137
timestamp 1649977179
transform 1 0 13708 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_149
timestamp 1649977179
transform 1 0 14812 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_161
timestamp 1649977179
transform 1 0 15916 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_167
timestamp 1649977179
transform 1 0 16468 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_169
timestamp 1649977179
transform 1 0 16652 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_181
timestamp 1649977179
transform 1 0 17756 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_193
timestamp 1649977179
transform 1 0 18860 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_205
timestamp 1649977179
transform 1 0 19964 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_217
timestamp 1649977179
transform 1 0 21068 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_223
timestamp 1649977179
transform 1 0 21620 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_225
timestamp 1649977179
transform 1 0 21804 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_237
timestamp 1649977179
transform 1 0 22908 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_249
timestamp 1649977179
transform 1 0 24012 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_261
timestamp 1649977179
transform 1 0 25116 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_273
timestamp 1649977179
transform 1 0 26220 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_279
timestamp 1649977179
transform 1 0 26772 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_281
timestamp 1649977179
transform 1 0 26956 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_293
timestamp 1649977179
transform 1 0 28060 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_305
timestamp 1649977179
transform 1 0 29164 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_317
timestamp 1649977179
transform 1 0 30268 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_329
timestamp 1649977179
transform 1 0 31372 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_335
timestamp 1649977179
transform 1 0 31924 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_337
timestamp 1649977179
transform 1 0 32108 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_349
timestamp 1649977179
transform 1 0 33212 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_361
timestamp 1649977179
transform 1 0 34316 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_373
timestamp 1649977179
transform 1 0 35420 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_385
timestamp 1649977179
transform 1 0 36524 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_391
timestamp 1649977179
transform 1 0 37076 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_393
timestamp 1649977179
transform 1 0 37260 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_405
timestamp 1649977179
transform 1 0 38364 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_417
timestamp 1649977179
transform 1 0 39468 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_429
timestamp 1649977179
transform 1 0 40572 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_441
timestamp 1649977179
transform 1 0 41676 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_447
timestamp 1649977179
transform 1 0 42228 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_449
timestamp 1649977179
transform 1 0 42412 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_461
timestamp 1649977179
transform 1 0 43516 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_473
timestamp 1649977179
transform 1 0 44620 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_485
timestamp 1649977179
transform 1 0 45724 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_497
timestamp 1649977179
transform 1 0 46828 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_503
timestamp 1649977179
transform 1 0 47380 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_505
timestamp 1649977179
transform 1 0 47564 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_517
timestamp 1649977179
transform 1 0 48668 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_529
timestamp 1649977179
transform 1 0 49772 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_541
timestamp 1649977179
transform 1 0 50876 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_553
timestamp 1649977179
transform 1 0 51980 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_559
timestamp 1649977179
transform 1 0 52532 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_561
timestamp 1649977179
transform 1 0 52716 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_573
timestamp 1649977179
transform 1 0 53820 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_585
timestamp 1649977179
transform 1 0 54924 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_597
timestamp 1649977179
transform 1 0 56028 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_609
timestamp 1649977179
transform 1 0 57132 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_615
timestamp 1649977179
transform 1 0 57684 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_617
timestamp 1649977179
transform 1 0 57868 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_629
timestamp 1649977179
transform 1 0 58972 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_641
timestamp 1649977179
transform 1 0 60076 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_653
timestamp 1649977179
transform 1 0 61180 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_665
timestamp 1649977179
transform 1 0 62284 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_671
timestamp 1649977179
transform 1 0 62836 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_673
timestamp 1649977179
transform 1 0 63020 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_685
timestamp 1649977179
transform 1 0 64124 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_697
timestamp 1649977179
transform 1 0 65228 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_709
timestamp 1649977179
transform 1 0 66332 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_721
timestamp 1649977179
transform 1 0 67436 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_727
timestamp 1649977179
transform 1 0 67988 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_729
timestamp 1649977179
transform 1 0 68172 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_741
timestamp 1649977179
transform 1 0 69276 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_753
timestamp 1649977179
transform 1 0 70380 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_765
timestamp 1649977179
transform 1 0 71484 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_777
timestamp 1649977179
transform 1 0 72588 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_783
timestamp 1649977179
transform 1 0 73140 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_785
timestamp 1649977179
transform 1 0 73324 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_797
timestamp 1649977179
transform 1 0 74428 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_809
timestamp 1649977179
transform 1 0 75532 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_821
timestamp 1649977179
transform 1 0 76636 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_825
timestamp 1649977179
transform 1 0 77004 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_131_828
timestamp 1649977179
transform 1 0 77280 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_131_836
timestamp 1649977179
transform 1 0 78016 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_841
timestamp 1649977179
transform 1 0 78476 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_5
timestamp 1649977179
transform 1 0 1564 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_17
timestamp 1649977179
transform 1 0 2668 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_132_25
timestamp 1649977179
transform 1 0 3404 0 1 73984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1649977179
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_41
timestamp 1649977179
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_53
timestamp 1649977179
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_65
timestamp 1649977179
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1649977179
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1649977179
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_85
timestamp 1649977179
transform 1 0 8924 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_97
timestamp 1649977179
transform 1 0 10028 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_109
timestamp 1649977179
transform 1 0 11132 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_121
timestamp 1649977179
transform 1 0 12236 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_133
timestamp 1649977179
transform 1 0 13340 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_139
timestamp 1649977179
transform 1 0 13892 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_141
timestamp 1649977179
transform 1 0 14076 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_153
timestamp 1649977179
transform 1 0 15180 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_165
timestamp 1649977179
transform 1 0 16284 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_177
timestamp 1649977179
transform 1 0 17388 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_189
timestamp 1649977179
transform 1 0 18492 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_195
timestamp 1649977179
transform 1 0 19044 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_197
timestamp 1649977179
transform 1 0 19228 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_209
timestamp 1649977179
transform 1 0 20332 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_221
timestamp 1649977179
transform 1 0 21436 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_233
timestamp 1649977179
transform 1 0 22540 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_245
timestamp 1649977179
transform 1 0 23644 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_251
timestamp 1649977179
transform 1 0 24196 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_253
timestamp 1649977179
transform 1 0 24380 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_265
timestamp 1649977179
transform 1 0 25484 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_277
timestamp 1649977179
transform 1 0 26588 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_289
timestamp 1649977179
transform 1 0 27692 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_301
timestamp 1649977179
transform 1 0 28796 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_307
timestamp 1649977179
transform 1 0 29348 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_309
timestamp 1649977179
transform 1 0 29532 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_321
timestamp 1649977179
transform 1 0 30636 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_333
timestamp 1649977179
transform 1 0 31740 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_345
timestamp 1649977179
transform 1 0 32844 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_357
timestamp 1649977179
transform 1 0 33948 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_363
timestamp 1649977179
transform 1 0 34500 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_365
timestamp 1649977179
transform 1 0 34684 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_377
timestamp 1649977179
transform 1 0 35788 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_389
timestamp 1649977179
transform 1 0 36892 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_401
timestamp 1649977179
transform 1 0 37996 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_413
timestamp 1649977179
transform 1 0 39100 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_419
timestamp 1649977179
transform 1 0 39652 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_421
timestamp 1649977179
transform 1 0 39836 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_433
timestamp 1649977179
transform 1 0 40940 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_445
timestamp 1649977179
transform 1 0 42044 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_457
timestamp 1649977179
transform 1 0 43148 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_469
timestamp 1649977179
transform 1 0 44252 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_475
timestamp 1649977179
transform 1 0 44804 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_477
timestamp 1649977179
transform 1 0 44988 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_489
timestamp 1649977179
transform 1 0 46092 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_501
timestamp 1649977179
transform 1 0 47196 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_513
timestamp 1649977179
transform 1 0 48300 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_525
timestamp 1649977179
transform 1 0 49404 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_531
timestamp 1649977179
transform 1 0 49956 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_533
timestamp 1649977179
transform 1 0 50140 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_545
timestamp 1649977179
transform 1 0 51244 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_557
timestamp 1649977179
transform 1 0 52348 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_569
timestamp 1649977179
transform 1 0 53452 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_581
timestamp 1649977179
transform 1 0 54556 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_587
timestamp 1649977179
transform 1 0 55108 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_589
timestamp 1649977179
transform 1 0 55292 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_601
timestamp 1649977179
transform 1 0 56396 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_613
timestamp 1649977179
transform 1 0 57500 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_625
timestamp 1649977179
transform 1 0 58604 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_637
timestamp 1649977179
transform 1 0 59708 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_643
timestamp 1649977179
transform 1 0 60260 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_645
timestamp 1649977179
transform 1 0 60444 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_657
timestamp 1649977179
transform 1 0 61548 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_669
timestamp 1649977179
transform 1 0 62652 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_681
timestamp 1649977179
transform 1 0 63756 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_693
timestamp 1649977179
transform 1 0 64860 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_699
timestamp 1649977179
transform 1 0 65412 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_701
timestamp 1649977179
transform 1 0 65596 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_713
timestamp 1649977179
transform 1 0 66700 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_725
timestamp 1649977179
transform 1 0 67804 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_737
timestamp 1649977179
transform 1 0 68908 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_749
timestamp 1649977179
transform 1 0 70012 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_755
timestamp 1649977179
transform 1 0 70564 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_757
timestamp 1649977179
transform 1 0 70748 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_769
timestamp 1649977179
transform 1 0 71852 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_781
timestamp 1649977179
transform 1 0 72956 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_793
timestamp 1649977179
transform 1 0 74060 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_805
timestamp 1649977179
transform 1 0 75164 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_811
timestamp 1649977179
transform 1 0 75716 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_813
timestamp 1649977179
transform 1 0 75900 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_825
timestamp 1649977179
transform 1 0 77004 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_132_833
timestamp 1649977179
transform 1 0 77740 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_838
timestamp 1649977179
transform 1 0 78200 0 1 73984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_133_7
timestamp 1649977179
transform 1 0 1748 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_19
timestamp 1649977179
transform 1 0 2852 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_31
timestamp 1649977179
transform 1 0 3956 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_43
timestamp 1649977179
transform 1 0 5060 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_133_55
timestamp 1649977179
transform 1 0 6164 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_57
timestamp 1649977179
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_69
timestamp 1649977179
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_81
timestamp 1649977179
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_93
timestamp 1649977179
transform 1 0 9660 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_105
timestamp 1649977179
transform 1 0 10764 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_111
timestamp 1649977179
transform 1 0 11316 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_113
timestamp 1649977179
transform 1 0 11500 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_125
timestamp 1649977179
transform 1 0 12604 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_137
timestamp 1649977179
transform 1 0 13708 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_149
timestamp 1649977179
transform 1 0 14812 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_161
timestamp 1649977179
transform 1 0 15916 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_167
timestamp 1649977179
transform 1 0 16468 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_169
timestamp 1649977179
transform 1 0 16652 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_181
timestamp 1649977179
transform 1 0 17756 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_193
timestamp 1649977179
transform 1 0 18860 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_205
timestamp 1649977179
transform 1 0 19964 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_217
timestamp 1649977179
transform 1 0 21068 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_223
timestamp 1649977179
transform 1 0 21620 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_225
timestamp 1649977179
transform 1 0 21804 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_237
timestamp 1649977179
transform 1 0 22908 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_249
timestamp 1649977179
transform 1 0 24012 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_261
timestamp 1649977179
transform 1 0 25116 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_273
timestamp 1649977179
transform 1 0 26220 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_279
timestamp 1649977179
transform 1 0 26772 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_281
timestamp 1649977179
transform 1 0 26956 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_293
timestamp 1649977179
transform 1 0 28060 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_305
timestamp 1649977179
transform 1 0 29164 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_317
timestamp 1649977179
transform 1 0 30268 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_329
timestamp 1649977179
transform 1 0 31372 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_335
timestamp 1649977179
transform 1 0 31924 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_337
timestamp 1649977179
transform 1 0 32108 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_349
timestamp 1649977179
transform 1 0 33212 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_361
timestamp 1649977179
transform 1 0 34316 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_373
timestamp 1649977179
transform 1 0 35420 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_385
timestamp 1649977179
transform 1 0 36524 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_391
timestamp 1649977179
transform 1 0 37076 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_393
timestamp 1649977179
transform 1 0 37260 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_405
timestamp 1649977179
transform 1 0 38364 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_417
timestamp 1649977179
transform 1 0 39468 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_429
timestamp 1649977179
transform 1 0 40572 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_441
timestamp 1649977179
transform 1 0 41676 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_447
timestamp 1649977179
transform 1 0 42228 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_449
timestamp 1649977179
transform 1 0 42412 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_461
timestamp 1649977179
transform 1 0 43516 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_473
timestamp 1649977179
transform 1 0 44620 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_485
timestamp 1649977179
transform 1 0 45724 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_497
timestamp 1649977179
transform 1 0 46828 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_503
timestamp 1649977179
transform 1 0 47380 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_505
timestamp 1649977179
transform 1 0 47564 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_517
timestamp 1649977179
transform 1 0 48668 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_529
timestamp 1649977179
transform 1 0 49772 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_541
timestamp 1649977179
transform 1 0 50876 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_553
timestamp 1649977179
transform 1 0 51980 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_559
timestamp 1649977179
transform 1 0 52532 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_561
timestamp 1649977179
transform 1 0 52716 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_573
timestamp 1649977179
transform 1 0 53820 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_585
timestamp 1649977179
transform 1 0 54924 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_597
timestamp 1649977179
transform 1 0 56028 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_609
timestamp 1649977179
transform 1 0 57132 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_615
timestamp 1649977179
transform 1 0 57684 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_617
timestamp 1649977179
transform 1 0 57868 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_629
timestamp 1649977179
transform 1 0 58972 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_641
timestamp 1649977179
transform 1 0 60076 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_653
timestamp 1649977179
transform 1 0 61180 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_665
timestamp 1649977179
transform 1 0 62284 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_671
timestamp 1649977179
transform 1 0 62836 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_673
timestamp 1649977179
transform 1 0 63020 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_685
timestamp 1649977179
transform 1 0 64124 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_697
timestamp 1649977179
transform 1 0 65228 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_709
timestamp 1649977179
transform 1 0 66332 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_721
timestamp 1649977179
transform 1 0 67436 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_727
timestamp 1649977179
transform 1 0 67988 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_729
timestamp 1649977179
transform 1 0 68172 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_741
timestamp 1649977179
transform 1 0 69276 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_753
timestamp 1649977179
transform 1 0 70380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_765
timestamp 1649977179
transform 1 0 71484 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_777
timestamp 1649977179
transform 1 0 72588 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_783
timestamp 1649977179
transform 1 0 73140 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_785
timestamp 1649977179
transform 1 0 73324 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_797
timestamp 1649977179
transform 1 0 74428 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_809
timestamp 1649977179
transform 1 0 75532 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_821
timestamp 1649977179
transform 1 0 76636 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_133_829
timestamp 1649977179
transform 1 0 77372 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_133_836
timestamp 1649977179
transform 1 0 78016 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_841
timestamp 1649977179
transform 1 0 78476 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_134_7
timestamp 1649977179
transform 1 0 1748 0 1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_134_13
timestamp 1649977179
transform 1 0 2300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_134_25
timestamp 1649977179
transform 1 0 3404 0 1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1649977179
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_41
timestamp 1649977179
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_53
timestamp 1649977179
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_65
timestamp 1649977179
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1649977179
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1649977179
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_85
timestamp 1649977179
transform 1 0 8924 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_97
timestamp 1649977179
transform 1 0 10028 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_109
timestamp 1649977179
transform 1 0 11132 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_121
timestamp 1649977179
transform 1 0 12236 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_133
timestamp 1649977179
transform 1 0 13340 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_139
timestamp 1649977179
transform 1 0 13892 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_141
timestamp 1649977179
transform 1 0 14076 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_153
timestamp 1649977179
transform 1 0 15180 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_165
timestamp 1649977179
transform 1 0 16284 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_177
timestamp 1649977179
transform 1 0 17388 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_189
timestamp 1649977179
transform 1 0 18492 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_195
timestamp 1649977179
transform 1 0 19044 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_197
timestamp 1649977179
transform 1 0 19228 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_209
timestamp 1649977179
transform 1 0 20332 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_221
timestamp 1649977179
transform 1 0 21436 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_233
timestamp 1649977179
transform 1 0 22540 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_245
timestamp 1649977179
transform 1 0 23644 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_251
timestamp 1649977179
transform 1 0 24196 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_253
timestamp 1649977179
transform 1 0 24380 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_265
timestamp 1649977179
transform 1 0 25484 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_277
timestamp 1649977179
transform 1 0 26588 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_289
timestamp 1649977179
transform 1 0 27692 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_301
timestamp 1649977179
transform 1 0 28796 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_307
timestamp 1649977179
transform 1 0 29348 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_309
timestamp 1649977179
transform 1 0 29532 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_321
timestamp 1649977179
transform 1 0 30636 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_333
timestamp 1649977179
transform 1 0 31740 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_345
timestamp 1649977179
transform 1 0 32844 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_357
timestamp 1649977179
transform 1 0 33948 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_363
timestamp 1649977179
transform 1 0 34500 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_365
timestamp 1649977179
transform 1 0 34684 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_377
timestamp 1649977179
transform 1 0 35788 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_389
timestamp 1649977179
transform 1 0 36892 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_401
timestamp 1649977179
transform 1 0 37996 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_413
timestamp 1649977179
transform 1 0 39100 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_419
timestamp 1649977179
transform 1 0 39652 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_421
timestamp 1649977179
transform 1 0 39836 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_433
timestamp 1649977179
transform 1 0 40940 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_445
timestamp 1649977179
transform 1 0 42044 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_457
timestamp 1649977179
transform 1 0 43148 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_469
timestamp 1649977179
transform 1 0 44252 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_475
timestamp 1649977179
transform 1 0 44804 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_477
timestamp 1649977179
transform 1 0 44988 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_489
timestamp 1649977179
transform 1 0 46092 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_501
timestamp 1649977179
transform 1 0 47196 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_513
timestamp 1649977179
transform 1 0 48300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_525
timestamp 1649977179
transform 1 0 49404 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_531
timestamp 1649977179
transform 1 0 49956 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_533
timestamp 1649977179
transform 1 0 50140 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_545
timestamp 1649977179
transform 1 0 51244 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_557
timestamp 1649977179
transform 1 0 52348 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_569
timestamp 1649977179
transform 1 0 53452 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_581
timestamp 1649977179
transform 1 0 54556 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_587
timestamp 1649977179
transform 1 0 55108 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_589
timestamp 1649977179
transform 1 0 55292 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_601
timestamp 1649977179
transform 1 0 56396 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_613
timestamp 1649977179
transform 1 0 57500 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_625
timestamp 1649977179
transform 1 0 58604 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_637
timestamp 1649977179
transform 1 0 59708 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_643
timestamp 1649977179
transform 1 0 60260 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_645
timestamp 1649977179
transform 1 0 60444 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_657
timestamp 1649977179
transform 1 0 61548 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_669
timestamp 1649977179
transform 1 0 62652 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_681
timestamp 1649977179
transform 1 0 63756 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_693
timestamp 1649977179
transform 1 0 64860 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_699
timestamp 1649977179
transform 1 0 65412 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_701
timestamp 1649977179
transform 1 0 65596 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_713
timestamp 1649977179
transform 1 0 66700 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_725
timestamp 1649977179
transform 1 0 67804 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_737
timestamp 1649977179
transform 1 0 68908 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_749
timestamp 1649977179
transform 1 0 70012 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_755
timestamp 1649977179
transform 1 0 70564 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_757
timestamp 1649977179
transform 1 0 70748 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_769
timestamp 1649977179
transform 1 0 71852 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_781
timestamp 1649977179
transform 1 0 72956 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_793
timestamp 1649977179
transform 1 0 74060 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_805
timestamp 1649977179
transform 1 0 75164 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_811
timestamp 1649977179
transform 1 0 75716 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_813
timestamp 1649977179
transform 1 0 75900 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_134_825
timestamp 1649977179
transform 1 0 77004 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_830
timestamp 1649977179
transform 1 0 77464 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_134_838
timestamp 1649977179
transform 1 0 78200 0 1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_135_3
timestamp 1649977179
transform 1 0 1380 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_15
timestamp 1649977179
transform 1 0 2484 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_27
timestamp 1649977179
transform 1 0 3588 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_39
timestamp 1649977179
transform 1 0 4692 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_51
timestamp 1649977179
transform 1 0 5796 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_55
timestamp 1649977179
transform 1 0 6164 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_57
timestamp 1649977179
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_69
timestamp 1649977179
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_81
timestamp 1649977179
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_93
timestamp 1649977179
transform 1 0 9660 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_105
timestamp 1649977179
transform 1 0 10764 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_111
timestamp 1649977179
transform 1 0 11316 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_113
timestamp 1649977179
transform 1 0 11500 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_125
timestamp 1649977179
transform 1 0 12604 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_137
timestamp 1649977179
transform 1 0 13708 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_149
timestamp 1649977179
transform 1 0 14812 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_161
timestamp 1649977179
transform 1 0 15916 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_167
timestamp 1649977179
transform 1 0 16468 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_169
timestamp 1649977179
transform 1 0 16652 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_181
timestamp 1649977179
transform 1 0 17756 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_193
timestamp 1649977179
transform 1 0 18860 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_205
timestamp 1649977179
transform 1 0 19964 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_217
timestamp 1649977179
transform 1 0 21068 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_223
timestamp 1649977179
transform 1 0 21620 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_225
timestamp 1649977179
transform 1 0 21804 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_237
timestamp 1649977179
transform 1 0 22908 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_249
timestamp 1649977179
transform 1 0 24012 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_261
timestamp 1649977179
transform 1 0 25116 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_273
timestamp 1649977179
transform 1 0 26220 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_279
timestamp 1649977179
transform 1 0 26772 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_281
timestamp 1649977179
transform 1 0 26956 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_293
timestamp 1649977179
transform 1 0 28060 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_305
timestamp 1649977179
transform 1 0 29164 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_317
timestamp 1649977179
transform 1 0 30268 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_329
timestamp 1649977179
transform 1 0 31372 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_335
timestamp 1649977179
transform 1 0 31924 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_337
timestamp 1649977179
transform 1 0 32108 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_349
timestamp 1649977179
transform 1 0 33212 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_361
timestamp 1649977179
transform 1 0 34316 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_373
timestamp 1649977179
transform 1 0 35420 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_385
timestamp 1649977179
transform 1 0 36524 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_391
timestamp 1649977179
transform 1 0 37076 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_393
timestamp 1649977179
transform 1 0 37260 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_405
timestamp 1649977179
transform 1 0 38364 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_417
timestamp 1649977179
transform 1 0 39468 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_429
timestamp 1649977179
transform 1 0 40572 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_441
timestamp 1649977179
transform 1 0 41676 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_447
timestamp 1649977179
transform 1 0 42228 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_449
timestamp 1649977179
transform 1 0 42412 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_461
timestamp 1649977179
transform 1 0 43516 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_473
timestamp 1649977179
transform 1 0 44620 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_485
timestamp 1649977179
transform 1 0 45724 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_497
timestamp 1649977179
transform 1 0 46828 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_503
timestamp 1649977179
transform 1 0 47380 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_505
timestamp 1649977179
transform 1 0 47564 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_517
timestamp 1649977179
transform 1 0 48668 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_529
timestamp 1649977179
transform 1 0 49772 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_541
timestamp 1649977179
transform 1 0 50876 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_553
timestamp 1649977179
transform 1 0 51980 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_559
timestamp 1649977179
transform 1 0 52532 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_561
timestamp 1649977179
transform 1 0 52716 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_573
timestamp 1649977179
transform 1 0 53820 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_585
timestamp 1649977179
transform 1 0 54924 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_597
timestamp 1649977179
transform 1 0 56028 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_609
timestamp 1649977179
transform 1 0 57132 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_615
timestamp 1649977179
transform 1 0 57684 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_617
timestamp 1649977179
transform 1 0 57868 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_629
timestamp 1649977179
transform 1 0 58972 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_641
timestamp 1649977179
transform 1 0 60076 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_653
timestamp 1649977179
transform 1 0 61180 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_665
timestamp 1649977179
transform 1 0 62284 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_671
timestamp 1649977179
transform 1 0 62836 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_673
timestamp 1649977179
transform 1 0 63020 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_685
timestamp 1649977179
transform 1 0 64124 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_697
timestamp 1649977179
transform 1 0 65228 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_709
timestamp 1649977179
transform 1 0 66332 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_721
timestamp 1649977179
transform 1 0 67436 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_727
timestamp 1649977179
transform 1 0 67988 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_729
timestamp 1649977179
transform 1 0 68172 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_741
timestamp 1649977179
transform 1 0 69276 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_753
timestamp 1649977179
transform 1 0 70380 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_765
timestamp 1649977179
transform 1 0 71484 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_777
timestamp 1649977179
transform 1 0 72588 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_783
timestamp 1649977179
transform 1 0 73140 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_785
timestamp 1649977179
transform 1 0 73324 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_797
timestamp 1649977179
transform 1 0 74428 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_809
timestamp 1649977179
transform 1 0 75532 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_821
timestamp 1649977179
transform 1 0 76636 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_833
timestamp 1649977179
transform 1 0 77740 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_839
timestamp 1649977179
transform 1 0 78292 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_135_841
timestamp 1649977179
transform 1 0 78476 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_3
timestamp 1649977179
transform 1 0 1380 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_15
timestamp 1649977179
transform 1 0 2484 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1649977179
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1649977179
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_41
timestamp 1649977179
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_53
timestamp 1649977179
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_65
timestamp 1649977179
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1649977179
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1649977179
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_85
timestamp 1649977179
transform 1 0 8924 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_97
timestamp 1649977179
transform 1 0 10028 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_109
timestamp 1649977179
transform 1 0 11132 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_121
timestamp 1649977179
transform 1 0 12236 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_133
timestamp 1649977179
transform 1 0 13340 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_139
timestamp 1649977179
transform 1 0 13892 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_141
timestamp 1649977179
transform 1 0 14076 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_153
timestamp 1649977179
transform 1 0 15180 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_165
timestamp 1649977179
transform 1 0 16284 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_177
timestamp 1649977179
transform 1 0 17388 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_189
timestamp 1649977179
transform 1 0 18492 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_195
timestamp 1649977179
transform 1 0 19044 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_197
timestamp 1649977179
transform 1 0 19228 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_209
timestamp 1649977179
transform 1 0 20332 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_221
timestamp 1649977179
transform 1 0 21436 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_233
timestamp 1649977179
transform 1 0 22540 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_245
timestamp 1649977179
transform 1 0 23644 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_251
timestamp 1649977179
transform 1 0 24196 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_253
timestamp 1649977179
transform 1 0 24380 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_265
timestamp 1649977179
transform 1 0 25484 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_277
timestamp 1649977179
transform 1 0 26588 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_289
timestamp 1649977179
transform 1 0 27692 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_301
timestamp 1649977179
transform 1 0 28796 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_307
timestamp 1649977179
transform 1 0 29348 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_309
timestamp 1649977179
transform 1 0 29532 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_321
timestamp 1649977179
transform 1 0 30636 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_333
timestamp 1649977179
transform 1 0 31740 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_345
timestamp 1649977179
transform 1 0 32844 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_357
timestamp 1649977179
transform 1 0 33948 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_363
timestamp 1649977179
transform 1 0 34500 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_365
timestamp 1649977179
transform 1 0 34684 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_377
timestamp 1649977179
transform 1 0 35788 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_389
timestamp 1649977179
transform 1 0 36892 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_401
timestamp 1649977179
transform 1 0 37996 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_413
timestamp 1649977179
transform 1 0 39100 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_419
timestamp 1649977179
transform 1 0 39652 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_421
timestamp 1649977179
transform 1 0 39836 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_433
timestamp 1649977179
transform 1 0 40940 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_445
timestamp 1649977179
transform 1 0 42044 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_457
timestamp 1649977179
transform 1 0 43148 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_469
timestamp 1649977179
transform 1 0 44252 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_475
timestamp 1649977179
transform 1 0 44804 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_477
timestamp 1649977179
transform 1 0 44988 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_489
timestamp 1649977179
transform 1 0 46092 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_501
timestamp 1649977179
transform 1 0 47196 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_513
timestamp 1649977179
transform 1 0 48300 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_525
timestamp 1649977179
transform 1 0 49404 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_531
timestamp 1649977179
transform 1 0 49956 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_533
timestamp 1649977179
transform 1 0 50140 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_545
timestamp 1649977179
transform 1 0 51244 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_557
timestamp 1649977179
transform 1 0 52348 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_569
timestamp 1649977179
transform 1 0 53452 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_581
timestamp 1649977179
transform 1 0 54556 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_587
timestamp 1649977179
transform 1 0 55108 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_589
timestamp 1649977179
transform 1 0 55292 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_601
timestamp 1649977179
transform 1 0 56396 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_613
timestamp 1649977179
transform 1 0 57500 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_625
timestamp 1649977179
transform 1 0 58604 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_637
timestamp 1649977179
transform 1 0 59708 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_643
timestamp 1649977179
transform 1 0 60260 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_645
timestamp 1649977179
transform 1 0 60444 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_657
timestamp 1649977179
transform 1 0 61548 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_669
timestamp 1649977179
transform 1 0 62652 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_681
timestamp 1649977179
transform 1 0 63756 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_693
timestamp 1649977179
transform 1 0 64860 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_699
timestamp 1649977179
transform 1 0 65412 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_701
timestamp 1649977179
transform 1 0 65596 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_713
timestamp 1649977179
transform 1 0 66700 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_725
timestamp 1649977179
transform 1 0 67804 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_737
timestamp 1649977179
transform 1 0 68908 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_749
timestamp 1649977179
transform 1 0 70012 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_755
timestamp 1649977179
transform 1 0 70564 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_757
timestamp 1649977179
transform 1 0 70748 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_769
timestamp 1649977179
transform 1 0 71852 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_781
timestamp 1649977179
transform 1 0 72956 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_793
timestamp 1649977179
transform 1 0 74060 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_805
timestamp 1649977179
transform 1 0 75164 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_811
timestamp 1649977179
transform 1 0 75716 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_813
timestamp 1649977179
transform 1 0 75900 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_825
timestamp 1649977179
transform 1 0 77004 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_837
timestamp 1649977179
transform 1 0 78108 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_841
timestamp 1649977179
transform 1 0 78476 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_3
timestamp 1649977179
transform 1 0 1380 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_15
timestamp 1649977179
transform 1 0 2484 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_27
timestamp 1649977179
transform 1 0 3588 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_39
timestamp 1649977179
transform 1 0 4692 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_51
timestamp 1649977179
transform 1 0 5796 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1649977179
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_57
timestamp 1649977179
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_69
timestamp 1649977179
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_81
timestamp 1649977179
transform 1 0 8556 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_93
timestamp 1649977179
transform 1 0 9660 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_105
timestamp 1649977179
transform 1 0 10764 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_111
timestamp 1649977179
transform 1 0 11316 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_113
timestamp 1649977179
transform 1 0 11500 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_125
timestamp 1649977179
transform 1 0 12604 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_137
timestamp 1649977179
transform 1 0 13708 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_149
timestamp 1649977179
transform 1 0 14812 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_161
timestamp 1649977179
transform 1 0 15916 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_167
timestamp 1649977179
transform 1 0 16468 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_169
timestamp 1649977179
transform 1 0 16652 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_181
timestamp 1649977179
transform 1 0 17756 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_193
timestamp 1649977179
transform 1 0 18860 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_205
timestamp 1649977179
transform 1 0 19964 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_217
timestamp 1649977179
transform 1 0 21068 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_223
timestamp 1649977179
transform 1 0 21620 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_225
timestamp 1649977179
transform 1 0 21804 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_237
timestamp 1649977179
transform 1 0 22908 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_249
timestamp 1649977179
transform 1 0 24012 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_261
timestamp 1649977179
transform 1 0 25116 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_273
timestamp 1649977179
transform 1 0 26220 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_279
timestamp 1649977179
transform 1 0 26772 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_281
timestamp 1649977179
transform 1 0 26956 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_293
timestamp 1649977179
transform 1 0 28060 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_305
timestamp 1649977179
transform 1 0 29164 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_317
timestamp 1649977179
transform 1 0 30268 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_329
timestamp 1649977179
transform 1 0 31372 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_335
timestamp 1649977179
transform 1 0 31924 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_337
timestamp 1649977179
transform 1 0 32108 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_349
timestamp 1649977179
transform 1 0 33212 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_361
timestamp 1649977179
transform 1 0 34316 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_373
timestamp 1649977179
transform 1 0 35420 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_385
timestamp 1649977179
transform 1 0 36524 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_391
timestamp 1649977179
transform 1 0 37076 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_393
timestamp 1649977179
transform 1 0 37260 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_405
timestamp 1649977179
transform 1 0 38364 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_417
timestamp 1649977179
transform 1 0 39468 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_429
timestamp 1649977179
transform 1 0 40572 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_441
timestamp 1649977179
transform 1 0 41676 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_447
timestamp 1649977179
transform 1 0 42228 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_449
timestamp 1649977179
transform 1 0 42412 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_461
timestamp 1649977179
transform 1 0 43516 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_473
timestamp 1649977179
transform 1 0 44620 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_485
timestamp 1649977179
transform 1 0 45724 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_497
timestamp 1649977179
transform 1 0 46828 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_503
timestamp 1649977179
transform 1 0 47380 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_505
timestamp 1649977179
transform 1 0 47564 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_517
timestamp 1649977179
transform 1 0 48668 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_529
timestamp 1649977179
transform 1 0 49772 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_541
timestamp 1649977179
transform 1 0 50876 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_553
timestamp 1649977179
transform 1 0 51980 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_559
timestamp 1649977179
transform 1 0 52532 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_561
timestamp 1649977179
transform 1 0 52716 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_573
timestamp 1649977179
transform 1 0 53820 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_585
timestamp 1649977179
transform 1 0 54924 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_597
timestamp 1649977179
transform 1 0 56028 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_609
timestamp 1649977179
transform 1 0 57132 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_615
timestamp 1649977179
transform 1 0 57684 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_617
timestamp 1649977179
transform 1 0 57868 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_629
timestamp 1649977179
transform 1 0 58972 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_641
timestamp 1649977179
transform 1 0 60076 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_653
timestamp 1649977179
transform 1 0 61180 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_665
timestamp 1649977179
transform 1 0 62284 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_671
timestamp 1649977179
transform 1 0 62836 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_673
timestamp 1649977179
transform 1 0 63020 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_685
timestamp 1649977179
transform 1 0 64124 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_697
timestamp 1649977179
transform 1 0 65228 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_709
timestamp 1649977179
transform 1 0 66332 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_721
timestamp 1649977179
transform 1 0 67436 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_727
timestamp 1649977179
transform 1 0 67988 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_729
timestamp 1649977179
transform 1 0 68172 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_741
timestamp 1649977179
transform 1 0 69276 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_753
timestamp 1649977179
transform 1 0 70380 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_765
timestamp 1649977179
transform 1 0 71484 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_777
timestamp 1649977179
transform 1 0 72588 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_783
timestamp 1649977179
transform 1 0 73140 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_785
timestamp 1649977179
transform 1 0 73324 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_797
timestamp 1649977179
transform 1 0 74428 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_809
timestamp 1649977179
transform 1 0 75532 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_821
timestamp 1649977179
transform 1 0 76636 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_833
timestamp 1649977179
transform 1 0 77740 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_839
timestamp 1649977179
transform 1 0 78292 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_137_841
timestamp 1649977179
transform 1 0 78476 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1649977179
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1649977179
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1649977179
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1649977179
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_41
timestamp 1649977179
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_53
timestamp 1649977179
transform 1 0 5980 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_57
timestamp 1649977179
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_69
timestamp 1649977179
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1649977179
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_85
timestamp 1649977179
transform 1 0 8924 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_97
timestamp 1649977179
transform 1 0 10028 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_109
timestamp 1649977179
transform 1 0 11132 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_113
timestamp 1649977179
transform 1 0 11500 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_125
timestamp 1649977179
transform 1 0 12604 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_137
timestamp 1649977179
transform 1 0 13708 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_141
timestamp 1649977179
transform 1 0 14076 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_153
timestamp 1649977179
transform 1 0 15180 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_165
timestamp 1649977179
transform 1 0 16284 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_169
timestamp 1649977179
transform 1 0 16652 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_181
timestamp 1649977179
transform 1 0 17756 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_193
timestamp 1649977179
transform 1 0 18860 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_197
timestamp 1649977179
transform 1 0 19228 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_209
timestamp 1649977179
transform 1 0 20332 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_221
timestamp 1649977179
transform 1 0 21436 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_225
timestamp 1649977179
transform 1 0 21804 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_237
timestamp 1649977179
transform 1 0 22908 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_249
timestamp 1649977179
transform 1 0 24012 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_253
timestamp 1649977179
transform 1 0 24380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_265
timestamp 1649977179
transform 1 0 25484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_277
timestamp 1649977179
transform 1 0 26588 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_281
timestamp 1649977179
transform 1 0 26956 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_293
timestamp 1649977179
transform 1 0 28060 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_305
timestamp 1649977179
transform 1 0 29164 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_309
timestamp 1649977179
transform 1 0 29532 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_321
timestamp 1649977179
transform 1 0 30636 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_333
timestamp 1649977179
transform 1 0 31740 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_337
timestamp 1649977179
transform 1 0 32108 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_349
timestamp 1649977179
transform 1 0 33212 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_361
timestamp 1649977179
transform 1 0 34316 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_365
timestamp 1649977179
transform 1 0 34684 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_377
timestamp 1649977179
transform 1 0 35788 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_389
timestamp 1649977179
transform 1 0 36892 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_393
timestamp 1649977179
transform 1 0 37260 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_405
timestamp 1649977179
transform 1 0 38364 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_417
timestamp 1649977179
transform 1 0 39468 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_421
timestamp 1649977179
transform 1 0 39836 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_433
timestamp 1649977179
transform 1 0 40940 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_445
timestamp 1649977179
transform 1 0 42044 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_449
timestamp 1649977179
transform 1 0 42412 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_461
timestamp 1649977179
transform 1 0 43516 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_473
timestamp 1649977179
transform 1 0 44620 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_477
timestamp 1649977179
transform 1 0 44988 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_489
timestamp 1649977179
transform 1 0 46092 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_501
timestamp 1649977179
transform 1 0 47196 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_505
timestamp 1649977179
transform 1 0 47564 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_517
timestamp 1649977179
transform 1 0 48668 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_529
timestamp 1649977179
transform 1 0 49772 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_533
timestamp 1649977179
transform 1 0 50140 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_545
timestamp 1649977179
transform 1 0 51244 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_557
timestamp 1649977179
transform 1 0 52348 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_561
timestamp 1649977179
transform 1 0 52716 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_573
timestamp 1649977179
transform 1 0 53820 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_585
timestamp 1649977179
transform 1 0 54924 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_589
timestamp 1649977179
transform 1 0 55292 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_601
timestamp 1649977179
transform 1 0 56396 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_613
timestamp 1649977179
transform 1 0 57500 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_617
timestamp 1649977179
transform 1 0 57868 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_629
timestamp 1649977179
transform 1 0 58972 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_641
timestamp 1649977179
transform 1 0 60076 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_645
timestamp 1649977179
transform 1 0 60444 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_657
timestamp 1649977179
transform 1 0 61548 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_669
timestamp 1649977179
transform 1 0 62652 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_673
timestamp 1649977179
transform 1 0 63020 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_685
timestamp 1649977179
transform 1 0 64124 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_697
timestamp 1649977179
transform 1 0 65228 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_701
timestamp 1649977179
transform 1 0 65596 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_713
timestamp 1649977179
transform 1 0 66700 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_725
timestamp 1649977179
transform 1 0 67804 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_729
timestamp 1649977179
transform 1 0 68172 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_741
timestamp 1649977179
transform 1 0 69276 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_753
timestamp 1649977179
transform 1 0 70380 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_757
timestamp 1649977179
transform 1 0 70748 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_769
timestamp 1649977179
transform 1 0 71852 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_781
timestamp 1649977179
transform 1 0 72956 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_785
timestamp 1649977179
transform 1 0 73324 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_797
timestamp 1649977179
transform 1 0 74428 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_809
timestamp 1649977179
transform 1 0 75532 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_813
timestamp 1649977179
transform 1 0 75900 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_825
timestamp 1649977179
transform 1 0 77004 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_837
timestamp 1649977179
transform 1 0 78108 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_138_841
timestamp 1649977179
transform 1 0 78476 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 78844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 78844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 78844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 78844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 78844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 78844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 78844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 78844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 78844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 78844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 78844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 78844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 78844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 78844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 78844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 78844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 78844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 78844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 78844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 78844 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 78844 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 78844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 78844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 78844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 78844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 78844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 78844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 78844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 78844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 78844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 78844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 78844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 78844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 78844 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 78844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 78844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 78844 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 78844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 78844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 78844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 78844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 78844 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 78844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 78844 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 78844 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 78844 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 78844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 78844 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 78844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 78844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 78844 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 78844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 78844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 78844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 78844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 78844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 78844 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 78844 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 78844 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 78844 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 78844 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 78844 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 78844 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 78844 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 78844 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 78844 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 78844 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 78844 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 78844 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 78844 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 78844 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 78844 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 78844 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 78844 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 78844 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 78844 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 78844 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 78844 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 78844 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 78844 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 78844 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 78844 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 78844 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 78844 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 78844 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 78844 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 78844 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 78844 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 78844 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 78844 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 78844 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 78844 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 78844 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 78844 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 78844 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 78844 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 78844 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 78844 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 78844 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 78844 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 78844 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 78844 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1649977179
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1649977179
transform -1 0 78844 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1649977179
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1649977179
transform -1 0 78844 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1649977179
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1649977179
transform -1 0 78844 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1649977179
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1649977179
transform -1 0 78844 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1649977179
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1649977179
transform -1 0 78844 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1649977179
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1649977179
transform -1 0 78844 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1649977179
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1649977179
transform -1 0 78844 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1649977179
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1649977179
transform -1 0 78844 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1649977179
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1649977179
transform -1 0 78844 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1649977179
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1649977179
transform -1 0 78844 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1649977179
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1649977179
transform -1 0 78844 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1649977179
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1649977179
transform -1 0 78844 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1649977179
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1649977179
transform -1 0 78844 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1649977179
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1649977179
transform -1 0 78844 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1649977179
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1649977179
transform -1 0 78844 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1649977179
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1649977179
transform -1 0 78844 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1649977179
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1649977179
transform -1 0 78844 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1649977179
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1649977179
transform -1 0 78844 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1649977179
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1649977179
transform -1 0 78844 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1649977179
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1649977179
transform -1 0 78844 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1649977179
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1649977179
transform -1 0 78844 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1649977179
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1649977179
transform -1 0 78844 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1649977179
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1649977179
transform -1 0 78844 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1649977179
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1649977179
transform -1 0 78844 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1649977179
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1649977179
transform -1 0 78844 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1649977179
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1649977179
transform -1 0 78844 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1649977179
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1649977179
transform -1 0 78844 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1649977179
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1649977179
transform -1 0 78844 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1649977179
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1649977179
transform -1 0 78844 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1649977179
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1649977179
transform -1 0 78844 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1649977179
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1649977179
transform -1 0 78844 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1649977179
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1649977179
transform -1 0 78844 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1649977179
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1649977179
transform -1 0 78844 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1649977179
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1649977179
transform -1 0 78844 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1649977179
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1649977179
transform -1 0 78844 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1649977179
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1649977179
transform -1 0 78844 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1649977179
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1649977179
transform -1 0 78844 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 70656 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 73232 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 75808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 78384 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 73232 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 78384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 70656 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 75808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 73232 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 78384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 70656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 75808 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 73232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 78384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 70656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 75808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 73232 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 78384 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 70656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 75808 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 73232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 78384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 70656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 75808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 73232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 78384 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 70656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 75808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 73232 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 78384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 70656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 75808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 73232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 78384 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 70656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 75808 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 73232 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 78384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 70656 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 75808 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 73232 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 78384 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 70656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 75808 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 73232 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 78384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 70656 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 75808 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 73232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 78384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 70656 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 75808 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 73232 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 78384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 70656 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 75808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 73232 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 78384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 70656 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 75808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 73232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 78384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 70656 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 75808 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 73232 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 78384 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 70656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 75808 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 73232 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 78384 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 70656 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 75808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 73232 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 78384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 70656 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 75808 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 73232 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 78384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 70656 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 75808 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 73232 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 78384 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 70656 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 75808 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 73232 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 78384 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 70656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 75808 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 73232 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 78384 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 70656 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 75808 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 73232 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 78384 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 70656 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 75808 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 73232 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 78384 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 70656 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 75808 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 73232 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 78384 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 70656 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 75808 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 73232 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 78384 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 70656 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 75808 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 73232 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 78384 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 70656 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 75808 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 73232 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 78384 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 70656 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 75808 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 73232 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 78384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 70656 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 75808 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 73232 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 78384 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 70656 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 75808 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 73232 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 78384 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 70656 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 75808 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 73232 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 78384 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 70656 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 75808 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 73232 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 78384 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 70656 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 75808 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 73232 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 78384 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 70656 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 75808 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 73232 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 78384 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1649977179
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1649977179
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1649977179
transform 1 0 70656 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1649977179
transform 1 0 75808 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1649977179
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1649977179
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1649977179
transform 1 0 73232 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1649977179
transform 1 0 78384 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1649977179
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1649977179
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1649977179
transform 1 0 70656 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1649977179
transform 1 0 75808 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1649977179
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1649977179
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1649977179
transform 1 0 73232 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1649977179
transform 1 0 78384 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1649977179
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1649977179
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1649977179
transform 1 0 70656 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1649977179
transform 1 0 75808 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1649977179
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1649977179
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1649977179
transform 1 0 73232 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1649977179
transform 1 0 78384 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1649977179
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1649977179
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1649977179
transform 1 0 70656 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1649977179
transform 1 0 75808 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1649977179
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1649977179
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1649977179
transform 1 0 73232 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1649977179
transform 1 0 78384 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1649977179
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1649977179
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1649977179
transform 1 0 70656 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1649977179
transform 1 0 75808 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1649977179
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1649977179
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1649977179
transform 1 0 73232 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1649977179
transform 1 0 78384 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1649977179
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1649977179
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1649977179
transform 1 0 70656 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1649977179
transform 1 0 75808 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1649977179
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1649977179
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1649977179
transform 1 0 73232 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1649977179
transform 1 0 78384 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1649977179
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1649977179
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1649977179
transform 1 0 70656 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1649977179
transform 1 0 75808 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1649977179
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1649977179
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1649977179
transform 1 0 73232 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1649977179
transform 1 0 78384 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1556
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1557
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1558
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1559
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1560
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1561
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1562
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1563
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1564
timestamp 1649977179
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1565
timestamp 1649977179
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1566
timestamp 1649977179
transform 1 0 70656 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1567
timestamp 1649977179
transform 1 0 75808 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1568
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1569
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1570
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1571
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1572
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1573
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1574
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1575
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1576
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1577
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1578
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1579
timestamp 1649977179
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1580
timestamp 1649977179
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1581
timestamp 1649977179
transform 1 0 73232 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1582
timestamp 1649977179
transform 1 0 78384 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1583
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1584
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1585
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1586
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1587
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1588
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1589
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1590
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1591
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1592
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1593
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1594
timestamp 1649977179
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1595
timestamp 1649977179
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1596
timestamp 1649977179
transform 1 0 70656 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1597
timestamp 1649977179
transform 1 0 75808 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1598
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1599
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1600
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1601
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1602
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1603
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1604
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1605
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1606
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1607
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1608
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1609
timestamp 1649977179
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1610
timestamp 1649977179
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1611
timestamp 1649977179
transform 1 0 73232 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1612
timestamp 1649977179
transform 1 0 78384 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1613
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1614
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1615
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1616
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1617
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1618
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1619
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1620
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1621
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1622
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1623
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1624
timestamp 1649977179
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1625
timestamp 1649977179
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1626
timestamp 1649977179
transform 1 0 70656 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1627
timestamp 1649977179
transform 1 0 75808 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1628
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1629
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1630
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1631
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1632
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1633
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1634
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1635
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1636
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1637
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1638
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1639
timestamp 1649977179
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1640
timestamp 1649977179
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1641
timestamp 1649977179
transform 1 0 73232 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1642
timestamp 1649977179
transform 1 0 78384 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1643
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1644
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1645
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1646
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1647
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1648
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1649
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1650
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1651
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1652
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1653
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1654
timestamp 1649977179
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1655
timestamp 1649977179
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1656
timestamp 1649977179
transform 1 0 70656 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1657
timestamp 1649977179
transform 1 0 75808 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1658
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1659
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1660
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1661
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1662
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1663
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1664
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1665
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1666
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1667
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1668
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1669
timestamp 1649977179
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1670
timestamp 1649977179
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1671
timestamp 1649977179
transform 1 0 73232 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1672
timestamp 1649977179
transform 1 0 78384 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1673
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1674
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1675
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1676
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1677
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1678
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1679
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1680
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1681
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1682
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1683
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1684
timestamp 1649977179
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1685
timestamp 1649977179
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1686
timestamp 1649977179
transform 1 0 70656 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1687
timestamp 1649977179
transform 1 0 75808 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1688
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1689
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1690
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1691
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1692
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1693
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1694
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1695
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1696
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1697
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1698
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1699
timestamp 1649977179
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1700
timestamp 1649977179
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1701
timestamp 1649977179
transform 1 0 73232 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1702
timestamp 1649977179
transform 1 0 78384 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1703
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1704
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1705
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1706
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1707
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1708
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1709
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1710
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1711
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1712
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1713
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1714
timestamp 1649977179
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1715
timestamp 1649977179
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1716
timestamp 1649977179
transform 1 0 70656 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1717
timestamp 1649977179
transform 1 0 75808 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1718
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1719
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1720
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1721
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1722
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1723
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1724
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1725
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1726
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1727
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1728
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1729
timestamp 1649977179
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1730
timestamp 1649977179
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1731
timestamp 1649977179
transform 1 0 73232 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1732
timestamp 1649977179
transform 1 0 78384 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1733
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1734
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1735
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1736
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1737
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1738
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1739
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1740
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1741
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1742
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1743
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1744
timestamp 1649977179
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1745
timestamp 1649977179
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1746
timestamp 1649977179
transform 1 0 70656 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1747
timestamp 1649977179
transform 1 0 75808 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1748
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1749
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1750
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1751
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1752
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1753
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1754
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1755
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1756
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1757
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1758
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1759
timestamp 1649977179
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1760
timestamp 1649977179
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1761
timestamp 1649977179
transform 1 0 73232 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1762
timestamp 1649977179
transform 1 0 78384 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1763
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1764
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1765
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1766
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1767
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1768
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1769
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1770
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1771
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1772
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1773
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1774
timestamp 1649977179
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1775
timestamp 1649977179
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1776
timestamp 1649977179
transform 1 0 70656 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1777
timestamp 1649977179
transform 1 0 75808 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1778
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1779
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1780
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1781
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1782
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1783
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1784
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1785
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1786
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1787
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1788
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1789
timestamp 1649977179
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1790
timestamp 1649977179
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1791
timestamp 1649977179
transform 1 0 73232 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1792
timestamp 1649977179
transform 1 0 78384 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1793
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1794
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1795
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1796
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1797
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1798
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1799
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1800
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1801
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1802
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1803
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1804
timestamp 1649977179
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1805
timestamp 1649977179
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1806
timestamp 1649977179
transform 1 0 70656 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1807
timestamp 1649977179
transform 1 0 75808 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1808
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1809
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1810
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1811
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1812
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1813
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1814
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1815
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1816
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1817
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1818
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1819
timestamp 1649977179
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1820
timestamp 1649977179
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1821
timestamp 1649977179
transform 1 0 73232 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1822
timestamp 1649977179
transform 1 0 78384 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1823
timestamp 1649977179
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1824
timestamp 1649977179
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1825
timestamp 1649977179
transform 1 0 13984 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1826
timestamp 1649977179
transform 1 0 19136 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1827
timestamp 1649977179
transform 1 0 24288 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1828
timestamp 1649977179
transform 1 0 29440 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1829
timestamp 1649977179
transform 1 0 34592 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1830
timestamp 1649977179
transform 1 0 39744 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1831
timestamp 1649977179
transform 1 0 44896 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1832
timestamp 1649977179
transform 1 0 50048 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1833
timestamp 1649977179
transform 1 0 55200 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1834
timestamp 1649977179
transform 1 0 60352 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1835
timestamp 1649977179
transform 1 0 65504 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1836
timestamp 1649977179
transform 1 0 70656 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1837
timestamp 1649977179
transform 1 0 75808 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1838
timestamp 1649977179
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1839
timestamp 1649977179
transform 1 0 11408 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1840
timestamp 1649977179
transform 1 0 16560 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1841
timestamp 1649977179
transform 1 0 21712 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1842
timestamp 1649977179
transform 1 0 26864 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1843
timestamp 1649977179
transform 1 0 32016 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1844
timestamp 1649977179
transform 1 0 37168 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1845
timestamp 1649977179
transform 1 0 42320 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1846
timestamp 1649977179
transform 1 0 47472 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1847
timestamp 1649977179
transform 1 0 52624 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1848
timestamp 1649977179
transform 1 0 57776 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1849
timestamp 1649977179
transform 1 0 62928 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1850
timestamp 1649977179
transform 1 0 68080 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1851
timestamp 1649977179
transform 1 0 73232 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1852
timestamp 1649977179
transform 1 0 78384 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1853
timestamp 1649977179
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1854
timestamp 1649977179
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1855
timestamp 1649977179
transform 1 0 13984 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1856
timestamp 1649977179
transform 1 0 19136 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1857
timestamp 1649977179
transform 1 0 24288 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1858
timestamp 1649977179
transform 1 0 29440 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1859
timestamp 1649977179
transform 1 0 34592 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1860
timestamp 1649977179
transform 1 0 39744 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1861
timestamp 1649977179
transform 1 0 44896 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1862
timestamp 1649977179
transform 1 0 50048 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1863
timestamp 1649977179
transform 1 0 55200 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1864
timestamp 1649977179
transform 1 0 60352 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1865
timestamp 1649977179
transform 1 0 65504 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1866
timestamp 1649977179
transform 1 0 70656 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1867
timestamp 1649977179
transform 1 0 75808 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1868
timestamp 1649977179
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1869
timestamp 1649977179
transform 1 0 11408 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1870
timestamp 1649977179
transform 1 0 16560 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1871
timestamp 1649977179
transform 1 0 21712 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1872
timestamp 1649977179
transform 1 0 26864 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1873
timestamp 1649977179
transform 1 0 32016 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1874
timestamp 1649977179
transform 1 0 37168 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1875
timestamp 1649977179
transform 1 0 42320 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1876
timestamp 1649977179
transform 1 0 47472 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1877
timestamp 1649977179
transform 1 0 52624 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1878
timestamp 1649977179
transform 1 0 57776 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1879
timestamp 1649977179
transform 1 0 62928 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1880
timestamp 1649977179
transform 1 0 68080 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1881
timestamp 1649977179
transform 1 0 73232 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1882
timestamp 1649977179
transform 1 0 78384 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1883
timestamp 1649977179
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1884
timestamp 1649977179
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1885
timestamp 1649977179
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1886
timestamp 1649977179
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1887
timestamp 1649977179
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1888
timestamp 1649977179
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1889
timestamp 1649977179
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1890
timestamp 1649977179
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1891
timestamp 1649977179
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1892
timestamp 1649977179
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1893
timestamp 1649977179
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1894
timestamp 1649977179
transform 1 0 60352 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1895
timestamp 1649977179
transform 1 0 65504 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1896
timestamp 1649977179
transform 1 0 70656 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1897
timestamp 1649977179
transform 1 0 75808 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1898
timestamp 1649977179
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1899
timestamp 1649977179
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1900
timestamp 1649977179
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1901
timestamp 1649977179
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1902
timestamp 1649977179
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1903
timestamp 1649977179
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1904
timestamp 1649977179
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1905
timestamp 1649977179
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1906
timestamp 1649977179
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1907
timestamp 1649977179
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1908
timestamp 1649977179
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1909
timestamp 1649977179
transform 1 0 62928 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1910
timestamp 1649977179
transform 1 0 68080 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1911
timestamp 1649977179
transform 1 0 73232 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1912
timestamp 1649977179
transform 1 0 78384 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1913
timestamp 1649977179
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1914
timestamp 1649977179
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1915
timestamp 1649977179
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1916
timestamp 1649977179
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1917
timestamp 1649977179
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1918
timestamp 1649977179
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1919
timestamp 1649977179
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1920
timestamp 1649977179
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1921
timestamp 1649977179
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1922
timestamp 1649977179
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1923
timestamp 1649977179
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1924
timestamp 1649977179
transform 1 0 60352 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1925
timestamp 1649977179
transform 1 0 65504 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1926
timestamp 1649977179
transform 1 0 70656 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1927
timestamp 1649977179
transform 1 0 75808 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1928
timestamp 1649977179
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1929
timestamp 1649977179
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1930
timestamp 1649977179
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1931
timestamp 1649977179
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1932
timestamp 1649977179
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1933
timestamp 1649977179
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1934
timestamp 1649977179
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1935
timestamp 1649977179
transform 1 0 42320 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1936
timestamp 1649977179
transform 1 0 47472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1937
timestamp 1649977179
transform 1 0 52624 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1938
timestamp 1649977179
transform 1 0 57776 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1939
timestamp 1649977179
transform 1 0 62928 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1940
timestamp 1649977179
transform 1 0 68080 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1941
timestamp 1649977179
transform 1 0 73232 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1942
timestamp 1649977179
transform 1 0 78384 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1943
timestamp 1649977179
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1944
timestamp 1649977179
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1945
timestamp 1649977179
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1946
timestamp 1649977179
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1947
timestamp 1649977179
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1948
timestamp 1649977179
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1949
timestamp 1649977179
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1950
timestamp 1649977179
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1951
timestamp 1649977179
transform 1 0 44896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1952
timestamp 1649977179
transform 1 0 50048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1953
timestamp 1649977179
transform 1 0 55200 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1954
timestamp 1649977179
transform 1 0 60352 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1955
timestamp 1649977179
transform 1 0 65504 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1956
timestamp 1649977179
transform 1 0 70656 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1957
timestamp 1649977179
transform 1 0 75808 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1958
timestamp 1649977179
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1959
timestamp 1649977179
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1960
timestamp 1649977179
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1961
timestamp 1649977179
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1962
timestamp 1649977179
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1963
timestamp 1649977179
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1964
timestamp 1649977179
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1965
timestamp 1649977179
transform 1 0 42320 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1966
timestamp 1649977179
transform 1 0 47472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1967
timestamp 1649977179
transform 1 0 52624 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1968
timestamp 1649977179
transform 1 0 57776 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1969
timestamp 1649977179
transform 1 0 62928 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1970
timestamp 1649977179
transform 1 0 68080 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1971
timestamp 1649977179
transform 1 0 73232 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1972
timestamp 1649977179
transform 1 0 78384 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1973
timestamp 1649977179
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1974
timestamp 1649977179
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1975
timestamp 1649977179
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1976
timestamp 1649977179
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1977
timestamp 1649977179
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1978
timestamp 1649977179
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1979
timestamp 1649977179
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1980
timestamp 1649977179
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1981
timestamp 1649977179
transform 1 0 44896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1982
timestamp 1649977179
transform 1 0 50048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1983
timestamp 1649977179
transform 1 0 55200 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1984
timestamp 1649977179
transform 1 0 60352 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1985
timestamp 1649977179
transform 1 0 65504 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1986
timestamp 1649977179
transform 1 0 70656 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1987
timestamp 1649977179
transform 1 0 75808 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1988
timestamp 1649977179
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1989
timestamp 1649977179
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1990
timestamp 1649977179
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1991
timestamp 1649977179
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1992
timestamp 1649977179
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1993
timestamp 1649977179
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1994
timestamp 1649977179
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1995
timestamp 1649977179
transform 1 0 42320 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1996
timestamp 1649977179
transform 1 0 47472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1997
timestamp 1649977179
transform 1 0 52624 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1998
timestamp 1649977179
transform 1 0 57776 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1999
timestamp 1649977179
transform 1 0 62928 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2000
timestamp 1649977179
transform 1 0 68080 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2001
timestamp 1649977179
transform 1 0 73232 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2002
timestamp 1649977179
transform 1 0 78384 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2003
timestamp 1649977179
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2004
timestamp 1649977179
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2005
timestamp 1649977179
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2006
timestamp 1649977179
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2007
timestamp 1649977179
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2008
timestamp 1649977179
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2009
timestamp 1649977179
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2010
timestamp 1649977179
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2011
timestamp 1649977179
transform 1 0 44896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2012
timestamp 1649977179
transform 1 0 50048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2013
timestamp 1649977179
transform 1 0 55200 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2014
timestamp 1649977179
transform 1 0 60352 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2015
timestamp 1649977179
transform 1 0 65504 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2016
timestamp 1649977179
transform 1 0 70656 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2017
timestamp 1649977179
transform 1 0 75808 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2018
timestamp 1649977179
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2019
timestamp 1649977179
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2020
timestamp 1649977179
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2021
timestamp 1649977179
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2022
timestamp 1649977179
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2023
timestamp 1649977179
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2024
timestamp 1649977179
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2025
timestamp 1649977179
transform 1 0 42320 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2026
timestamp 1649977179
transform 1 0 47472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2027
timestamp 1649977179
transform 1 0 52624 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2028
timestamp 1649977179
transform 1 0 57776 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2029
timestamp 1649977179
transform 1 0 62928 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2030
timestamp 1649977179
transform 1 0 68080 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2031
timestamp 1649977179
transform 1 0 73232 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2032
timestamp 1649977179
transform 1 0 78384 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2033
timestamp 1649977179
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2034
timestamp 1649977179
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2035
timestamp 1649977179
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2036
timestamp 1649977179
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2037
timestamp 1649977179
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2038
timestamp 1649977179
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2039
timestamp 1649977179
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2040
timestamp 1649977179
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2041
timestamp 1649977179
transform 1 0 44896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2042
timestamp 1649977179
transform 1 0 50048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2043
timestamp 1649977179
transform 1 0 55200 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2044
timestamp 1649977179
transform 1 0 60352 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2045
timestamp 1649977179
transform 1 0 65504 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2046
timestamp 1649977179
transform 1 0 70656 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2047
timestamp 1649977179
transform 1 0 75808 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2048
timestamp 1649977179
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2049
timestamp 1649977179
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2050
timestamp 1649977179
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2051
timestamp 1649977179
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2052
timestamp 1649977179
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2053
timestamp 1649977179
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2054
timestamp 1649977179
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2055
timestamp 1649977179
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2056
timestamp 1649977179
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2057
timestamp 1649977179
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2058
timestamp 1649977179
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2059
timestamp 1649977179
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2060
timestamp 1649977179
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2061
timestamp 1649977179
transform 1 0 73232 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2062
timestamp 1649977179
transform 1 0 78384 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2063
timestamp 1649977179
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2064
timestamp 1649977179
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2065
timestamp 1649977179
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2066
timestamp 1649977179
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2067
timestamp 1649977179
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2068
timestamp 1649977179
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2069
timestamp 1649977179
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2070
timestamp 1649977179
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2071
timestamp 1649977179
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2072
timestamp 1649977179
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2073
timestamp 1649977179
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2074
timestamp 1649977179
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2075
timestamp 1649977179
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2076
timestamp 1649977179
transform 1 0 70656 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2077
timestamp 1649977179
transform 1 0 75808 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2078
timestamp 1649977179
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2079
timestamp 1649977179
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2080
timestamp 1649977179
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2081
timestamp 1649977179
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2082
timestamp 1649977179
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2083
timestamp 1649977179
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2084
timestamp 1649977179
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2085
timestamp 1649977179
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2086
timestamp 1649977179
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2087
timestamp 1649977179
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2088
timestamp 1649977179
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2089
timestamp 1649977179
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2090
timestamp 1649977179
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2091
timestamp 1649977179
transform 1 0 73232 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2092
timestamp 1649977179
transform 1 0 78384 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2093
timestamp 1649977179
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2094
timestamp 1649977179
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2095
timestamp 1649977179
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2096
timestamp 1649977179
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2097
timestamp 1649977179
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2098
timestamp 1649977179
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2099
timestamp 1649977179
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2100
timestamp 1649977179
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2101
timestamp 1649977179
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2102
timestamp 1649977179
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2103
timestamp 1649977179
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2104
timestamp 1649977179
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2105
timestamp 1649977179
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2106
timestamp 1649977179
transform 1 0 70656 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2107
timestamp 1649977179
transform 1 0 75808 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2108
timestamp 1649977179
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2109
timestamp 1649977179
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2110
timestamp 1649977179
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2111
timestamp 1649977179
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2112
timestamp 1649977179
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2113
timestamp 1649977179
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2114
timestamp 1649977179
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2115
timestamp 1649977179
transform 1 0 42320 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2116
timestamp 1649977179
transform 1 0 47472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2117
timestamp 1649977179
transform 1 0 52624 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2118
timestamp 1649977179
transform 1 0 57776 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2119
timestamp 1649977179
transform 1 0 62928 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2120
timestamp 1649977179
transform 1 0 68080 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2121
timestamp 1649977179
transform 1 0 73232 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2122
timestamp 1649977179
transform 1 0 78384 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2123
timestamp 1649977179
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2124
timestamp 1649977179
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2125
timestamp 1649977179
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2126
timestamp 1649977179
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2127
timestamp 1649977179
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2128
timestamp 1649977179
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2129
timestamp 1649977179
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2130
timestamp 1649977179
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2131
timestamp 1649977179
transform 1 0 44896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2132
timestamp 1649977179
transform 1 0 50048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2133
timestamp 1649977179
transform 1 0 55200 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2134
timestamp 1649977179
transform 1 0 60352 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2135
timestamp 1649977179
transform 1 0 65504 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2136
timestamp 1649977179
transform 1 0 70656 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2137
timestamp 1649977179
transform 1 0 75808 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2138
timestamp 1649977179
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2139
timestamp 1649977179
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2140
timestamp 1649977179
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2141
timestamp 1649977179
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2142
timestamp 1649977179
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2143
timestamp 1649977179
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2144
timestamp 1649977179
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2145
timestamp 1649977179
transform 1 0 42320 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2146
timestamp 1649977179
transform 1 0 47472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2147
timestamp 1649977179
transform 1 0 52624 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2148
timestamp 1649977179
transform 1 0 57776 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2149
timestamp 1649977179
transform 1 0 62928 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2150
timestamp 1649977179
transform 1 0 68080 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2151
timestamp 1649977179
transform 1 0 73232 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2152
timestamp 1649977179
transform 1 0 78384 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2153
timestamp 1649977179
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2154
timestamp 1649977179
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2155
timestamp 1649977179
transform 1 0 13984 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2156
timestamp 1649977179
transform 1 0 19136 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2157
timestamp 1649977179
transform 1 0 24288 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2158
timestamp 1649977179
transform 1 0 29440 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2159
timestamp 1649977179
transform 1 0 34592 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2160
timestamp 1649977179
transform 1 0 39744 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2161
timestamp 1649977179
transform 1 0 44896 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2162
timestamp 1649977179
transform 1 0 50048 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2163
timestamp 1649977179
transform 1 0 55200 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2164
timestamp 1649977179
transform 1 0 60352 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2165
timestamp 1649977179
transform 1 0 65504 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2166
timestamp 1649977179
transform 1 0 70656 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2167
timestamp 1649977179
transform 1 0 75808 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2168
timestamp 1649977179
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2169
timestamp 1649977179
transform 1 0 11408 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2170
timestamp 1649977179
transform 1 0 16560 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2171
timestamp 1649977179
transform 1 0 21712 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2172
timestamp 1649977179
transform 1 0 26864 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2173
timestamp 1649977179
transform 1 0 32016 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2174
timestamp 1649977179
transform 1 0 37168 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2175
timestamp 1649977179
transform 1 0 42320 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2176
timestamp 1649977179
transform 1 0 47472 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2177
timestamp 1649977179
transform 1 0 52624 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2178
timestamp 1649977179
transform 1 0 57776 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2179
timestamp 1649977179
transform 1 0 62928 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2180
timestamp 1649977179
transform 1 0 68080 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2181
timestamp 1649977179
transform 1 0 73232 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2182
timestamp 1649977179
transform 1 0 78384 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2183
timestamp 1649977179
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2184
timestamp 1649977179
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2185
timestamp 1649977179
transform 1 0 13984 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2186
timestamp 1649977179
transform 1 0 19136 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2187
timestamp 1649977179
transform 1 0 24288 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2188
timestamp 1649977179
transform 1 0 29440 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2189
timestamp 1649977179
transform 1 0 34592 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2190
timestamp 1649977179
transform 1 0 39744 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2191
timestamp 1649977179
transform 1 0 44896 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2192
timestamp 1649977179
transform 1 0 50048 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2193
timestamp 1649977179
transform 1 0 55200 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2194
timestamp 1649977179
transform 1 0 60352 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2195
timestamp 1649977179
transform 1 0 65504 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2196
timestamp 1649977179
transform 1 0 70656 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2197
timestamp 1649977179
transform 1 0 75808 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2198
timestamp 1649977179
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2199
timestamp 1649977179
transform 1 0 11408 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2200
timestamp 1649977179
transform 1 0 16560 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2201
timestamp 1649977179
transform 1 0 21712 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2202
timestamp 1649977179
transform 1 0 26864 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2203
timestamp 1649977179
transform 1 0 32016 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2204
timestamp 1649977179
transform 1 0 37168 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2205
timestamp 1649977179
transform 1 0 42320 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2206
timestamp 1649977179
transform 1 0 47472 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2207
timestamp 1649977179
transform 1 0 52624 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2208
timestamp 1649977179
transform 1 0 57776 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2209
timestamp 1649977179
transform 1 0 62928 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2210
timestamp 1649977179
transform 1 0 68080 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2211
timestamp 1649977179
transform 1 0 73232 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2212
timestamp 1649977179
transform 1 0 78384 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2213
timestamp 1649977179
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2214
timestamp 1649977179
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2215
timestamp 1649977179
transform 1 0 13984 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2216
timestamp 1649977179
transform 1 0 19136 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2217
timestamp 1649977179
transform 1 0 24288 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2218
timestamp 1649977179
transform 1 0 29440 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2219
timestamp 1649977179
transform 1 0 34592 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2220
timestamp 1649977179
transform 1 0 39744 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2221
timestamp 1649977179
transform 1 0 44896 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2222
timestamp 1649977179
transform 1 0 50048 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2223
timestamp 1649977179
transform 1 0 55200 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2224
timestamp 1649977179
transform 1 0 60352 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2225
timestamp 1649977179
transform 1 0 65504 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2226
timestamp 1649977179
transform 1 0 70656 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2227
timestamp 1649977179
transform 1 0 75808 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2228
timestamp 1649977179
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2229
timestamp 1649977179
transform 1 0 11408 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2230
timestamp 1649977179
transform 1 0 16560 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2231
timestamp 1649977179
transform 1 0 21712 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2232
timestamp 1649977179
transform 1 0 26864 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2233
timestamp 1649977179
transform 1 0 32016 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2234
timestamp 1649977179
transform 1 0 37168 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2235
timestamp 1649977179
transform 1 0 42320 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2236
timestamp 1649977179
transform 1 0 47472 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2237
timestamp 1649977179
transform 1 0 52624 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2238
timestamp 1649977179
transform 1 0 57776 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2239
timestamp 1649977179
transform 1 0 62928 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2240
timestamp 1649977179
transform 1 0 68080 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2241
timestamp 1649977179
transform 1 0 73232 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2242
timestamp 1649977179
transform 1 0 78384 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2243
timestamp 1649977179
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2244
timestamp 1649977179
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2245
timestamp 1649977179
transform 1 0 13984 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2246
timestamp 1649977179
transform 1 0 19136 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2247
timestamp 1649977179
transform 1 0 24288 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2248
timestamp 1649977179
transform 1 0 29440 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2249
timestamp 1649977179
transform 1 0 34592 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2250
timestamp 1649977179
transform 1 0 39744 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2251
timestamp 1649977179
transform 1 0 44896 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2252
timestamp 1649977179
transform 1 0 50048 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2253
timestamp 1649977179
transform 1 0 55200 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2254
timestamp 1649977179
transform 1 0 60352 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2255
timestamp 1649977179
transform 1 0 65504 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2256
timestamp 1649977179
transform 1 0 70656 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2257
timestamp 1649977179
transform 1 0 75808 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2258
timestamp 1649977179
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2259
timestamp 1649977179
transform 1 0 11408 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2260
timestamp 1649977179
transform 1 0 16560 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2261
timestamp 1649977179
transform 1 0 21712 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2262
timestamp 1649977179
transform 1 0 26864 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2263
timestamp 1649977179
transform 1 0 32016 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2264
timestamp 1649977179
transform 1 0 37168 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2265
timestamp 1649977179
transform 1 0 42320 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2266
timestamp 1649977179
transform 1 0 47472 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2267
timestamp 1649977179
transform 1 0 52624 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2268
timestamp 1649977179
transform 1 0 57776 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2269
timestamp 1649977179
transform 1 0 62928 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2270
timestamp 1649977179
transform 1 0 68080 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2271
timestamp 1649977179
transform 1 0 73232 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2272
timestamp 1649977179
transform 1 0 78384 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2273
timestamp 1649977179
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2274
timestamp 1649977179
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2275
timestamp 1649977179
transform 1 0 13984 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2276
timestamp 1649977179
transform 1 0 19136 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2277
timestamp 1649977179
transform 1 0 24288 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2278
timestamp 1649977179
transform 1 0 29440 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2279
timestamp 1649977179
transform 1 0 34592 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2280
timestamp 1649977179
transform 1 0 39744 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2281
timestamp 1649977179
transform 1 0 44896 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2282
timestamp 1649977179
transform 1 0 50048 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2283
timestamp 1649977179
transform 1 0 55200 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2284
timestamp 1649977179
transform 1 0 60352 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2285
timestamp 1649977179
transform 1 0 65504 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2286
timestamp 1649977179
transform 1 0 70656 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2287
timestamp 1649977179
transform 1 0 75808 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2288
timestamp 1649977179
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2289
timestamp 1649977179
transform 1 0 11408 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2290
timestamp 1649977179
transform 1 0 16560 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2291
timestamp 1649977179
transform 1 0 21712 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2292
timestamp 1649977179
transform 1 0 26864 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2293
timestamp 1649977179
transform 1 0 32016 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2294
timestamp 1649977179
transform 1 0 37168 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2295
timestamp 1649977179
transform 1 0 42320 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2296
timestamp 1649977179
transform 1 0 47472 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2297
timestamp 1649977179
transform 1 0 52624 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2298
timestamp 1649977179
transform 1 0 57776 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2299
timestamp 1649977179
transform 1 0 62928 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2300
timestamp 1649977179
transform 1 0 68080 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2301
timestamp 1649977179
transform 1 0 73232 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2302
timestamp 1649977179
transform 1 0 78384 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2303
timestamp 1649977179
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2304
timestamp 1649977179
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2305
timestamp 1649977179
transform 1 0 13984 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2306
timestamp 1649977179
transform 1 0 19136 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2307
timestamp 1649977179
transform 1 0 24288 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2308
timestamp 1649977179
transform 1 0 29440 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2309
timestamp 1649977179
transform 1 0 34592 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2310
timestamp 1649977179
transform 1 0 39744 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2311
timestamp 1649977179
transform 1 0 44896 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2312
timestamp 1649977179
transform 1 0 50048 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2313
timestamp 1649977179
transform 1 0 55200 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2314
timestamp 1649977179
transform 1 0 60352 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2315
timestamp 1649977179
transform 1 0 65504 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2316
timestamp 1649977179
transform 1 0 70656 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2317
timestamp 1649977179
transform 1 0 75808 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2318
timestamp 1649977179
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2319
timestamp 1649977179
transform 1 0 11408 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2320
timestamp 1649977179
transform 1 0 16560 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2321
timestamp 1649977179
transform 1 0 21712 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2322
timestamp 1649977179
transform 1 0 26864 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2323
timestamp 1649977179
transform 1 0 32016 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2324
timestamp 1649977179
transform 1 0 37168 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2325
timestamp 1649977179
transform 1 0 42320 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2326
timestamp 1649977179
transform 1 0 47472 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2327
timestamp 1649977179
transform 1 0 52624 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2328
timestamp 1649977179
transform 1 0 57776 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2329
timestamp 1649977179
transform 1 0 62928 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2330
timestamp 1649977179
transform 1 0 68080 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2331
timestamp 1649977179
transform 1 0 73232 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2332
timestamp 1649977179
transform 1 0 78384 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2333
timestamp 1649977179
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2334
timestamp 1649977179
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2335
timestamp 1649977179
transform 1 0 13984 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2336
timestamp 1649977179
transform 1 0 19136 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2337
timestamp 1649977179
transform 1 0 24288 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2338
timestamp 1649977179
transform 1 0 29440 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2339
timestamp 1649977179
transform 1 0 34592 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2340
timestamp 1649977179
transform 1 0 39744 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2341
timestamp 1649977179
transform 1 0 44896 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2342
timestamp 1649977179
transform 1 0 50048 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2343
timestamp 1649977179
transform 1 0 55200 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2344
timestamp 1649977179
transform 1 0 60352 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2345
timestamp 1649977179
transform 1 0 65504 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2346
timestamp 1649977179
transform 1 0 70656 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2347
timestamp 1649977179
transform 1 0 75808 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2348
timestamp 1649977179
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2349
timestamp 1649977179
transform 1 0 11408 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2350
timestamp 1649977179
transform 1 0 16560 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2351
timestamp 1649977179
transform 1 0 21712 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2352
timestamp 1649977179
transform 1 0 26864 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2353
timestamp 1649977179
transform 1 0 32016 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2354
timestamp 1649977179
transform 1 0 37168 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2355
timestamp 1649977179
transform 1 0 42320 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2356
timestamp 1649977179
transform 1 0 47472 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2357
timestamp 1649977179
transform 1 0 52624 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2358
timestamp 1649977179
transform 1 0 57776 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2359
timestamp 1649977179
transform 1 0 62928 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2360
timestamp 1649977179
transform 1 0 68080 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2361
timestamp 1649977179
transform 1 0 73232 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2362
timestamp 1649977179
transform 1 0 78384 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2363
timestamp 1649977179
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2364
timestamp 1649977179
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2365
timestamp 1649977179
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2366
timestamp 1649977179
transform 1 0 11408 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2367
timestamp 1649977179
transform 1 0 13984 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2368
timestamp 1649977179
transform 1 0 16560 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2369
timestamp 1649977179
transform 1 0 19136 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2370
timestamp 1649977179
transform 1 0 21712 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2371
timestamp 1649977179
transform 1 0 24288 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2372
timestamp 1649977179
transform 1 0 26864 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2373
timestamp 1649977179
transform 1 0 29440 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2374
timestamp 1649977179
transform 1 0 32016 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2375
timestamp 1649977179
transform 1 0 34592 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2376
timestamp 1649977179
transform 1 0 37168 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2377
timestamp 1649977179
transform 1 0 39744 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2378
timestamp 1649977179
transform 1 0 42320 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2379
timestamp 1649977179
transform 1 0 44896 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2380
timestamp 1649977179
transform 1 0 47472 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2381
timestamp 1649977179
transform 1 0 50048 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2382
timestamp 1649977179
transform 1 0 52624 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2383
timestamp 1649977179
transform 1 0 55200 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2384
timestamp 1649977179
transform 1 0 57776 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2385
timestamp 1649977179
transform 1 0 60352 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2386
timestamp 1649977179
transform 1 0 62928 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2387
timestamp 1649977179
transform 1 0 65504 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2388
timestamp 1649977179
transform 1 0 68080 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2389
timestamp 1649977179
transform 1 0 70656 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2390
timestamp 1649977179
transform 1 0 73232 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2391
timestamp 1649977179
transform 1 0 75808 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_2392
timestamp 1649977179
transform 1 0 78384 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__or4_1  _029_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31096 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _030_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32200 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _031_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 31648 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _032_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _033_
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _034_
timestamp 1649977179
transform 1 0 27048 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _035_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27232 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_2  _036_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 41216 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _037_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 60720 0 1 55488
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _038_
timestamp 1649977179
transform 1 0 53176 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _039_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 41492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _040_
timestamp 1649977179
transform 1 0 61180 0 -1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _041_
timestamp 1649977179
transform 1 0 52900 0 1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _042_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 52808 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _043_
timestamp 1649977179
transform 1 0 50140 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _044_
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _045_
timestamp 1649977179
transform 1 0 50324 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _046_
timestamp 1649977179
transform 1 0 50784 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _047_
timestamp 1649977179
transform 1 0 53360 0 1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _048_
timestamp 1649977179
transform 1 0 53084 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _049_
timestamp 1649977179
transform 1 0 51796 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _050_
timestamp 1649977179
transform -1 0 55108 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _051_
timestamp 1649977179
transform 1 0 52992 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _052_
timestamp 1649977179
transform 1 0 51520 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _053_
timestamp 1649977179
transform 1 0 54096 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _054_
timestamp 1649977179
transform 1 0 57592 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _055_
timestamp 1649977179
transform 1 0 56304 0 1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _056_
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _057_
timestamp 1649977179
transform 1 0 56212 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _058_
timestamp 1649977179
transform 1 0 56488 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _059_
timestamp 1649977179
transform 1 0 57592 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _060_
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _061_
timestamp 1649977179
transform -1 0 60812 0 -1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _062_
timestamp 1649977179
transform 1 0 60444 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _063_
timestamp 1649977179
transform 1 0 59340 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _064_
timestamp 1649977179
transform -1 0 61180 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _065_
timestamp 1649977179
transform 1 0 59984 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _066_
timestamp 1649977179
transform 1 0 59248 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _067_
timestamp 1649977179
transform 1 0 59248 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _068_
timestamp 1649977179
transform 1 0 61732 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _069_
timestamp 1649977179
transform -1 0 61732 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _070_
timestamp 1649977179
transform 1 0 61824 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _071_
timestamp 1649977179
transform 1 0 63020 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _072_
timestamp 1649977179
transform 1 0 62836 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _073_
timestamp 1649977179
transform 1 0 61824 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _074_
timestamp 1649977179
transform 1 0 61732 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _075_
timestamp 1649977179
transform -1 0 65044 0 -1 58752
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _076_
timestamp 1649977179
transform -1 0 64676 0 1 58752
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_2  _077_
timestamp 1649977179
transform 1 0 64400 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _078_
timestamp 1649977179
transform 1 0 64400 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _079_
timestamp 1649977179
transform 1 0 64400 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _080_
timestamp 1649977179
transform 1 0 63296 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _081_
timestamp 1649977179
transform 1 0 65504 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _082_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 65872 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 63388 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _084_
timestamp 1649977179
transform 1 0 65596 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _085_
timestamp 1649977179
transform 1 0 65596 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _086_
timestamp 1649977179
transform 1 0 64400 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _087_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 67160 0 1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 66976 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _089_
timestamp 1649977179
transform 1 0 65504 0 -1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _090_
timestamp 1649977179
transform 1 0 66332 0 -1 60928
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _091_
timestamp 1649977179
transform 1 0 63572 0 -1 60928
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _092_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 64124 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _093_
timestamp 1649977179
transform 1 0 63572 0 1 59840
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1649977179
transform -1 0 64032 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1649977179
transform 1 0 6440 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1649977179
transform 1 0 6900 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1649977179
transform 1 0 7452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1649977179
transform 1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1649977179
transform 1 0 10672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1649977179
transform 1 0 11960 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1649977179
transform 1 0 27784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1649977179
transform 1 0 27232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1649977179
transform 1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1649977179
transform 1 0 27876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1649977179
transform 1 0 27968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1649977179
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1649977179
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1649977179
transform 1 0 32016 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1649977179
transform 1 0 31464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1649977179
transform 1 0 27876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1649977179
transform 1 0 27692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1649977179
transform 1 0 27692 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1649977179
transform 1 0 31924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1649977179
transform 1 0 32476 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1649977179
transform 1 0 32568 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1649977179
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1649977179
transform 1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1649977179
transform 1 0 3220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1649977179
transform 1 0 3864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1649977179
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1649977179
transform 1 0 6716 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1649977179
transform 1 0 7544 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1649977179
transform 1 0 9384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1649977179
transform 1 0 10396 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1649977179
transform 1 0 13432 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1649977179
transform 1 0 12696 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _145_
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1649977179
transform 1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1649977179
transform 1 0 16100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1649977179
transform 1 0 18492 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1649977179
transform 1 0 17848 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1649977179
transform 1 0 19044 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1649977179
transform 1 0 19688 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1649977179
transform 1 0 22264 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1649977179
transform 1 0 22264 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1649977179
transform -1 0 23184 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1649977179
transform 1 0 27324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1649977179
transform 1 0 28704 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1649977179
transform 1 0 29440 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1649977179
transform 1 0 30084 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _165_
timestamp 1649977179
transform 1 0 30820 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1649977179
transform 1 0 32200 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1649977179
transform 1 0 32844 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1649977179
transform 1 0 33580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1649977179
transform 1 0 34960 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1649977179
transform 1 0 35696 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1649977179
transform 1 0 36432 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1649977179
transform 1 0 37812 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1649977179
transform 1 0 38548 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1649977179
transform 1 0 39284 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1649977179
transform 1 0 40020 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1649977179
transform 1 0 40756 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1649977179
transform 1 0 41492 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1649977179
transform 1 0 42228 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1649977179
transform 1 0 43148 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _183_
timestamp 1649977179
transform 1 0 43608 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1649977179
transform 1 0 44344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1649977179
transform 1 0 45080 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1649977179
transform 1 0 45816 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1649977179
transform 1 0 46552 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1649977179
transform 1 0 47288 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1649977179
transform 1 0 48024 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1649977179
transform 1 0 48760 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1649977179
transform -1 0 25484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1649977179
transform -1 0 26312 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1649977179
transform -1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1649977179
transform -1 0 27784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _195_
timestamp 1649977179
transform -1 0 28520 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _196_
timestamp 1649977179
transform -1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _197_
timestamp 1649977179
transform -1 0 29992 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1649977179
transform -1 0 30728 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _199_
timestamp 1649977179
transform -1 0 31464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _200_
timestamp 1649977179
transform -1 0 32476 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _201_
timestamp 1649977179
transform -1 0 32936 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _202_
timestamp 1649977179
transform -1 0 33672 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _203_
timestamp 1649977179
transform -1 0 34408 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _204_
timestamp 1649977179
transform -1 0 35144 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _205_
timestamp 1649977179
transform -1 0 35880 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _206_
timestamp 1649977179
transform -1 0 36524 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _207_
timestamp 1649977179
transform -1 0 37260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _208_
timestamp 1649977179
transform -1 0 37996 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _209_
timestamp 1649977179
transform -1 0 38732 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _210_
timestamp 1649977179
transform -1 0 39376 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _211_
timestamp 1649977179
transform -1 0 40204 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _212_
timestamp 1649977179
transform -1 0 40940 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _213_
timestamp 1649977179
transform -1 0 41676 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _214_
timestamp 1649977179
transform -1 0 42780 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _215_
timestamp 1649977179
transform -1 0 43056 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _216_
timestamp 1649977179
transform -1 0 43792 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _217_
timestamp 1649977179
transform -1 0 44528 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _218_
timestamp 1649977179
transform -1 0 45356 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _219_
timestamp 1649977179
transform -1 0 45908 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _220_
timestamp 1649977179
transform -1 0 46644 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _221_
timestamp 1649977179
transform -1 0 47380 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _222_
timestamp 1649977179
transform -1 0 48024 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1649977179
transform -1 0 74152 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _224_
timestamp 1649977179
transform -1 0 74888 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1649977179
transform -1 0 76176 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _226_
timestamp 1649977179
transform -1 0 76268 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _227_
timestamp 1649977179
transform -1 0 71116 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _228_
timestamp 1649977179
transform -1 0 71484 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _229_
timestamp 1649977179
transform -1 0 72128 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _230_
timestamp 1649977179
transform -1 0 72680 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _231_
timestamp 1649977179
transform -1 0 73416 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _232_
timestamp 1649977179
transform -1 0 70196 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1649977179
transform -1 0 78016 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1649977179
transform 1 0 1380 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 2392 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform -1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform -1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1649977179
transform -1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform -1 0 19872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform -1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform -1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1649977179
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 22724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1649977179
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 24196 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform -1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 5612 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input35
timestamp 1649977179
transform -1 0 78016 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1649977179
transform 1 0 77096 0 -1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 77924 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform 1 0 77740 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 77924 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform 1 0 77740 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 77740 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 77924 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform 1 0 77740 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform 1 0 77924 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 77924 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform 1 0 77740 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1649977179
transform -1 0 78200 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform 1 0 77924 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform 1 0 77740 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform 1 0 77740 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform 1 0 77924 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform 1 0 77740 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 77924 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform 1 0 77924 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform 1 0 77740 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform 1 0 77924 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform 1 0 77740 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1649977179
transform 1 0 77280 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform 1 0 77740 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform 1 0 77924 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1649977179
transform 1 0 77096 0 -1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1649977179
transform 1 0 77280 0 1 51136
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1649977179
transform -1 0 78016 0 -1 52224
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1649977179
transform -1 0 78016 0 -1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1649977179
transform 1 0 77280 0 1 53312
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1649977179
transform -1 0 78016 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1649977179
transform 1 0 77924 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1649977179
transform 1 0 1380 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1649977179
transform 1 0 1380 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1649977179
transform 1 0 1380 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1649977179
transform 1 0 1380 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1649977179
transform 1 0 1380 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1649977179
transform 1 0 1380 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1649977179
transform 1 0 1380 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input81
timestamp 1649977179
transform 1 0 1380 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input82
timestamp 1649977179
transform 1 0 1380 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input83
timestamp 1649977179
transform 1 0 1380 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input84
timestamp 1649977179
transform 1 0 1380 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input85
timestamp 1649977179
transform 1 0 1380 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1649977179
transform 1 0 1380 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input87
timestamp 1649977179
transform 1 0 1380 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1649977179
transform 1 0 1380 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1649977179
transform 1 0 1380 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1649977179
transform 1 0 1380 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1649977179
transform 1 0 1380 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input94
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input95
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input96
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input99
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input100
timestamp 1649977179
transform -1 0 26496 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1649977179
transform 1 0 33028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1649977179
transform 1 0 33764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input103
timestamp 1649977179
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1649977179
transform -1 0 35328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input105
timestamp 1649977179
transform -1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1649977179
transform -1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1649977179
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1649977179
transform 1 0 38916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1649977179
transform 1 0 39652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input111
timestamp 1649977179
transform -1 0 26496 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1649977179
transform 1 0 40388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input113
timestamp 1649977179
transform 1 0 41124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input114
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1649977179
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1649977179
transform 1 0 43884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 1649977179
transform 1 0 44068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1649977179
transform 1 0 45724 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1649977179
transform 1 0 46460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input122
timestamp 1649977179
transform 1 0 27140 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input123
timestamp 1649977179
transform 1 0 48300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input124
timestamp 1649977179
transform 1 0 49036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input125
timestamp 1649977179
transform -1 0 28428 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input126
timestamp 1649977179
transform -1 0 29072 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input127
timestamp 1649977179
transform -1 0 29716 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input128
timestamp 1649977179
transform 1 0 30084 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input129
timestamp 1649977179
transform 1 0 30728 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input130
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 1649977179
transform 1 0 32292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input132
timestamp 1649977179
transform 1 0 74060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input133
timestamp 1649977179
transform 1 0 74796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input134
timestamp 1649977179
transform 1 0 74980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input135
timestamp 1649977179
transform 1 0 75900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input136
timestamp 1649977179
transform 1 0 76636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input137
timestamp 1649977179
transform 1 0 73324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform 1 0 77372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform 1 0 77648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform 1 0 77832 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform 1 0 77648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform 1 0 77832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 77648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 77648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 77832 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 77648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 77832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 77832 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1649977179
transform 1 0 77648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1649977179
transform 1 0 77832 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1649977179
transform 1 0 77832 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1649977179
transform 1 0 77648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1649977179
transform 1 0 77648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1649977179
transform 1 0 77832 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1649977179
transform 1 0 77648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1649977179
transform 1 0 77832 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1649977179
transform 1 0 77832 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1649977179
transform 1 0 77648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1649977179
transform 1 0 77832 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1649977179
transform 1 0 77648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1649977179
transform 1 0 77832 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1649977179
transform 1 0 77648 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1649977179
transform 1 0 77832 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1649977179
transform 1 0 77648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1649977179
transform 1 0 77832 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1649977179
transform 1 0 77648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1649977179
transform 1 0 77648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1649977179
transform 1 0 77832 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1649977179
transform 1 0 77648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1649977179
transform 1 0 77832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1649977179
transform -1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1649977179
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1649977179
transform -1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1649977179
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1649977179
transform -1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1649977179
transform -1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1649977179
transform -1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1649977179
transform -1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1649977179
transform -1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1649977179
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1649977179
transform -1 0 1748 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1649977179
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1649977179
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1649977179
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1649977179
transform -1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1649977179
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1649977179
transform -1 0 1748 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1649977179
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1649977179
transform 1 0 77832 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1649977179
transform -1 0 1748 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1649977179
transform -1 0 49588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1649977179
transform -1 0 57132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1649977179
transform 1 0 57868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1649977179
transform 1 0 58604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1649977179
transform 1 0 59340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1649977179
transform -1 0 59892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1649977179
transform -1 0 60812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1649977179
transform -1 0 61548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1649977179
transform 1 0 61916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1649977179
transform 1 0 63020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1649977179
transform 1 0 63756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1649977179
transform -1 0 50508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1649977179
transform 1 0 64492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1649977179
transform 1 0 64676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1649977179
transform 1 0 66332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1649977179
transform 1 0 67068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1649977179
transform 1 0 68908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1649977179
transform 1 0 69644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1649977179
transform 1 0 69828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1649977179
transform 1 0 70748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1649977179
transform -1 0 51244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1649977179
transform 1 0 71484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1649977179
transform 1 0 72220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1649977179
transform -1 0 51980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1649977179
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1649977179
transform -1 0 53820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1649977179
transform 1 0 54188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1649977179
transform 1 0 54372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1649977179
transform 1 0 55292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1649977179
transform -1 0 56396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1649977179
transform 1 0 77648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1649977179
transform 1 0 77832 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1649977179
transform 1 0 77648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1649977179
transform 1 0 77832 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1649977179
transform 1 0 77648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1649977179
transform 1 0 77648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1649977179
transform 1 0 77832 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1649977179
transform 1 0 77648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1649977179
transform 1 0 77832 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1649977179
transform 1 0 77832 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1649977179
transform 1 0 77648 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1649977179
transform 1 0 77832 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1649977179
transform 1 0 77832 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1649977179
transform 1 0 77648 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1649977179
transform 1 0 77648 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1649977179
transform 1 0 77832 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1649977179
transform 1 0 77648 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1649977179
transform 1 0 77832 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1649977179
transform 1 0 77832 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1649977179
transform 1 0 77648 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1649977179
transform 1 0 77832 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1649977179
transform 1 0 77648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1649977179
transform 1 0 77832 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1649977179
transform 1 0 77648 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1649977179
transform 1 0 77832 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1649977179
transform 1 0 77648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1649977179
transform 1 0 77832 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1649977179
transform 1 0 77648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1649977179
transform 1 0 77648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1649977179
transform 1 0 77832 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1649977179
transform 1 0 77648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1649977179
transform 1 0 77832 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1649977179
transform -1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1649977179
transform -1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1649977179
transform -1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1649977179
transform -1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1649977179
transform -1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1649977179
transform -1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1649977179
transform -1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1649977179
transform -1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1649977179
transform -1 0 1748 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1649977179
transform -1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1649977179
transform -1 0 1748 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output280
timestamp 1649977179
transform -1 0 1748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1649977179
transform -1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output282
timestamp 1649977179
transform -1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output283
timestamp 1649977179
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output284
timestamp 1649977179
transform -1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output285
timestamp 1649977179
transform -1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output286
timestamp 1649977179
transform -1 0 1748 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output287
timestamp 1649977179
transform -1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output288
timestamp 1649977179
transform -1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output289
timestamp 1649977179
transform -1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output290
timestamp 1649977179
transform -1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output291
timestamp 1649977179
transform -1 0 1748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output292
timestamp 1649977179
transform -1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output293
timestamp 1649977179
transform -1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output294
timestamp 1649977179
transform -1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output295
timestamp 1649977179
transform -1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output296
timestamp 1649977179
transform -1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output297
timestamp 1649977179
transform -1 0 1748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output298
timestamp 1649977179
transform -1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output299
timestamp 1649977179
transform -1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output300
timestamp 1649977179
transform -1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output301
timestamp 1649977179
transform 1 0 77832 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output302
timestamp 1649977179
transform 1 0 77832 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output303
timestamp 1649977179
transform 1 0 77648 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output304
timestamp 1649977179
transform 1 0 77832 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output305
timestamp 1649977179
transform -1 0 1748 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output306
timestamp 1649977179
transform -1 0 1748 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output307
timestamp 1649977179
transform -1 0 1748 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output308
timestamp 1649977179
transform -1 0 1748 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output309
timestamp 1649977179
transform 1 0 77648 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output310
timestamp 1649977179
transform -1 0 1748 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output311
timestamp 1649977179
transform 1 0 77648 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output312
timestamp 1649977179
transform -1 0 1748 0 -1 70720
box -38 -48 406 592
<< labels >>
flabel metal2 s 77114 0 77170 800 0 FreeSans 224 90 0 0 io_wbs_ack
port 0 nsew signal tristate
flabel metal3 s 79200 74264 80000 74384 0 FreeSans 480 0 0 0 io_wbs_ack_0
port 1 nsew signal input
flabel metal3 s 0 74264 800 74384 0 FreeSans 480 0 0 0 io_wbs_ack_1
port 2 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 io_wbs_adr[0]
port 3 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 io_wbs_adr[10]
port 4 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 io_wbs_adr[11]
port 5 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 io_wbs_adr[12]
port 6 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 io_wbs_adr[13]
port 7 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 io_wbs_adr[14]
port 8 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 io_wbs_adr[15]
port 9 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 io_wbs_adr[16]
port 10 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 io_wbs_adr[17]
port 11 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 io_wbs_adr[18]
port 12 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 io_wbs_adr[19]
port 13 nsew signal input
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 io_wbs_adr[1]
port 14 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 io_wbs_adr[20]
port 15 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 io_wbs_adr[21]
port 16 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 io_wbs_adr[22]
port 17 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 io_wbs_adr[23]
port 18 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 io_wbs_adr[24]
port 19 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 io_wbs_adr[25]
port 20 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 io_wbs_adr[26]
port 21 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 io_wbs_adr[27]
port 22 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 io_wbs_adr[28]
port 23 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 io_wbs_adr[29]
port 24 nsew signal input
flabel metal2 s 3514 0 3570 800 0 FreeSans 224 90 0 0 io_wbs_adr[2]
port 25 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 io_wbs_adr[30]
port 26 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 io_wbs_adr[31]
port 27 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 io_wbs_adr[3]
port 28 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 io_wbs_adr[4]
port 29 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 io_wbs_adr[5]
port 30 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 io_wbs_adr[6]
port 31 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 io_wbs_adr[7]
port 32 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 io_wbs_adr[8]
port 33 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 io_wbs_adr[9]
port 34 nsew signal input
flabel metal3 s 79200 4904 80000 5024 0 FreeSans 480 0 0 0 io_wbs_adr_0[0]
port 35 nsew signal tristate
flabel metal3 s 79200 11704 80000 11824 0 FreeSans 480 0 0 0 io_wbs_adr_0[10]
port 36 nsew signal tristate
flabel metal3 s 79200 12384 80000 12504 0 FreeSans 480 0 0 0 io_wbs_adr_0[11]
port 37 nsew signal tristate
flabel metal3 s 79200 13064 80000 13184 0 FreeSans 480 0 0 0 io_wbs_adr_0[12]
port 38 nsew signal tristate
flabel metal3 s 79200 13744 80000 13864 0 FreeSans 480 0 0 0 io_wbs_adr_0[13]
port 39 nsew signal tristate
flabel metal3 s 79200 14424 80000 14544 0 FreeSans 480 0 0 0 io_wbs_adr_0[14]
port 40 nsew signal tristate
flabel metal3 s 79200 15104 80000 15224 0 FreeSans 480 0 0 0 io_wbs_adr_0[15]
port 41 nsew signal tristate
flabel metal3 s 79200 15784 80000 15904 0 FreeSans 480 0 0 0 io_wbs_adr_0[16]
port 42 nsew signal tristate
flabel metal3 s 79200 16464 80000 16584 0 FreeSans 480 0 0 0 io_wbs_adr_0[17]
port 43 nsew signal tristate
flabel metal3 s 79200 17144 80000 17264 0 FreeSans 480 0 0 0 io_wbs_adr_0[18]
port 44 nsew signal tristate
flabel metal3 s 79200 17824 80000 17944 0 FreeSans 480 0 0 0 io_wbs_adr_0[19]
port 45 nsew signal tristate
flabel metal3 s 79200 5584 80000 5704 0 FreeSans 480 0 0 0 io_wbs_adr_0[1]
port 46 nsew signal tristate
flabel metal3 s 79200 18504 80000 18624 0 FreeSans 480 0 0 0 io_wbs_adr_0[20]
port 47 nsew signal tristate
flabel metal3 s 79200 19184 80000 19304 0 FreeSans 480 0 0 0 io_wbs_adr_0[21]
port 48 nsew signal tristate
flabel metal3 s 79200 19864 80000 19984 0 FreeSans 480 0 0 0 io_wbs_adr_0[22]
port 49 nsew signal tristate
flabel metal3 s 79200 20544 80000 20664 0 FreeSans 480 0 0 0 io_wbs_adr_0[23]
port 50 nsew signal tristate
flabel metal3 s 79200 21224 80000 21344 0 FreeSans 480 0 0 0 io_wbs_adr_0[24]
port 51 nsew signal tristate
flabel metal3 s 79200 21904 80000 22024 0 FreeSans 480 0 0 0 io_wbs_adr_0[25]
port 52 nsew signal tristate
flabel metal3 s 79200 22584 80000 22704 0 FreeSans 480 0 0 0 io_wbs_adr_0[26]
port 53 nsew signal tristate
flabel metal3 s 79200 23264 80000 23384 0 FreeSans 480 0 0 0 io_wbs_adr_0[27]
port 54 nsew signal tristate
flabel metal3 s 79200 23944 80000 24064 0 FreeSans 480 0 0 0 io_wbs_adr_0[28]
port 55 nsew signal tristate
flabel metal3 s 79200 24624 80000 24744 0 FreeSans 480 0 0 0 io_wbs_adr_0[29]
port 56 nsew signal tristate
flabel metal3 s 79200 6264 80000 6384 0 FreeSans 480 0 0 0 io_wbs_adr_0[2]
port 57 nsew signal tristate
flabel metal3 s 79200 25304 80000 25424 0 FreeSans 480 0 0 0 io_wbs_adr_0[30]
port 58 nsew signal tristate
flabel metal3 s 79200 25984 80000 26104 0 FreeSans 480 0 0 0 io_wbs_adr_0[31]
port 59 nsew signal tristate
flabel metal3 s 79200 6944 80000 7064 0 FreeSans 480 0 0 0 io_wbs_adr_0[3]
port 60 nsew signal tristate
flabel metal3 s 79200 7624 80000 7744 0 FreeSans 480 0 0 0 io_wbs_adr_0[4]
port 61 nsew signal tristate
flabel metal3 s 79200 8304 80000 8424 0 FreeSans 480 0 0 0 io_wbs_adr_0[5]
port 62 nsew signal tristate
flabel metal3 s 79200 8984 80000 9104 0 FreeSans 480 0 0 0 io_wbs_adr_0[6]
port 63 nsew signal tristate
flabel metal3 s 79200 9664 80000 9784 0 FreeSans 480 0 0 0 io_wbs_adr_0[7]
port 64 nsew signal tristate
flabel metal3 s 79200 10344 80000 10464 0 FreeSans 480 0 0 0 io_wbs_adr_0[8]
port 65 nsew signal tristate
flabel metal3 s 79200 11024 80000 11144 0 FreeSans 480 0 0 0 io_wbs_adr_0[9]
port 66 nsew signal tristate
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 io_wbs_adr_1[0]
port 67 nsew signal tristate
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 io_wbs_adr_1[10]
port 68 nsew signal tristate
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 io_wbs_adr_1[11]
port 69 nsew signal tristate
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 io_wbs_adr_1[12]
port 70 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 io_wbs_adr_1[13]
port 71 nsew signal tristate
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 io_wbs_adr_1[14]
port 72 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 io_wbs_adr_1[15]
port 73 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 io_wbs_adr_1[16]
port 74 nsew signal tristate
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 io_wbs_adr_1[17]
port 75 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 io_wbs_adr_1[18]
port 76 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 io_wbs_adr_1[19]
port 77 nsew signal tristate
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 io_wbs_adr_1[1]
port 78 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 io_wbs_adr_1[20]
port 79 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 io_wbs_adr_1[21]
port 80 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 io_wbs_adr_1[22]
port 81 nsew signal tristate
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 io_wbs_adr_1[23]
port 82 nsew signal tristate
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 io_wbs_adr_1[24]
port 83 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 io_wbs_adr_1[25]
port 84 nsew signal tristate
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 io_wbs_adr_1[26]
port 85 nsew signal tristate
flabel metal3 s 0 23264 800 23384 0 FreeSans 480 0 0 0 io_wbs_adr_1[27]
port 86 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 io_wbs_adr_1[28]
port 87 nsew signal tristate
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 io_wbs_adr_1[29]
port 88 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 io_wbs_adr_1[2]
port 89 nsew signal tristate
flabel metal3 s 0 25304 800 25424 0 FreeSans 480 0 0 0 io_wbs_adr_1[30]
port 90 nsew signal tristate
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 io_wbs_adr_1[31]
port 91 nsew signal tristate
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 io_wbs_adr_1[3]
port 92 nsew signal tristate
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 io_wbs_adr_1[4]
port 93 nsew signal tristate
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 io_wbs_adr_1[5]
port 94 nsew signal tristate
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 io_wbs_adr_1[6]
port 95 nsew signal tristate
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_wbs_adr_1[7]
port 96 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 io_wbs_adr_1[8]
port 97 nsew signal tristate
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 io_wbs_adr_1[9]
port 98 nsew signal tristate
flabel metal2 s 77850 0 77906 800 0 FreeSans 224 90 0 0 io_wbs_cyc
port 99 nsew signal input
flabel metal3 s 79200 74944 80000 75064 0 FreeSans 480 0 0 0 io_wbs_cyc_0
port 100 nsew signal tristate
flabel metal3 s 0 74944 800 75064 0 FreeSans 480 0 0 0 io_wbs_cyc_1
port 101 nsew signal tristate
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 io_wbs_datrd[0]
port 102 nsew signal tristate
flabel metal2 s 56506 0 56562 800 0 FreeSans 224 90 0 0 io_wbs_datrd[10]
port 103 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 io_wbs_datrd[11]
port 104 nsew signal tristate
flabel metal2 s 57978 0 58034 800 0 FreeSans 224 90 0 0 io_wbs_datrd[12]
port 105 nsew signal tristate
flabel metal2 s 58714 0 58770 800 0 FreeSans 224 90 0 0 io_wbs_datrd[13]
port 106 nsew signal tristate
flabel metal2 s 59450 0 59506 800 0 FreeSans 224 90 0 0 io_wbs_datrd[14]
port 107 nsew signal tristate
flabel metal2 s 60186 0 60242 800 0 FreeSans 224 90 0 0 io_wbs_datrd[15]
port 108 nsew signal tristate
flabel metal2 s 60922 0 60978 800 0 FreeSans 224 90 0 0 io_wbs_datrd[16]
port 109 nsew signal tristate
flabel metal2 s 61658 0 61714 800 0 FreeSans 224 90 0 0 io_wbs_datrd[17]
port 110 nsew signal tristate
flabel metal2 s 62394 0 62450 800 0 FreeSans 224 90 0 0 io_wbs_datrd[18]
port 111 nsew signal tristate
flabel metal2 s 63130 0 63186 800 0 FreeSans 224 90 0 0 io_wbs_datrd[19]
port 112 nsew signal tristate
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 io_wbs_datrd[1]
port 113 nsew signal tristate
flabel metal2 s 63866 0 63922 800 0 FreeSans 224 90 0 0 io_wbs_datrd[20]
port 114 nsew signal tristate
flabel metal2 s 64602 0 64658 800 0 FreeSans 224 90 0 0 io_wbs_datrd[21]
port 115 nsew signal tristate
flabel metal2 s 65338 0 65394 800 0 FreeSans 224 90 0 0 io_wbs_datrd[22]
port 116 nsew signal tristate
flabel metal2 s 66074 0 66130 800 0 FreeSans 224 90 0 0 io_wbs_datrd[23]
port 117 nsew signal tristate
flabel metal2 s 66810 0 66866 800 0 FreeSans 224 90 0 0 io_wbs_datrd[24]
port 118 nsew signal tristate
flabel metal2 s 67546 0 67602 800 0 FreeSans 224 90 0 0 io_wbs_datrd[25]
port 119 nsew signal tristate
flabel metal2 s 68282 0 68338 800 0 FreeSans 224 90 0 0 io_wbs_datrd[26]
port 120 nsew signal tristate
flabel metal2 s 69018 0 69074 800 0 FreeSans 224 90 0 0 io_wbs_datrd[27]
port 121 nsew signal tristate
flabel metal2 s 69754 0 69810 800 0 FreeSans 224 90 0 0 io_wbs_datrd[28]
port 122 nsew signal tristate
flabel metal2 s 70490 0 70546 800 0 FreeSans 224 90 0 0 io_wbs_datrd[29]
port 123 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 io_wbs_datrd[2]
port 124 nsew signal tristate
flabel metal2 s 71226 0 71282 800 0 FreeSans 224 90 0 0 io_wbs_datrd[30]
port 125 nsew signal tristate
flabel metal2 s 71962 0 72018 800 0 FreeSans 224 90 0 0 io_wbs_datrd[31]
port 126 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 io_wbs_datrd[3]
port 127 nsew signal tristate
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 io_wbs_datrd[4]
port 128 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 io_wbs_datrd[5]
port 129 nsew signal tristate
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 io_wbs_datrd[6]
port 130 nsew signal tristate
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 io_wbs_datrd[7]
port 131 nsew signal tristate
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 io_wbs_datrd[8]
port 132 nsew signal tristate
flabel metal2 s 55770 0 55826 800 0 FreeSans 224 90 0 0 io_wbs_datrd[9]
port 133 nsew signal tristate
flabel metal3 s 79200 48424 80000 48544 0 FreeSans 480 0 0 0 io_wbs_datrd_0[0]
port 134 nsew signal input
flabel metal3 s 79200 55224 80000 55344 0 FreeSans 480 0 0 0 io_wbs_datrd_0[10]
port 135 nsew signal input
flabel metal3 s 79200 55904 80000 56024 0 FreeSans 480 0 0 0 io_wbs_datrd_0[11]
port 136 nsew signal input
flabel metal3 s 79200 56584 80000 56704 0 FreeSans 480 0 0 0 io_wbs_datrd_0[12]
port 137 nsew signal input
flabel metal3 s 79200 57264 80000 57384 0 FreeSans 480 0 0 0 io_wbs_datrd_0[13]
port 138 nsew signal input
flabel metal3 s 79200 57944 80000 58064 0 FreeSans 480 0 0 0 io_wbs_datrd_0[14]
port 139 nsew signal input
flabel metal3 s 79200 58624 80000 58744 0 FreeSans 480 0 0 0 io_wbs_datrd_0[15]
port 140 nsew signal input
flabel metal3 s 79200 59304 80000 59424 0 FreeSans 480 0 0 0 io_wbs_datrd_0[16]
port 141 nsew signal input
flabel metal3 s 79200 59984 80000 60104 0 FreeSans 480 0 0 0 io_wbs_datrd_0[17]
port 142 nsew signal input
flabel metal3 s 79200 60664 80000 60784 0 FreeSans 480 0 0 0 io_wbs_datrd_0[18]
port 143 nsew signal input
flabel metal3 s 79200 61344 80000 61464 0 FreeSans 480 0 0 0 io_wbs_datrd_0[19]
port 144 nsew signal input
flabel metal3 s 79200 49104 80000 49224 0 FreeSans 480 0 0 0 io_wbs_datrd_0[1]
port 145 nsew signal input
flabel metal3 s 79200 62024 80000 62144 0 FreeSans 480 0 0 0 io_wbs_datrd_0[20]
port 146 nsew signal input
flabel metal3 s 79200 62704 80000 62824 0 FreeSans 480 0 0 0 io_wbs_datrd_0[21]
port 147 nsew signal input
flabel metal3 s 79200 63384 80000 63504 0 FreeSans 480 0 0 0 io_wbs_datrd_0[22]
port 148 nsew signal input
flabel metal3 s 79200 64064 80000 64184 0 FreeSans 480 0 0 0 io_wbs_datrd_0[23]
port 149 nsew signal input
flabel metal3 s 79200 64744 80000 64864 0 FreeSans 480 0 0 0 io_wbs_datrd_0[24]
port 150 nsew signal input
flabel metal3 s 79200 65424 80000 65544 0 FreeSans 480 0 0 0 io_wbs_datrd_0[25]
port 151 nsew signal input
flabel metal3 s 79200 66104 80000 66224 0 FreeSans 480 0 0 0 io_wbs_datrd_0[26]
port 152 nsew signal input
flabel metal3 s 79200 66784 80000 66904 0 FreeSans 480 0 0 0 io_wbs_datrd_0[27]
port 153 nsew signal input
flabel metal3 s 79200 67464 80000 67584 0 FreeSans 480 0 0 0 io_wbs_datrd_0[28]
port 154 nsew signal input
flabel metal3 s 79200 68144 80000 68264 0 FreeSans 480 0 0 0 io_wbs_datrd_0[29]
port 155 nsew signal input
flabel metal3 s 79200 49784 80000 49904 0 FreeSans 480 0 0 0 io_wbs_datrd_0[2]
port 156 nsew signal input
flabel metal3 s 79200 68824 80000 68944 0 FreeSans 480 0 0 0 io_wbs_datrd_0[30]
port 157 nsew signal input
flabel metal3 s 79200 69504 80000 69624 0 FreeSans 480 0 0 0 io_wbs_datrd_0[31]
port 158 nsew signal input
flabel metal3 s 79200 50464 80000 50584 0 FreeSans 480 0 0 0 io_wbs_datrd_0[3]
port 159 nsew signal input
flabel metal3 s 79200 51144 80000 51264 0 FreeSans 480 0 0 0 io_wbs_datrd_0[4]
port 160 nsew signal input
flabel metal3 s 79200 51824 80000 51944 0 FreeSans 480 0 0 0 io_wbs_datrd_0[5]
port 161 nsew signal input
flabel metal3 s 79200 52504 80000 52624 0 FreeSans 480 0 0 0 io_wbs_datrd_0[6]
port 162 nsew signal input
flabel metal3 s 79200 53184 80000 53304 0 FreeSans 480 0 0 0 io_wbs_datrd_0[7]
port 163 nsew signal input
flabel metal3 s 79200 53864 80000 53984 0 FreeSans 480 0 0 0 io_wbs_datrd_0[8]
port 164 nsew signal input
flabel metal3 s 79200 54544 80000 54664 0 FreeSans 480 0 0 0 io_wbs_datrd_0[9]
port 165 nsew signal input
flabel metal3 s 0 48424 800 48544 0 FreeSans 480 0 0 0 io_wbs_datrd_1[0]
port 166 nsew signal input
flabel metal3 s 0 55224 800 55344 0 FreeSans 480 0 0 0 io_wbs_datrd_1[10]
port 167 nsew signal input
flabel metal3 s 0 55904 800 56024 0 FreeSans 480 0 0 0 io_wbs_datrd_1[11]
port 168 nsew signal input
flabel metal3 s 0 56584 800 56704 0 FreeSans 480 0 0 0 io_wbs_datrd_1[12]
port 169 nsew signal input
flabel metal3 s 0 57264 800 57384 0 FreeSans 480 0 0 0 io_wbs_datrd_1[13]
port 170 nsew signal input
flabel metal3 s 0 57944 800 58064 0 FreeSans 480 0 0 0 io_wbs_datrd_1[14]
port 171 nsew signal input
flabel metal3 s 0 58624 800 58744 0 FreeSans 480 0 0 0 io_wbs_datrd_1[15]
port 172 nsew signal input
flabel metal3 s 0 59304 800 59424 0 FreeSans 480 0 0 0 io_wbs_datrd_1[16]
port 173 nsew signal input
flabel metal3 s 0 59984 800 60104 0 FreeSans 480 0 0 0 io_wbs_datrd_1[17]
port 174 nsew signal input
flabel metal3 s 0 60664 800 60784 0 FreeSans 480 0 0 0 io_wbs_datrd_1[18]
port 175 nsew signal input
flabel metal3 s 0 61344 800 61464 0 FreeSans 480 0 0 0 io_wbs_datrd_1[19]
port 176 nsew signal input
flabel metal3 s 0 49104 800 49224 0 FreeSans 480 0 0 0 io_wbs_datrd_1[1]
port 177 nsew signal input
flabel metal3 s 0 62024 800 62144 0 FreeSans 480 0 0 0 io_wbs_datrd_1[20]
port 178 nsew signal input
flabel metal3 s 0 62704 800 62824 0 FreeSans 480 0 0 0 io_wbs_datrd_1[21]
port 179 nsew signal input
flabel metal3 s 0 63384 800 63504 0 FreeSans 480 0 0 0 io_wbs_datrd_1[22]
port 180 nsew signal input
flabel metal3 s 0 64064 800 64184 0 FreeSans 480 0 0 0 io_wbs_datrd_1[23]
port 181 nsew signal input
flabel metal3 s 0 64744 800 64864 0 FreeSans 480 0 0 0 io_wbs_datrd_1[24]
port 182 nsew signal input
flabel metal3 s 0 65424 800 65544 0 FreeSans 480 0 0 0 io_wbs_datrd_1[25]
port 183 nsew signal input
flabel metal3 s 0 66104 800 66224 0 FreeSans 480 0 0 0 io_wbs_datrd_1[26]
port 184 nsew signal input
flabel metal3 s 0 66784 800 66904 0 FreeSans 480 0 0 0 io_wbs_datrd_1[27]
port 185 nsew signal input
flabel metal3 s 0 67464 800 67584 0 FreeSans 480 0 0 0 io_wbs_datrd_1[28]
port 186 nsew signal input
flabel metal3 s 0 68144 800 68264 0 FreeSans 480 0 0 0 io_wbs_datrd_1[29]
port 187 nsew signal input
flabel metal3 s 0 49784 800 49904 0 FreeSans 480 0 0 0 io_wbs_datrd_1[2]
port 188 nsew signal input
flabel metal3 s 0 68824 800 68944 0 FreeSans 480 0 0 0 io_wbs_datrd_1[30]
port 189 nsew signal input
flabel metal3 s 0 69504 800 69624 0 FreeSans 480 0 0 0 io_wbs_datrd_1[31]
port 190 nsew signal input
flabel metal3 s 0 50464 800 50584 0 FreeSans 480 0 0 0 io_wbs_datrd_1[3]
port 191 nsew signal input
flabel metal3 s 0 51144 800 51264 0 FreeSans 480 0 0 0 io_wbs_datrd_1[4]
port 192 nsew signal input
flabel metal3 s 0 51824 800 51944 0 FreeSans 480 0 0 0 io_wbs_datrd_1[5]
port 193 nsew signal input
flabel metal3 s 0 52504 800 52624 0 FreeSans 480 0 0 0 io_wbs_datrd_1[6]
port 194 nsew signal input
flabel metal3 s 0 53184 800 53304 0 FreeSans 480 0 0 0 io_wbs_datrd_1[7]
port 195 nsew signal input
flabel metal3 s 0 53864 800 53984 0 FreeSans 480 0 0 0 io_wbs_datrd_1[8]
port 196 nsew signal input
flabel metal3 s 0 54544 800 54664 0 FreeSans 480 0 0 0 io_wbs_datrd_1[9]
port 197 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 io_wbs_datwr[0]
port 198 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 io_wbs_datwr[10]
port 199 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 io_wbs_datwr[11]
port 200 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 io_wbs_datwr[12]
port 201 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 io_wbs_datwr[13]
port 202 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 io_wbs_datwr[14]
port 203 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 io_wbs_datwr[15]
port 204 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 io_wbs_datwr[16]
port 205 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 io_wbs_datwr[17]
port 206 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 io_wbs_datwr[18]
port 207 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 io_wbs_datwr[19]
port 208 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 io_wbs_datwr[1]
port 209 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 io_wbs_datwr[20]
port 210 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 io_wbs_datwr[21]
port 211 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 io_wbs_datwr[22]
port 212 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 io_wbs_datwr[23]
port 213 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 io_wbs_datwr[24]
port 214 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 io_wbs_datwr[25]
port 215 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 io_wbs_datwr[26]
port 216 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 io_wbs_datwr[27]
port 217 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 io_wbs_datwr[28]
port 218 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 io_wbs_datwr[29]
port 219 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 io_wbs_datwr[2]
port 220 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 io_wbs_datwr[30]
port 221 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 io_wbs_datwr[31]
port 222 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 io_wbs_datwr[3]
port 223 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 io_wbs_datwr[4]
port 224 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 io_wbs_datwr[5]
port 225 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 io_wbs_datwr[6]
port 226 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 io_wbs_datwr[7]
port 227 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 io_wbs_datwr[8]
port 228 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 io_wbs_datwr[9]
port 229 nsew signal input
flabel metal3 s 79200 26664 80000 26784 0 FreeSans 480 0 0 0 io_wbs_datwr_0[0]
port 230 nsew signal tristate
flabel metal3 s 79200 33464 80000 33584 0 FreeSans 480 0 0 0 io_wbs_datwr_0[10]
port 231 nsew signal tristate
flabel metal3 s 79200 34144 80000 34264 0 FreeSans 480 0 0 0 io_wbs_datwr_0[11]
port 232 nsew signal tristate
flabel metal3 s 79200 34824 80000 34944 0 FreeSans 480 0 0 0 io_wbs_datwr_0[12]
port 233 nsew signal tristate
flabel metal3 s 79200 35504 80000 35624 0 FreeSans 480 0 0 0 io_wbs_datwr_0[13]
port 234 nsew signal tristate
flabel metal3 s 79200 36184 80000 36304 0 FreeSans 480 0 0 0 io_wbs_datwr_0[14]
port 235 nsew signal tristate
flabel metal3 s 79200 36864 80000 36984 0 FreeSans 480 0 0 0 io_wbs_datwr_0[15]
port 236 nsew signal tristate
flabel metal3 s 79200 37544 80000 37664 0 FreeSans 480 0 0 0 io_wbs_datwr_0[16]
port 237 nsew signal tristate
flabel metal3 s 79200 38224 80000 38344 0 FreeSans 480 0 0 0 io_wbs_datwr_0[17]
port 238 nsew signal tristate
flabel metal3 s 79200 38904 80000 39024 0 FreeSans 480 0 0 0 io_wbs_datwr_0[18]
port 239 nsew signal tristate
flabel metal3 s 79200 39584 80000 39704 0 FreeSans 480 0 0 0 io_wbs_datwr_0[19]
port 240 nsew signal tristate
flabel metal3 s 79200 27344 80000 27464 0 FreeSans 480 0 0 0 io_wbs_datwr_0[1]
port 241 nsew signal tristate
flabel metal3 s 79200 40264 80000 40384 0 FreeSans 480 0 0 0 io_wbs_datwr_0[20]
port 242 nsew signal tristate
flabel metal3 s 79200 40944 80000 41064 0 FreeSans 480 0 0 0 io_wbs_datwr_0[21]
port 243 nsew signal tristate
flabel metal3 s 79200 41624 80000 41744 0 FreeSans 480 0 0 0 io_wbs_datwr_0[22]
port 244 nsew signal tristate
flabel metal3 s 79200 42304 80000 42424 0 FreeSans 480 0 0 0 io_wbs_datwr_0[23]
port 245 nsew signal tristate
flabel metal3 s 79200 42984 80000 43104 0 FreeSans 480 0 0 0 io_wbs_datwr_0[24]
port 246 nsew signal tristate
flabel metal3 s 79200 43664 80000 43784 0 FreeSans 480 0 0 0 io_wbs_datwr_0[25]
port 247 nsew signal tristate
flabel metal3 s 79200 44344 80000 44464 0 FreeSans 480 0 0 0 io_wbs_datwr_0[26]
port 248 nsew signal tristate
flabel metal3 s 79200 45024 80000 45144 0 FreeSans 480 0 0 0 io_wbs_datwr_0[27]
port 249 nsew signal tristate
flabel metal3 s 79200 45704 80000 45824 0 FreeSans 480 0 0 0 io_wbs_datwr_0[28]
port 250 nsew signal tristate
flabel metal3 s 79200 46384 80000 46504 0 FreeSans 480 0 0 0 io_wbs_datwr_0[29]
port 251 nsew signal tristate
flabel metal3 s 79200 28024 80000 28144 0 FreeSans 480 0 0 0 io_wbs_datwr_0[2]
port 252 nsew signal tristate
flabel metal3 s 79200 47064 80000 47184 0 FreeSans 480 0 0 0 io_wbs_datwr_0[30]
port 253 nsew signal tristate
flabel metal3 s 79200 47744 80000 47864 0 FreeSans 480 0 0 0 io_wbs_datwr_0[31]
port 254 nsew signal tristate
flabel metal3 s 79200 28704 80000 28824 0 FreeSans 480 0 0 0 io_wbs_datwr_0[3]
port 255 nsew signal tristate
flabel metal3 s 79200 29384 80000 29504 0 FreeSans 480 0 0 0 io_wbs_datwr_0[4]
port 256 nsew signal tristate
flabel metal3 s 79200 30064 80000 30184 0 FreeSans 480 0 0 0 io_wbs_datwr_0[5]
port 257 nsew signal tristate
flabel metal3 s 79200 30744 80000 30864 0 FreeSans 480 0 0 0 io_wbs_datwr_0[6]
port 258 nsew signal tristate
flabel metal3 s 79200 31424 80000 31544 0 FreeSans 480 0 0 0 io_wbs_datwr_0[7]
port 259 nsew signal tristate
flabel metal3 s 79200 32104 80000 32224 0 FreeSans 480 0 0 0 io_wbs_datwr_0[8]
port 260 nsew signal tristate
flabel metal3 s 79200 32784 80000 32904 0 FreeSans 480 0 0 0 io_wbs_datwr_0[9]
port 261 nsew signal tristate
flabel metal3 s 0 26664 800 26784 0 FreeSans 480 0 0 0 io_wbs_datwr_1[0]
port 262 nsew signal tristate
flabel metal3 s 0 33464 800 33584 0 FreeSans 480 0 0 0 io_wbs_datwr_1[10]
port 263 nsew signal tristate
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 io_wbs_datwr_1[11]
port 264 nsew signal tristate
flabel metal3 s 0 34824 800 34944 0 FreeSans 480 0 0 0 io_wbs_datwr_1[12]
port 265 nsew signal tristate
flabel metal3 s 0 35504 800 35624 0 FreeSans 480 0 0 0 io_wbs_datwr_1[13]
port 266 nsew signal tristate
flabel metal3 s 0 36184 800 36304 0 FreeSans 480 0 0 0 io_wbs_datwr_1[14]
port 267 nsew signal tristate
flabel metal3 s 0 36864 800 36984 0 FreeSans 480 0 0 0 io_wbs_datwr_1[15]
port 268 nsew signal tristate
flabel metal3 s 0 37544 800 37664 0 FreeSans 480 0 0 0 io_wbs_datwr_1[16]
port 269 nsew signal tristate
flabel metal3 s 0 38224 800 38344 0 FreeSans 480 0 0 0 io_wbs_datwr_1[17]
port 270 nsew signal tristate
flabel metal3 s 0 38904 800 39024 0 FreeSans 480 0 0 0 io_wbs_datwr_1[18]
port 271 nsew signal tristate
flabel metal3 s 0 39584 800 39704 0 FreeSans 480 0 0 0 io_wbs_datwr_1[19]
port 272 nsew signal tristate
flabel metal3 s 0 27344 800 27464 0 FreeSans 480 0 0 0 io_wbs_datwr_1[1]
port 273 nsew signal tristate
flabel metal3 s 0 40264 800 40384 0 FreeSans 480 0 0 0 io_wbs_datwr_1[20]
port 274 nsew signal tristate
flabel metal3 s 0 40944 800 41064 0 FreeSans 480 0 0 0 io_wbs_datwr_1[21]
port 275 nsew signal tristate
flabel metal3 s 0 41624 800 41744 0 FreeSans 480 0 0 0 io_wbs_datwr_1[22]
port 276 nsew signal tristate
flabel metal3 s 0 42304 800 42424 0 FreeSans 480 0 0 0 io_wbs_datwr_1[23]
port 277 nsew signal tristate
flabel metal3 s 0 42984 800 43104 0 FreeSans 480 0 0 0 io_wbs_datwr_1[24]
port 278 nsew signal tristate
flabel metal3 s 0 43664 800 43784 0 FreeSans 480 0 0 0 io_wbs_datwr_1[25]
port 279 nsew signal tristate
flabel metal3 s 0 44344 800 44464 0 FreeSans 480 0 0 0 io_wbs_datwr_1[26]
port 280 nsew signal tristate
flabel metal3 s 0 45024 800 45144 0 FreeSans 480 0 0 0 io_wbs_datwr_1[27]
port 281 nsew signal tristate
flabel metal3 s 0 45704 800 45824 0 FreeSans 480 0 0 0 io_wbs_datwr_1[28]
port 282 nsew signal tristate
flabel metal3 s 0 46384 800 46504 0 FreeSans 480 0 0 0 io_wbs_datwr_1[29]
port 283 nsew signal tristate
flabel metal3 s 0 28024 800 28144 0 FreeSans 480 0 0 0 io_wbs_datwr_1[2]
port 284 nsew signal tristate
flabel metal3 s 0 47064 800 47184 0 FreeSans 480 0 0 0 io_wbs_datwr_1[30]
port 285 nsew signal tristate
flabel metal3 s 0 47744 800 47864 0 FreeSans 480 0 0 0 io_wbs_datwr_1[31]
port 286 nsew signal tristate
flabel metal3 s 0 28704 800 28824 0 FreeSans 480 0 0 0 io_wbs_datwr_1[3]
port 287 nsew signal tristate
flabel metal3 s 0 29384 800 29504 0 FreeSans 480 0 0 0 io_wbs_datwr_1[4]
port 288 nsew signal tristate
flabel metal3 s 0 30064 800 30184 0 FreeSans 480 0 0 0 io_wbs_datwr_1[5]
port 289 nsew signal tristate
flabel metal3 s 0 30744 800 30864 0 FreeSans 480 0 0 0 io_wbs_datwr_1[6]
port 290 nsew signal tristate
flabel metal3 s 0 31424 800 31544 0 FreeSans 480 0 0 0 io_wbs_datwr_1[7]
port 291 nsew signal tristate
flabel metal3 s 0 32104 800 32224 0 FreeSans 480 0 0 0 io_wbs_datwr_1[8]
port 292 nsew signal tristate
flabel metal3 s 0 32784 800 32904 0 FreeSans 480 0 0 0 io_wbs_datwr_1[9]
port 293 nsew signal tristate
flabel metal2 s 73434 0 73490 800 0 FreeSans 224 90 0 0 io_wbs_sel[0]
port 294 nsew signal input
flabel metal2 s 74170 0 74226 800 0 FreeSans 224 90 0 0 io_wbs_sel[1]
port 295 nsew signal input
flabel metal2 s 74906 0 74962 800 0 FreeSans 224 90 0 0 io_wbs_sel[2]
port 296 nsew signal input
flabel metal2 s 75642 0 75698 800 0 FreeSans 224 90 0 0 io_wbs_sel[3]
port 297 nsew signal input
flabel metal3 s 79200 70864 80000 70984 0 FreeSans 480 0 0 0 io_wbs_sel_0[0]
port 298 nsew signal tristate
flabel metal3 s 79200 71544 80000 71664 0 FreeSans 480 0 0 0 io_wbs_sel_0[1]
port 299 nsew signal tristate
flabel metal3 s 79200 72224 80000 72344 0 FreeSans 480 0 0 0 io_wbs_sel_0[2]
port 300 nsew signal tristate
flabel metal3 s 79200 72904 80000 73024 0 FreeSans 480 0 0 0 io_wbs_sel_0[3]
port 301 nsew signal tristate
flabel metal3 s 0 70864 800 70984 0 FreeSans 480 0 0 0 io_wbs_sel_1[0]
port 302 nsew signal tristate
flabel metal3 s 0 71544 800 71664 0 FreeSans 480 0 0 0 io_wbs_sel_1[1]
port 303 nsew signal tristate
flabel metal3 s 0 72224 800 72344 0 FreeSans 480 0 0 0 io_wbs_sel_1[2]
port 304 nsew signal tristate
flabel metal3 s 0 72904 800 73024 0 FreeSans 480 0 0 0 io_wbs_sel_1[3]
port 305 nsew signal tristate
flabel metal2 s 76378 0 76434 800 0 FreeSans 224 90 0 0 io_wbs_stb
port 306 nsew signal input
flabel metal3 s 79200 73584 80000 73704 0 FreeSans 480 0 0 0 io_wbs_stb_0
port 307 nsew signal tristate
flabel metal3 s 0 73584 800 73704 0 FreeSans 480 0 0 0 io_wbs_stb_1
port 308 nsew signal tristate
flabel metal2 s 72698 0 72754 800 0 FreeSans 224 90 0 0 io_wbs_we
port 309 nsew signal input
flabel metal3 s 79200 70184 80000 70304 0 FreeSans 480 0 0 0 io_wbs_we_0
port 310 nsew signal tristate
flabel metal3 s 0 70184 800 70304 0 FreeSans 480 0 0 0 io_wbs_we_1
port 311 nsew signal tristate
flabel metal4 s 4208 2128 4528 77840 0 FreeSans 1920 90 0 0 vccd1
port 312 nsew power bidirectional
flabel metal4 s 34928 2128 35248 77840 0 FreeSans 1920 90 0 0 vccd1
port 312 nsew power bidirectional
flabel metal4 s 65648 2128 65968 77840 0 FreeSans 1920 90 0 0 vccd1
port 312 nsew power bidirectional
flabel metal4 s 19568 2128 19888 77840 0 FreeSans 1920 90 0 0 vssd1
port 313 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 77840 0 FreeSans 1920 90 0 0 vssd1
port 313 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>
