magic
tech sky130A
magscale 1 2
timestamp 1657014069
<< obsli1 >>
rect 1104 2159 78844 37553
<< obsm1 >>
rect 934 1912 79106 37584
<< metal2 >>
rect 938 39200 994 40000
rect 2778 39200 2834 40000
rect 4710 39200 4766 40000
rect 6642 39200 6698 40000
rect 8482 39200 8538 40000
rect 10414 39200 10470 40000
rect 12346 39200 12402 40000
rect 14278 39200 14334 40000
rect 16118 39200 16174 40000
rect 18050 39200 18106 40000
rect 19982 39200 20038 40000
rect 21822 39200 21878 40000
rect 23754 39200 23810 40000
rect 25686 39200 25742 40000
rect 27618 39200 27674 40000
rect 29458 39200 29514 40000
rect 31390 39200 31446 40000
rect 33322 39200 33378 40000
rect 35162 39200 35218 40000
rect 37094 39200 37150 40000
rect 39026 39200 39082 40000
rect 40958 39200 41014 40000
rect 42798 39200 42854 40000
rect 44730 39200 44786 40000
rect 46662 39200 46718 40000
rect 48502 39200 48558 40000
rect 50434 39200 50490 40000
rect 52366 39200 52422 40000
rect 54298 39200 54354 40000
rect 56138 39200 56194 40000
rect 58070 39200 58126 40000
rect 60002 39200 60058 40000
rect 61842 39200 61898 40000
rect 63774 39200 63830 40000
rect 65706 39200 65762 40000
rect 67638 39200 67694 40000
rect 69478 39200 69534 40000
rect 71410 39200 71466 40000
rect 73342 39200 73398 40000
rect 75182 39200 75238 40000
rect 77114 39200 77170 40000
rect 79046 39200 79102 40000
rect 938 0 994 800
rect 2778 0 2834 800
rect 4710 0 4766 800
rect 6642 0 6698 800
rect 8482 0 8538 800
rect 10414 0 10470 800
rect 12346 0 12402 800
rect 14278 0 14334 800
rect 16118 0 16174 800
rect 18050 0 18106 800
rect 19982 0 20038 800
rect 21822 0 21878 800
rect 23754 0 23810 800
rect 25686 0 25742 800
rect 27618 0 27674 800
rect 29458 0 29514 800
rect 31390 0 31446 800
rect 33322 0 33378 800
rect 35162 0 35218 800
rect 37094 0 37150 800
rect 39026 0 39082 800
rect 40958 0 41014 800
rect 42798 0 42854 800
rect 44730 0 44786 800
rect 46662 0 46718 800
rect 48502 0 48558 800
rect 50434 0 50490 800
rect 52366 0 52422 800
rect 54298 0 54354 800
rect 56138 0 56194 800
rect 58070 0 58126 800
rect 60002 0 60058 800
rect 61842 0 61898 800
rect 63774 0 63830 800
rect 65706 0 65762 800
rect 67638 0 67694 800
rect 69478 0 69534 800
rect 71410 0 71466 800
rect 73342 0 73398 800
rect 75182 0 75238 800
rect 77114 0 77170 800
rect 79046 0 79102 800
<< obsm2 >>
rect 1050 39144 2722 39545
rect 2890 39144 4654 39545
rect 4822 39144 6586 39545
rect 6754 39144 8426 39545
rect 8594 39144 10358 39545
rect 10526 39144 12290 39545
rect 12458 39144 14222 39545
rect 14390 39144 16062 39545
rect 16230 39144 17994 39545
rect 18162 39144 19926 39545
rect 20094 39144 21766 39545
rect 21934 39144 23698 39545
rect 23866 39144 25630 39545
rect 25798 39144 27562 39545
rect 27730 39144 29402 39545
rect 29570 39144 31334 39545
rect 31502 39144 33266 39545
rect 33434 39144 35106 39545
rect 35274 39144 37038 39545
rect 37206 39144 38970 39545
rect 39138 39144 40902 39545
rect 41070 39144 42742 39545
rect 42910 39144 44674 39545
rect 44842 39144 46606 39545
rect 46774 39144 48446 39545
rect 48614 39144 50378 39545
rect 50546 39144 52310 39545
rect 52478 39144 54242 39545
rect 54410 39144 56082 39545
rect 56250 39144 58014 39545
rect 58182 39144 59946 39545
rect 60114 39144 61786 39545
rect 61954 39144 63718 39545
rect 63886 39144 65650 39545
rect 65818 39144 67582 39545
rect 67750 39144 69422 39545
rect 69590 39144 71354 39545
rect 71522 39144 73286 39545
rect 73454 39144 75126 39545
rect 75294 39144 77058 39545
rect 77226 39144 78990 39545
rect 940 856 79100 39144
rect 1050 439 2722 856
rect 2890 439 4654 856
rect 4822 439 6586 856
rect 6754 439 8426 856
rect 8594 439 10358 856
rect 10526 439 12290 856
rect 12458 439 14222 856
rect 14390 439 16062 856
rect 16230 439 17994 856
rect 18162 439 19926 856
rect 20094 439 21766 856
rect 21934 439 23698 856
rect 23866 439 25630 856
rect 25798 439 27562 856
rect 27730 439 29402 856
rect 29570 439 31334 856
rect 31502 439 33266 856
rect 33434 439 35106 856
rect 35274 439 37038 856
rect 37206 439 38970 856
rect 39138 439 40902 856
rect 41070 439 42742 856
rect 42910 439 44674 856
rect 44842 439 46606 856
rect 46774 439 48446 856
rect 48614 439 50378 856
rect 50546 439 52310 856
rect 52478 439 54242 856
rect 54410 439 56082 856
rect 56250 439 58014 856
rect 58182 439 59946 856
rect 60114 439 61786 856
rect 61954 439 63718 856
rect 63886 439 65650 856
rect 65818 439 67582 856
rect 67750 439 69422 856
rect 69590 439 71354 856
rect 71522 439 73286 856
rect 73454 439 75126 856
rect 75294 439 77058 856
rect 77226 439 78990 856
<< metal3 >>
rect 79200 39448 80000 39568
rect 79200 38496 80000 38616
rect 79200 37544 80000 37664
rect 79200 36592 80000 36712
rect 79200 35640 80000 35760
rect 79200 34688 80000 34808
rect 79200 33872 80000 33992
rect 79200 32920 80000 33040
rect 79200 31968 80000 32088
rect 79200 31016 80000 31136
rect 79200 30064 80000 30184
rect 79200 29112 80000 29232
rect 79200 28296 80000 28416
rect 79200 27344 80000 27464
rect 79200 26392 80000 26512
rect 79200 25440 80000 25560
rect 79200 24488 80000 24608
rect 79200 23536 80000 23656
rect 79200 22720 80000 22840
rect 79200 21768 80000 21888
rect 79200 20816 80000 20936
rect 79200 19864 80000 19984
rect 79200 18912 80000 19032
rect 79200 17960 80000 18080
rect 79200 17144 80000 17264
rect 79200 16192 80000 16312
rect 79200 15240 80000 15360
rect 79200 14288 80000 14408
rect 79200 13336 80000 13456
rect 79200 12384 80000 12504
rect 79200 11568 80000 11688
rect 79200 10616 80000 10736
rect 79200 9664 80000 9784
rect 79200 8712 80000 8832
rect 79200 7760 80000 7880
rect 79200 6808 80000 6928
rect 79200 5992 80000 6112
rect 79200 5040 80000 5160
rect 79200 4088 80000 4208
rect 79200 3136 80000 3256
rect 79200 2184 80000 2304
rect 79200 1232 80000 1352
rect 79200 416 80000 536
<< obsm3 >>
rect 4208 39368 79120 39541
rect 4208 38696 79200 39368
rect 4208 38416 79120 38696
rect 4208 37744 79200 38416
rect 4208 37464 79120 37744
rect 4208 36792 79200 37464
rect 4208 36512 79120 36792
rect 4208 35840 79200 36512
rect 4208 35560 79120 35840
rect 4208 34888 79200 35560
rect 4208 34608 79120 34888
rect 4208 34072 79200 34608
rect 4208 33792 79120 34072
rect 4208 33120 79200 33792
rect 4208 32840 79120 33120
rect 4208 32168 79200 32840
rect 4208 31888 79120 32168
rect 4208 31216 79200 31888
rect 4208 30936 79120 31216
rect 4208 30264 79200 30936
rect 4208 29984 79120 30264
rect 4208 29312 79200 29984
rect 4208 29032 79120 29312
rect 4208 28496 79200 29032
rect 4208 28216 79120 28496
rect 4208 27544 79200 28216
rect 4208 27264 79120 27544
rect 4208 26592 79200 27264
rect 4208 26312 79120 26592
rect 4208 25640 79200 26312
rect 4208 25360 79120 25640
rect 4208 24688 79200 25360
rect 4208 24408 79120 24688
rect 4208 23736 79200 24408
rect 4208 23456 79120 23736
rect 4208 22920 79200 23456
rect 4208 22640 79120 22920
rect 4208 21968 79200 22640
rect 4208 21688 79120 21968
rect 4208 21016 79200 21688
rect 4208 20736 79120 21016
rect 4208 20064 79200 20736
rect 4208 19784 79120 20064
rect 4208 19112 79200 19784
rect 4208 18832 79120 19112
rect 4208 18160 79200 18832
rect 4208 17880 79120 18160
rect 4208 17344 79200 17880
rect 4208 17064 79120 17344
rect 4208 16392 79200 17064
rect 4208 16112 79120 16392
rect 4208 15440 79200 16112
rect 4208 15160 79120 15440
rect 4208 14488 79200 15160
rect 4208 14208 79120 14488
rect 4208 13536 79200 14208
rect 4208 13256 79120 13536
rect 4208 12584 79200 13256
rect 4208 12304 79120 12584
rect 4208 11768 79200 12304
rect 4208 11488 79120 11768
rect 4208 10816 79200 11488
rect 4208 10536 79120 10816
rect 4208 9864 79200 10536
rect 4208 9584 79120 9864
rect 4208 8912 79200 9584
rect 4208 8632 79120 8912
rect 4208 7960 79200 8632
rect 4208 7680 79120 7960
rect 4208 7008 79200 7680
rect 4208 6728 79120 7008
rect 4208 6192 79200 6728
rect 4208 5912 79120 6192
rect 4208 5240 79200 5912
rect 4208 4960 79120 5240
rect 4208 4288 79200 4960
rect 4208 4008 79120 4288
rect 4208 3336 79200 4008
rect 4208 3056 79120 3336
rect 4208 2384 79200 3056
rect 4208 2104 79120 2384
rect 4208 1432 79200 2104
rect 4208 1152 79120 1432
rect 4208 616 79200 1152
rect 4208 443 79120 616
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
rect 65648 2128 65968 37584
<< labels >>
rlabel metal3 s 79200 1232 80000 1352 6 addr[0]
port 1 nsew signal input
rlabel metal3 s 79200 2184 80000 2304 6 addr[1]
port 2 nsew signal input
rlabel metal3 s 79200 3136 80000 3256 6 addr[2]
port 3 nsew signal input
rlabel metal3 s 79200 4088 80000 4208 6 addr[3]
port 4 nsew signal input
rlabel metal3 s 79200 5040 80000 5160 6 addr[4]
port 5 nsew signal input
rlabel metal3 s 79200 5992 80000 6112 6 addr[5]
port 6 nsew signal input
rlabel metal3 s 79200 6808 80000 6928 6 addr[6]
port 7 nsew signal input
rlabel metal3 s 79200 7760 80000 7880 6 addr[7]
port 8 nsew signal input
rlabel metal3 s 79200 8712 80000 8832 6 addr[8]
port 9 nsew signal input
rlabel metal3 s 79200 9664 80000 9784 6 addr[9]
port 10 nsew signal input
rlabel metal2 s 2778 39200 2834 40000 6 addr_mem0[0]
port 11 nsew signal output
rlabel metal2 s 4710 39200 4766 40000 6 addr_mem0[1]
port 12 nsew signal output
rlabel metal2 s 6642 39200 6698 40000 6 addr_mem0[2]
port 13 nsew signal output
rlabel metal2 s 8482 39200 8538 40000 6 addr_mem0[3]
port 14 nsew signal output
rlabel metal2 s 10414 39200 10470 40000 6 addr_mem0[4]
port 15 nsew signal output
rlabel metal2 s 12346 39200 12402 40000 6 addr_mem0[5]
port 16 nsew signal output
rlabel metal2 s 14278 39200 14334 40000 6 addr_mem0[6]
port 17 nsew signal output
rlabel metal2 s 16118 39200 16174 40000 6 addr_mem0[7]
port 18 nsew signal output
rlabel metal2 s 18050 39200 18106 40000 6 addr_mem0[8]
port 19 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 addr_mem1[0]
port 20 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 addr_mem1[1]
port 21 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 addr_mem1[2]
port 22 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 addr_mem1[3]
port 23 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 addr_mem1[4]
port 24 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 addr_mem1[5]
port 25 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 addr_mem1[6]
port 26 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 addr_mem1[7]
port 27 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 addr_mem1[8]
port 28 nsew signal output
rlabel metal3 s 79200 416 80000 536 6 csb
port 29 nsew signal input
rlabel metal2 s 938 39200 994 40000 6 csb_mem0
port 30 nsew signal output
rlabel metal2 s 938 0 994 800 6 csb_mem1
port 31 nsew signal output
rlabel metal3 s 79200 10616 80000 10736 6 dout[0]
port 32 nsew signal output
rlabel metal3 s 79200 19864 80000 19984 6 dout[10]
port 33 nsew signal output
rlabel metal3 s 79200 20816 80000 20936 6 dout[11]
port 34 nsew signal output
rlabel metal3 s 79200 21768 80000 21888 6 dout[12]
port 35 nsew signal output
rlabel metal3 s 79200 22720 80000 22840 6 dout[13]
port 36 nsew signal output
rlabel metal3 s 79200 23536 80000 23656 6 dout[14]
port 37 nsew signal output
rlabel metal3 s 79200 24488 80000 24608 6 dout[15]
port 38 nsew signal output
rlabel metal3 s 79200 25440 80000 25560 6 dout[16]
port 39 nsew signal output
rlabel metal3 s 79200 26392 80000 26512 6 dout[17]
port 40 nsew signal output
rlabel metal3 s 79200 27344 80000 27464 6 dout[18]
port 41 nsew signal output
rlabel metal3 s 79200 28296 80000 28416 6 dout[19]
port 42 nsew signal output
rlabel metal3 s 79200 11568 80000 11688 6 dout[1]
port 43 nsew signal output
rlabel metal3 s 79200 29112 80000 29232 6 dout[20]
port 44 nsew signal output
rlabel metal3 s 79200 30064 80000 30184 6 dout[21]
port 45 nsew signal output
rlabel metal3 s 79200 31016 80000 31136 6 dout[22]
port 46 nsew signal output
rlabel metal3 s 79200 31968 80000 32088 6 dout[23]
port 47 nsew signal output
rlabel metal3 s 79200 32920 80000 33040 6 dout[24]
port 48 nsew signal output
rlabel metal3 s 79200 33872 80000 33992 6 dout[25]
port 49 nsew signal output
rlabel metal3 s 79200 34688 80000 34808 6 dout[26]
port 50 nsew signal output
rlabel metal3 s 79200 35640 80000 35760 6 dout[27]
port 51 nsew signal output
rlabel metal3 s 79200 36592 80000 36712 6 dout[28]
port 52 nsew signal output
rlabel metal3 s 79200 37544 80000 37664 6 dout[29]
port 53 nsew signal output
rlabel metal3 s 79200 12384 80000 12504 6 dout[2]
port 54 nsew signal output
rlabel metal3 s 79200 38496 80000 38616 6 dout[30]
port 55 nsew signal output
rlabel metal3 s 79200 39448 80000 39568 6 dout[31]
port 56 nsew signal output
rlabel metal3 s 79200 13336 80000 13456 6 dout[3]
port 57 nsew signal output
rlabel metal3 s 79200 14288 80000 14408 6 dout[4]
port 58 nsew signal output
rlabel metal3 s 79200 15240 80000 15360 6 dout[5]
port 59 nsew signal output
rlabel metal3 s 79200 16192 80000 16312 6 dout[6]
port 60 nsew signal output
rlabel metal3 s 79200 17144 80000 17264 6 dout[7]
port 61 nsew signal output
rlabel metal3 s 79200 17960 80000 18080 6 dout[8]
port 62 nsew signal output
rlabel metal3 s 79200 18912 80000 19032 6 dout[9]
port 63 nsew signal output
rlabel metal2 s 19982 39200 20038 40000 6 dout_mem0[0]
port 64 nsew signal input
rlabel metal2 s 39026 39200 39082 40000 6 dout_mem0[10]
port 65 nsew signal input
rlabel metal2 s 40958 39200 41014 40000 6 dout_mem0[11]
port 66 nsew signal input
rlabel metal2 s 42798 39200 42854 40000 6 dout_mem0[12]
port 67 nsew signal input
rlabel metal2 s 44730 39200 44786 40000 6 dout_mem0[13]
port 68 nsew signal input
rlabel metal2 s 46662 39200 46718 40000 6 dout_mem0[14]
port 69 nsew signal input
rlabel metal2 s 48502 39200 48558 40000 6 dout_mem0[15]
port 70 nsew signal input
rlabel metal2 s 50434 39200 50490 40000 6 dout_mem0[16]
port 71 nsew signal input
rlabel metal2 s 52366 39200 52422 40000 6 dout_mem0[17]
port 72 nsew signal input
rlabel metal2 s 54298 39200 54354 40000 6 dout_mem0[18]
port 73 nsew signal input
rlabel metal2 s 56138 39200 56194 40000 6 dout_mem0[19]
port 74 nsew signal input
rlabel metal2 s 21822 39200 21878 40000 6 dout_mem0[1]
port 75 nsew signal input
rlabel metal2 s 58070 39200 58126 40000 6 dout_mem0[20]
port 76 nsew signal input
rlabel metal2 s 60002 39200 60058 40000 6 dout_mem0[21]
port 77 nsew signal input
rlabel metal2 s 61842 39200 61898 40000 6 dout_mem0[22]
port 78 nsew signal input
rlabel metal2 s 63774 39200 63830 40000 6 dout_mem0[23]
port 79 nsew signal input
rlabel metal2 s 65706 39200 65762 40000 6 dout_mem0[24]
port 80 nsew signal input
rlabel metal2 s 67638 39200 67694 40000 6 dout_mem0[25]
port 81 nsew signal input
rlabel metal2 s 69478 39200 69534 40000 6 dout_mem0[26]
port 82 nsew signal input
rlabel metal2 s 71410 39200 71466 40000 6 dout_mem0[27]
port 83 nsew signal input
rlabel metal2 s 73342 39200 73398 40000 6 dout_mem0[28]
port 84 nsew signal input
rlabel metal2 s 75182 39200 75238 40000 6 dout_mem0[29]
port 85 nsew signal input
rlabel metal2 s 23754 39200 23810 40000 6 dout_mem0[2]
port 86 nsew signal input
rlabel metal2 s 77114 39200 77170 40000 6 dout_mem0[30]
port 87 nsew signal input
rlabel metal2 s 79046 39200 79102 40000 6 dout_mem0[31]
port 88 nsew signal input
rlabel metal2 s 25686 39200 25742 40000 6 dout_mem0[3]
port 89 nsew signal input
rlabel metal2 s 27618 39200 27674 40000 6 dout_mem0[4]
port 90 nsew signal input
rlabel metal2 s 29458 39200 29514 40000 6 dout_mem0[5]
port 91 nsew signal input
rlabel metal2 s 31390 39200 31446 40000 6 dout_mem0[6]
port 92 nsew signal input
rlabel metal2 s 33322 39200 33378 40000 6 dout_mem0[7]
port 93 nsew signal input
rlabel metal2 s 35162 39200 35218 40000 6 dout_mem0[8]
port 94 nsew signal input
rlabel metal2 s 37094 39200 37150 40000 6 dout_mem0[9]
port 95 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 dout_mem1[0]
port 96 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 dout_mem1[10]
port 97 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 dout_mem1[11]
port 98 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 dout_mem1[12]
port 99 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 dout_mem1[13]
port 100 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 dout_mem1[14]
port 101 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 dout_mem1[15]
port 102 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 dout_mem1[16]
port 103 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 dout_mem1[17]
port 104 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 dout_mem1[18]
port 105 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 dout_mem1[19]
port 106 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 dout_mem1[1]
port 107 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 dout_mem1[20]
port 108 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 dout_mem1[21]
port 109 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 dout_mem1[22]
port 110 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 dout_mem1[23]
port 111 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 dout_mem1[24]
port 112 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 dout_mem1[25]
port 113 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 dout_mem1[26]
port 114 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 dout_mem1[27]
port 115 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 dout_mem1[28]
port 116 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 dout_mem1[29]
port 117 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 dout_mem1[2]
port 118 nsew signal input
rlabel metal2 s 77114 0 77170 800 6 dout_mem1[30]
port 119 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 dout_mem1[31]
port 120 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 dout_mem1[3]
port 121 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 dout_mem1[4]
port 122 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 dout_mem1[5]
port 123 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 dout_mem1[6]
port 124 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 dout_mem1[7]
port 125 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 dout_mem1[8]
port 126 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 dout_mem1[9]
port 127 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 128 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 128 nsew power input
rlabel metal4 s 65648 2128 65968 37584 6 vccd1
port 128 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 129 nsew ground input
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 129 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 80000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1179284
string GDS_FILE /home/leo/Dokumente/caravel_workspace/caravel_wfg/openlane/merge_memory/runs/merge_memory/results/finishing/merge_memory.magic.gds
string GDS_START 81792
<< end >>

