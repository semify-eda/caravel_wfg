VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wfg_top
  CLASS BLOCK ;
  FOREIGN wfg_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 350.000 ;
  PIN addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END addr1[0]
  PIN addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END addr1[1]
  PIN addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END addr1[2]
  PIN addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END addr1[3]
  PIN addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END addr1[4]
  PIN addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END addr1[5]
  PIN addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END addr1[6]
  PIN addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END addr1[7]
  PIN addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END addr1[8]
  PIN addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END addr1[9]
  PIN csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END csb1
  PIN dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END dout1[0]
  PIN dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END dout1[10]
  PIN dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END dout1[11]
  PIN dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END dout1[12]
  PIN dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END dout1[13]
  PIN dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END dout1[14]
  PIN dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END dout1[15]
  PIN dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END dout1[16]
  PIN dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END dout1[17]
  PIN dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END dout1[18]
  PIN dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END dout1[19]
  PIN dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END dout1[1]
  PIN dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END dout1[20]
  PIN dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END dout1[21]
  PIN dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END dout1[22]
  PIN dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END dout1[23]
  PIN dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END dout1[24]
  PIN dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END dout1[25]
  PIN dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END dout1[26]
  PIN dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END dout1[27]
  PIN dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END dout1[28]
  PIN dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END dout1[29]
  PIN dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END dout1[2]
  PIN dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END dout1[30]
  PIN dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END dout1[31]
  PIN dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END dout1[3]
  PIN dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END dout1[4]
  PIN dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END dout1[5]
  PIN dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END dout1[6]
  PIN dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END dout1[7]
  PIN dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END dout1[8]
  PIN dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END dout1[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 346.000 463.130 350.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 346.000 593.310 350.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 346.000 476.010 350.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 346.000 488.890 350.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 346.000 502.230 350.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 346.000 515.110 350.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 346.000 527.990 350.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 346.000 541.330 350.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 346.000 554.210 350.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 346.000 567.090 350.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 346.000 580.430 350.000 ;
    END
  END io_oeb[9]
  PIN io_wbs_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END io_wbs_ack
  PIN io_wbs_adr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END io_wbs_adr[0]
  PIN io_wbs_adr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END io_wbs_adr[10]
  PIN io_wbs_adr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END io_wbs_adr[11]
  PIN io_wbs_adr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END io_wbs_adr[12]
  PIN io_wbs_adr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END io_wbs_adr[13]
  PIN io_wbs_adr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END io_wbs_adr[14]
  PIN io_wbs_adr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END io_wbs_adr[15]
  PIN io_wbs_adr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END io_wbs_adr[16]
  PIN io_wbs_adr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 0.000 338.010 4.000 ;
    END
  END io_wbs_adr[17]
  PIN io_wbs_adr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 0.000 355.950 4.000 ;
    END
  END io_wbs_adr[18]
  PIN io_wbs_adr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END io_wbs_adr[19]
  PIN io_wbs_adr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END io_wbs_adr[1]
  PIN io_wbs_adr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END io_wbs_adr[20]
  PIN io_wbs_adr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END io_wbs_adr[21]
  PIN io_wbs_adr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END io_wbs_adr[22]
  PIN io_wbs_adr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END io_wbs_adr[23]
  PIN io_wbs_adr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END io_wbs_adr[24]
  PIN io_wbs_adr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END io_wbs_adr[25]
  PIN io_wbs_adr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END io_wbs_adr[26]
  PIN io_wbs_adr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.370 0.000 514.650 4.000 ;
    END
  END io_wbs_adr[27]
  PIN io_wbs_adr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END io_wbs_adr[28]
  PIN io_wbs_adr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END io_wbs_adr[29]
  PIN io_wbs_adr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END io_wbs_adr[2]
  PIN io_wbs_adr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 0.000 567.550 4.000 ;
    END
  END io_wbs_adr[30]
  PIN io_wbs_adr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END io_wbs_adr[31]
  PIN io_wbs_adr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END io_wbs_adr[3]
  PIN io_wbs_adr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END io_wbs_adr[4]
  PIN io_wbs_adr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END io_wbs_adr[5]
  PIN io_wbs_adr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END io_wbs_adr[6]
  PIN io_wbs_adr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END io_wbs_adr[7]
  PIN io_wbs_adr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END io_wbs_adr[8]
  PIN io_wbs_adr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END io_wbs_adr[9]
  PIN io_wbs_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END io_wbs_clk
  PIN io_wbs_cyc
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END io_wbs_cyc
  PIN io_wbs_datrd[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END io_wbs_datrd[0]
  PIN io_wbs_datrd[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END io_wbs_datrd[10]
  PIN io_wbs_datrd[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END io_wbs_datrd[11]
  PIN io_wbs_datrd[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END io_wbs_datrd[12]
  PIN io_wbs_datrd[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END io_wbs_datrd[13]
  PIN io_wbs_datrd[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END io_wbs_datrd[14]
  PIN io_wbs_datrd[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END io_wbs_datrd[15]
  PIN io_wbs_datrd[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 0.000 326.510 4.000 ;
    END
  END io_wbs_datrd[16]
  PIN io_wbs_datrd[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END io_wbs_datrd[17]
  PIN io_wbs_datrd[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END io_wbs_datrd[18]
  PIN io_wbs_datrd[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END io_wbs_datrd[19]
  PIN io_wbs_datrd[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_wbs_datrd[1]
  PIN io_wbs_datrd[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END io_wbs_datrd[20]
  PIN io_wbs_datrd[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END io_wbs_datrd[21]
  PIN io_wbs_datrd[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END io_wbs_datrd[22]
  PIN io_wbs_datrd[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END io_wbs_datrd[23]
  PIN io_wbs_datrd[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END io_wbs_datrd[24]
  PIN io_wbs_datrd[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END io_wbs_datrd[25]
  PIN io_wbs_datrd[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END io_wbs_datrd[26]
  PIN io_wbs_datrd[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END io_wbs_datrd[27]
  PIN io_wbs_datrd[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END io_wbs_datrd[28]
  PIN io_wbs_datrd[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END io_wbs_datrd[29]
  PIN io_wbs_datrd[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END io_wbs_datrd[2]
  PIN io_wbs_datrd[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END io_wbs_datrd[30]
  PIN io_wbs_datrd[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END io_wbs_datrd[31]
  PIN io_wbs_datrd[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_wbs_datrd[3]
  PIN io_wbs_datrd[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END io_wbs_datrd[4]
  PIN io_wbs_datrd[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END io_wbs_datrd[5]
  PIN io_wbs_datrd[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END io_wbs_datrd[6]
  PIN io_wbs_datrd[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END io_wbs_datrd[7]
  PIN io_wbs_datrd[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END io_wbs_datrd[8]
  PIN io_wbs_datrd[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END io_wbs_datrd[9]
  PIN io_wbs_datwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END io_wbs_datwr[0]
  PIN io_wbs_datwr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END io_wbs_datwr[10]
  PIN io_wbs_datwr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END io_wbs_datwr[11]
  PIN io_wbs_datwr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END io_wbs_datwr[12]
  PIN io_wbs_datwr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END io_wbs_datwr[13]
  PIN io_wbs_datwr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END io_wbs_datwr[14]
  PIN io_wbs_datwr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END io_wbs_datwr[15]
  PIN io_wbs_datwr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END io_wbs_datwr[16]
  PIN io_wbs_datwr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END io_wbs_datwr[17]
  PIN io_wbs_datwr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END io_wbs_datwr[18]
  PIN io_wbs_datwr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 0.000 384.930 4.000 ;
    END
  END io_wbs_datwr[19]
  PIN io_wbs_datwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END io_wbs_datwr[1]
  PIN io_wbs_datwr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END io_wbs_datwr[20]
  PIN io_wbs_datwr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END io_wbs_datwr[21]
  PIN io_wbs_datwr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END io_wbs_datwr[22]
  PIN io_wbs_datwr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END io_wbs_datwr[23]
  PIN io_wbs_datwr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END io_wbs_datwr[24]
  PIN io_wbs_datwr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END io_wbs_datwr[25]
  PIN io_wbs_datwr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END io_wbs_datwr[26]
  PIN io_wbs_datwr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 4.000 ;
    END
  END io_wbs_datwr[27]
  PIN io_wbs_datwr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END io_wbs_datwr[28]
  PIN io_wbs_datwr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END io_wbs_datwr[29]
  PIN io_wbs_datwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END io_wbs_datwr[2]
  PIN io_wbs_datwr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END io_wbs_datwr[30]
  PIN io_wbs_datwr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END io_wbs_datwr[31]
  PIN io_wbs_datwr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END io_wbs_datwr[3]
  PIN io_wbs_datwr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END io_wbs_datwr[4]
  PIN io_wbs_datwr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END io_wbs_datwr[5]
  PIN io_wbs_datwr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END io_wbs_datwr[6]
  PIN io_wbs_datwr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END io_wbs_datwr[7]
  PIN io_wbs_datwr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END io_wbs_datwr[8]
  PIN io_wbs_datwr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END io_wbs_datwr[9]
  PIN io_wbs_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 4.000 ;
    END
  END io_wbs_rst
  PIN io_wbs_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END io_wbs_stb
  PIN io_wbs_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END io_wbs_we
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 337.520 ;
    END
  END vssd1
  PIN wfg_drive_pat_dout_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 346.000 45.910 350.000 ;
    END
  END wfg_drive_pat_dout_o[0]
  PIN wfg_drive_pat_dout_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 346.000 176.090 350.000 ;
    END
  END wfg_drive_pat_dout_o[10]
  PIN wfg_drive_pat_dout_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 346.000 188.970 350.000 ;
    END
  END wfg_drive_pat_dout_o[11]
  PIN wfg_drive_pat_dout_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 346.000 202.310 350.000 ;
    END
  END wfg_drive_pat_dout_o[12]
  PIN wfg_drive_pat_dout_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 346.000 215.190 350.000 ;
    END
  END wfg_drive_pat_dout_o[13]
  PIN wfg_drive_pat_dout_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 346.000 228.070 350.000 ;
    END
  END wfg_drive_pat_dout_o[14]
  PIN wfg_drive_pat_dout_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 346.000 241.410 350.000 ;
    END
  END wfg_drive_pat_dout_o[15]
  PIN wfg_drive_pat_dout_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 346.000 254.290 350.000 ;
    END
  END wfg_drive_pat_dout_o[16]
  PIN wfg_drive_pat_dout_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 346.000 267.170 350.000 ;
    END
  END wfg_drive_pat_dout_o[17]
  PIN wfg_drive_pat_dout_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 346.000 280.510 350.000 ;
    END
  END wfg_drive_pat_dout_o[18]
  PIN wfg_drive_pat_dout_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 346.000 293.390 350.000 ;
    END
  END wfg_drive_pat_dout_o[19]
  PIN wfg_drive_pat_dout_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 346.000 58.790 350.000 ;
    END
  END wfg_drive_pat_dout_o[1]
  PIN wfg_drive_pat_dout_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 346.000 306.730 350.000 ;
    END
  END wfg_drive_pat_dout_o[20]
  PIN wfg_drive_pat_dout_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 346.000 319.610 350.000 ;
    END
  END wfg_drive_pat_dout_o[21]
  PIN wfg_drive_pat_dout_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 346.000 332.490 350.000 ;
    END
  END wfg_drive_pat_dout_o[22]
  PIN wfg_drive_pat_dout_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 346.000 345.830 350.000 ;
    END
  END wfg_drive_pat_dout_o[23]
  PIN wfg_drive_pat_dout_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 346.000 358.710 350.000 ;
    END
  END wfg_drive_pat_dout_o[24]
  PIN wfg_drive_pat_dout_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 346.000 371.590 350.000 ;
    END
  END wfg_drive_pat_dout_o[25]
  PIN wfg_drive_pat_dout_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.650 346.000 384.930 350.000 ;
    END
  END wfg_drive_pat_dout_o[26]
  PIN wfg_drive_pat_dout_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 346.000 397.810 350.000 ;
    END
  END wfg_drive_pat_dout_o[27]
  PIN wfg_drive_pat_dout_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.410 346.000 410.690 350.000 ;
    END
  END wfg_drive_pat_dout_o[28]
  PIN wfg_drive_pat_dout_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 346.000 424.030 350.000 ;
    END
  END wfg_drive_pat_dout_o[29]
  PIN wfg_drive_pat_dout_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 346.000 71.670 350.000 ;
    END
  END wfg_drive_pat_dout_o[2]
  PIN wfg_drive_pat_dout_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 346.000 436.910 350.000 ;
    END
  END wfg_drive_pat_dout_o[30]
  PIN wfg_drive_pat_dout_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 346.000 449.790 350.000 ;
    END
  END wfg_drive_pat_dout_o[31]
  PIN wfg_drive_pat_dout_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 346.000 85.010 350.000 ;
    END
  END wfg_drive_pat_dout_o[3]
  PIN wfg_drive_pat_dout_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 346.000 97.890 350.000 ;
    END
  END wfg_drive_pat_dout_o[4]
  PIN wfg_drive_pat_dout_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 346.000 110.770 350.000 ;
    END
  END wfg_drive_pat_dout_o[5]
  PIN wfg_drive_pat_dout_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 346.000 124.110 350.000 ;
    END
  END wfg_drive_pat_dout_o[6]
  PIN wfg_drive_pat_dout_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 346.000 136.990 350.000 ;
    END
  END wfg_drive_pat_dout_o[7]
  PIN wfg_drive_pat_dout_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 346.000 149.870 350.000 ;
    END
  END wfg_drive_pat_dout_o[8]
  PIN wfg_drive_pat_dout_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 346.000 163.210 350.000 ;
    END
  END wfg_drive_pat_dout_o[9]
  PIN wfg_drive_spi_cs_no
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 346.000 6.810 350.000 ;
    END
  END wfg_drive_spi_cs_no
  PIN wfg_drive_spi_sclk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 346.000 19.690 350.000 ;
    END
  END wfg_drive_spi_sclk_o
  PIN wfg_drive_spi_sdo_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 346.000 32.570 350.000 ;
    END
  END wfg_drive_spi_sdo_o
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 337.365 ;
      LAYER met1 ;
        RECT 2.830 0.040 597.010 337.920 ;
      LAYER met2 ;
        RECT 2.860 345.720 6.250 346.530 ;
        RECT 7.090 345.720 19.130 346.530 ;
        RECT 19.970 345.720 32.010 346.530 ;
        RECT 32.850 345.720 45.350 346.530 ;
        RECT 46.190 345.720 58.230 346.530 ;
        RECT 59.070 345.720 71.110 346.530 ;
        RECT 71.950 345.720 84.450 346.530 ;
        RECT 85.290 345.720 97.330 346.530 ;
        RECT 98.170 345.720 110.210 346.530 ;
        RECT 111.050 345.720 123.550 346.530 ;
        RECT 124.390 345.720 136.430 346.530 ;
        RECT 137.270 345.720 149.310 346.530 ;
        RECT 150.150 345.720 162.650 346.530 ;
        RECT 163.490 345.720 175.530 346.530 ;
        RECT 176.370 345.720 188.410 346.530 ;
        RECT 189.250 345.720 201.750 346.530 ;
        RECT 202.590 345.720 214.630 346.530 ;
        RECT 215.470 345.720 227.510 346.530 ;
        RECT 228.350 345.720 240.850 346.530 ;
        RECT 241.690 345.720 253.730 346.530 ;
        RECT 254.570 345.720 266.610 346.530 ;
        RECT 267.450 345.720 279.950 346.530 ;
        RECT 280.790 345.720 292.830 346.530 ;
        RECT 293.670 345.720 306.170 346.530 ;
        RECT 307.010 345.720 319.050 346.530 ;
        RECT 319.890 345.720 331.930 346.530 ;
        RECT 332.770 345.720 345.270 346.530 ;
        RECT 346.110 345.720 358.150 346.530 ;
        RECT 358.990 345.720 371.030 346.530 ;
        RECT 371.870 345.720 384.370 346.530 ;
        RECT 385.210 345.720 397.250 346.530 ;
        RECT 398.090 345.720 410.130 346.530 ;
        RECT 410.970 345.720 423.470 346.530 ;
        RECT 424.310 345.720 436.350 346.530 ;
        RECT 437.190 345.720 449.230 346.530 ;
        RECT 450.070 345.720 462.570 346.530 ;
        RECT 463.410 345.720 475.450 346.530 ;
        RECT 476.290 345.720 488.330 346.530 ;
        RECT 489.170 345.720 501.670 346.530 ;
        RECT 502.510 345.720 514.550 346.530 ;
        RECT 515.390 345.720 527.430 346.530 ;
        RECT 528.270 345.720 540.770 346.530 ;
        RECT 541.610 345.720 553.650 346.530 ;
        RECT 554.490 345.720 566.530 346.530 ;
        RECT 567.370 345.720 579.870 346.530 ;
        RECT 580.710 345.720 592.750 346.530 ;
        RECT 593.590 345.720 596.980 346.530 ;
        RECT 2.860 4.280 596.980 345.720 ;
        RECT 3.410 0.010 8.090 4.280 ;
        RECT 8.930 0.010 14.070 4.280 ;
        RECT 14.910 0.010 20.050 4.280 ;
        RECT 20.890 0.010 26.030 4.280 ;
        RECT 26.870 0.010 31.550 4.280 ;
        RECT 32.390 0.010 37.530 4.280 ;
        RECT 38.370 0.010 43.510 4.280 ;
        RECT 44.350 0.010 49.490 4.280 ;
        RECT 50.330 0.010 55.470 4.280 ;
        RECT 56.310 0.010 60.990 4.280 ;
        RECT 61.830 0.010 66.970 4.280 ;
        RECT 67.810 0.010 72.950 4.280 ;
        RECT 73.790 0.010 78.930 4.280 ;
        RECT 79.770 0.010 84.450 4.280 ;
        RECT 85.290 0.010 90.430 4.280 ;
        RECT 91.270 0.010 96.410 4.280 ;
        RECT 97.250 0.010 102.390 4.280 ;
        RECT 103.230 0.010 108.370 4.280 ;
        RECT 109.210 0.010 113.890 4.280 ;
        RECT 114.730 0.010 119.870 4.280 ;
        RECT 120.710 0.010 125.850 4.280 ;
        RECT 126.690 0.010 131.830 4.280 ;
        RECT 132.670 0.010 137.810 4.280 ;
        RECT 138.650 0.010 143.330 4.280 ;
        RECT 144.170 0.010 149.310 4.280 ;
        RECT 150.150 0.010 155.290 4.280 ;
        RECT 156.130 0.010 161.270 4.280 ;
        RECT 162.110 0.010 166.790 4.280 ;
        RECT 167.630 0.010 172.770 4.280 ;
        RECT 173.610 0.010 178.750 4.280 ;
        RECT 179.590 0.010 184.730 4.280 ;
        RECT 185.570 0.010 190.710 4.280 ;
        RECT 191.550 0.010 196.230 4.280 ;
        RECT 197.070 0.010 202.210 4.280 ;
        RECT 203.050 0.010 208.190 4.280 ;
        RECT 209.030 0.010 214.170 4.280 ;
        RECT 215.010 0.010 220.150 4.280 ;
        RECT 220.990 0.010 225.670 4.280 ;
        RECT 226.510 0.010 231.650 4.280 ;
        RECT 232.490 0.010 237.630 4.280 ;
        RECT 238.470 0.010 243.610 4.280 ;
        RECT 244.450 0.010 249.130 4.280 ;
        RECT 249.970 0.010 255.110 4.280 ;
        RECT 255.950 0.010 261.090 4.280 ;
        RECT 261.930 0.010 267.070 4.280 ;
        RECT 267.910 0.010 273.050 4.280 ;
        RECT 273.890 0.010 278.570 4.280 ;
        RECT 279.410 0.010 284.550 4.280 ;
        RECT 285.390 0.010 290.530 4.280 ;
        RECT 291.370 0.010 296.510 4.280 ;
        RECT 297.350 0.010 302.490 4.280 ;
        RECT 303.330 0.010 308.010 4.280 ;
        RECT 308.850 0.010 313.990 4.280 ;
        RECT 314.830 0.010 319.970 4.280 ;
        RECT 320.810 0.010 325.950 4.280 ;
        RECT 326.790 0.010 331.470 4.280 ;
        RECT 332.310 0.010 337.450 4.280 ;
        RECT 338.290 0.010 343.430 4.280 ;
        RECT 344.270 0.010 349.410 4.280 ;
        RECT 350.250 0.010 355.390 4.280 ;
        RECT 356.230 0.010 360.910 4.280 ;
        RECT 361.750 0.010 366.890 4.280 ;
        RECT 367.730 0.010 372.870 4.280 ;
        RECT 373.710 0.010 378.850 4.280 ;
        RECT 379.690 0.010 384.370 4.280 ;
        RECT 385.210 0.010 390.350 4.280 ;
        RECT 391.190 0.010 396.330 4.280 ;
        RECT 397.170 0.010 402.310 4.280 ;
        RECT 403.150 0.010 408.290 4.280 ;
        RECT 409.130 0.010 413.810 4.280 ;
        RECT 414.650 0.010 419.790 4.280 ;
        RECT 420.630 0.010 425.770 4.280 ;
        RECT 426.610 0.010 431.750 4.280 ;
        RECT 432.590 0.010 437.730 4.280 ;
        RECT 438.570 0.010 443.250 4.280 ;
        RECT 444.090 0.010 449.230 4.280 ;
        RECT 450.070 0.010 455.210 4.280 ;
        RECT 456.050 0.010 461.190 4.280 ;
        RECT 462.030 0.010 466.710 4.280 ;
        RECT 467.550 0.010 472.690 4.280 ;
        RECT 473.530 0.010 478.670 4.280 ;
        RECT 479.510 0.010 484.650 4.280 ;
        RECT 485.490 0.010 490.630 4.280 ;
        RECT 491.470 0.010 496.150 4.280 ;
        RECT 496.990 0.010 502.130 4.280 ;
        RECT 502.970 0.010 508.110 4.280 ;
        RECT 508.950 0.010 514.090 4.280 ;
        RECT 514.930 0.010 520.070 4.280 ;
        RECT 520.910 0.010 525.590 4.280 ;
        RECT 526.430 0.010 531.570 4.280 ;
        RECT 532.410 0.010 537.550 4.280 ;
        RECT 538.390 0.010 543.530 4.280 ;
        RECT 544.370 0.010 549.050 4.280 ;
        RECT 549.890 0.010 555.030 4.280 ;
        RECT 555.870 0.010 561.010 4.280 ;
        RECT 561.850 0.010 566.990 4.280 ;
        RECT 567.830 0.010 572.970 4.280 ;
        RECT 573.810 0.010 578.490 4.280 ;
        RECT 579.330 0.010 584.470 4.280 ;
        RECT 585.310 0.010 590.450 4.280 ;
        RECT 591.290 0.010 596.430 4.280 ;
      LAYER met3 ;
        RECT 4.400 345.080 580.915 345.945 ;
        RECT 4.000 338.320 580.915 345.080 ;
        RECT 4.400 336.920 580.915 338.320 ;
        RECT 4.000 330.160 580.915 336.920 ;
        RECT 4.400 328.760 580.915 330.160 ;
        RECT 4.000 322.000 580.915 328.760 ;
        RECT 4.400 320.600 580.915 322.000 ;
        RECT 4.000 313.840 580.915 320.600 ;
        RECT 4.400 312.440 580.915 313.840 ;
        RECT 4.000 305.680 580.915 312.440 ;
        RECT 4.400 304.280 580.915 305.680 ;
        RECT 4.000 297.520 580.915 304.280 ;
        RECT 4.400 296.120 580.915 297.520 ;
        RECT 4.000 289.360 580.915 296.120 ;
        RECT 4.400 287.960 580.915 289.360 ;
        RECT 4.000 281.200 580.915 287.960 ;
        RECT 4.400 279.800 580.915 281.200 ;
        RECT 4.000 273.040 580.915 279.800 ;
        RECT 4.400 271.640 580.915 273.040 ;
        RECT 4.000 264.880 580.915 271.640 ;
        RECT 4.400 263.480 580.915 264.880 ;
        RECT 4.000 256.720 580.915 263.480 ;
        RECT 4.400 255.320 580.915 256.720 ;
        RECT 4.000 248.560 580.915 255.320 ;
        RECT 4.400 247.160 580.915 248.560 ;
        RECT 4.000 240.400 580.915 247.160 ;
        RECT 4.400 239.000 580.915 240.400 ;
        RECT 4.000 232.240 580.915 239.000 ;
        RECT 4.400 230.840 580.915 232.240 ;
        RECT 4.000 224.080 580.915 230.840 ;
        RECT 4.400 222.680 580.915 224.080 ;
        RECT 4.000 215.920 580.915 222.680 ;
        RECT 4.400 214.520 580.915 215.920 ;
        RECT 4.000 207.760 580.915 214.520 ;
        RECT 4.400 206.360 580.915 207.760 ;
        RECT 4.000 199.600 580.915 206.360 ;
        RECT 4.400 198.200 580.915 199.600 ;
        RECT 4.000 191.440 580.915 198.200 ;
        RECT 4.400 190.040 580.915 191.440 ;
        RECT 4.000 183.280 580.915 190.040 ;
        RECT 4.400 181.880 580.915 183.280 ;
        RECT 4.000 175.120 580.915 181.880 ;
        RECT 4.400 173.720 580.915 175.120 ;
        RECT 4.000 166.960 580.915 173.720 ;
        RECT 4.400 165.560 580.915 166.960 ;
        RECT 4.000 158.800 580.915 165.560 ;
        RECT 4.400 157.400 580.915 158.800 ;
        RECT 4.000 150.640 580.915 157.400 ;
        RECT 4.400 149.240 580.915 150.640 ;
        RECT 4.000 142.480 580.915 149.240 ;
        RECT 4.400 141.080 580.915 142.480 ;
        RECT 4.000 134.320 580.915 141.080 ;
        RECT 4.400 132.920 580.915 134.320 ;
        RECT 4.000 126.160 580.915 132.920 ;
        RECT 4.400 124.760 580.915 126.160 ;
        RECT 4.000 118.000 580.915 124.760 ;
        RECT 4.400 116.600 580.915 118.000 ;
        RECT 4.000 109.840 580.915 116.600 ;
        RECT 4.400 108.440 580.915 109.840 ;
        RECT 4.000 101.680 580.915 108.440 ;
        RECT 4.400 100.280 580.915 101.680 ;
        RECT 4.000 93.520 580.915 100.280 ;
        RECT 4.400 92.120 580.915 93.520 ;
        RECT 4.000 85.360 580.915 92.120 ;
        RECT 4.400 83.960 580.915 85.360 ;
        RECT 4.000 77.200 580.915 83.960 ;
        RECT 4.400 75.800 580.915 77.200 ;
        RECT 4.000 69.040 580.915 75.800 ;
        RECT 4.400 67.640 580.915 69.040 ;
        RECT 4.000 60.880 580.915 67.640 ;
        RECT 4.400 59.480 580.915 60.880 ;
        RECT 4.000 52.720 580.915 59.480 ;
        RECT 4.400 51.320 580.915 52.720 ;
        RECT 4.000 44.560 580.915 51.320 ;
        RECT 4.400 43.160 580.915 44.560 ;
        RECT 4.000 36.400 580.915 43.160 ;
        RECT 4.400 35.000 580.915 36.400 ;
        RECT 4.000 28.240 580.915 35.000 ;
        RECT 4.400 26.840 580.915 28.240 ;
        RECT 4.000 20.080 580.915 26.840 ;
        RECT 4.400 18.680 580.915 20.080 ;
        RECT 4.000 11.920 580.915 18.680 ;
        RECT 4.400 10.520 580.915 11.920 ;
        RECT 4.000 4.440 580.915 10.520 ;
        RECT 4.400 3.575 580.915 4.440 ;
      LAYER met4 ;
        RECT 96.895 22.615 97.440 336.425 ;
        RECT 99.840 22.615 174.240 336.425 ;
        RECT 176.640 22.615 251.040 336.425 ;
        RECT 253.440 22.615 327.840 336.425 ;
        RECT 330.240 22.615 404.640 336.425 ;
        RECT 407.040 22.615 481.440 336.425 ;
        RECT 483.840 22.615 516.745 336.425 ;
  END
END wfg_top
END LIBRARY

