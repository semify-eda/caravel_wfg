magic
tech sky130A
magscale 1 2
timestamp 1657525571
<< obsli1 >>
rect 1104 2159 148856 107729
<< obsm1 >>
rect 1104 1640 148856 107840
<< metal2 >>
rect 2502 109200 2558 110000
rect 5722 109200 5778 110000
rect 8942 109200 8998 110000
rect 12162 109200 12218 110000
rect 15382 109200 15438 110000
rect 18602 109200 18658 110000
rect 21822 109200 21878 110000
rect 25042 109200 25098 110000
rect 28262 109200 28318 110000
rect 31482 109200 31538 110000
rect 34702 109200 34758 110000
rect 37922 109200 37978 110000
rect 41142 109200 41198 110000
rect 44362 109200 44418 110000
rect 47582 109200 47638 110000
rect 50802 109200 50858 110000
rect 54022 109200 54078 110000
rect 57242 109200 57298 110000
rect 60462 109200 60518 110000
rect 63682 109200 63738 110000
rect 66902 109200 66958 110000
rect 70122 109200 70178 110000
rect 73342 109200 73398 110000
rect 76562 109200 76618 110000
rect 79782 109200 79838 110000
rect 83002 109200 83058 110000
rect 86222 109200 86278 110000
rect 89442 109200 89498 110000
rect 92662 109200 92718 110000
rect 95882 109200 95938 110000
rect 99102 109200 99158 110000
rect 102322 109200 102378 110000
rect 105542 109200 105598 110000
rect 108762 109200 108818 110000
rect 111982 109200 112038 110000
rect 115202 109200 115258 110000
rect 118422 109200 118478 110000
rect 121642 109200 121698 110000
rect 124862 109200 124918 110000
rect 128082 109200 128138 110000
rect 131302 109200 131358 110000
rect 134522 109200 134578 110000
rect 137742 109200 137798 110000
rect 140962 109200 141018 110000
rect 144182 109200 144238 110000
rect 147402 109200 147458 110000
rect 5262 0 5318 800
rect 6642 0 6698 800
rect 8022 0 8078 800
rect 9402 0 9458 800
rect 10782 0 10838 800
rect 12162 0 12218 800
rect 13542 0 13598 800
rect 14922 0 14978 800
rect 16302 0 16358 800
rect 17682 0 17738 800
rect 19062 0 19118 800
rect 20442 0 20498 800
rect 21822 0 21878 800
rect 23202 0 23258 800
rect 24582 0 24638 800
rect 25962 0 26018 800
rect 27342 0 27398 800
rect 28722 0 28778 800
rect 30102 0 30158 800
rect 31482 0 31538 800
rect 32862 0 32918 800
rect 34242 0 34298 800
rect 35622 0 35678 800
rect 37002 0 37058 800
rect 38382 0 38438 800
rect 39762 0 39818 800
rect 41142 0 41198 800
rect 42522 0 42578 800
rect 43902 0 43958 800
rect 45282 0 45338 800
rect 46662 0 46718 800
rect 48042 0 48098 800
rect 49422 0 49478 800
rect 50802 0 50858 800
rect 52182 0 52238 800
rect 53562 0 53618 800
rect 54942 0 54998 800
rect 56322 0 56378 800
rect 57702 0 57758 800
rect 59082 0 59138 800
rect 60462 0 60518 800
rect 61842 0 61898 800
rect 63222 0 63278 800
rect 64602 0 64658 800
rect 65982 0 66038 800
rect 67362 0 67418 800
rect 68742 0 68798 800
rect 70122 0 70178 800
rect 71502 0 71558 800
rect 72882 0 72938 800
rect 74262 0 74318 800
rect 75642 0 75698 800
rect 77022 0 77078 800
rect 78402 0 78458 800
rect 79782 0 79838 800
rect 81162 0 81218 800
rect 82542 0 82598 800
rect 83922 0 83978 800
rect 85302 0 85358 800
rect 86682 0 86738 800
rect 88062 0 88118 800
rect 89442 0 89498 800
rect 90822 0 90878 800
rect 92202 0 92258 800
rect 93582 0 93638 800
rect 94962 0 95018 800
rect 96342 0 96398 800
rect 97722 0 97778 800
rect 99102 0 99158 800
rect 100482 0 100538 800
rect 101862 0 101918 800
rect 103242 0 103298 800
rect 104622 0 104678 800
rect 106002 0 106058 800
rect 107382 0 107438 800
rect 108762 0 108818 800
rect 110142 0 110198 800
rect 111522 0 111578 800
rect 112902 0 112958 800
rect 114282 0 114338 800
rect 115662 0 115718 800
rect 117042 0 117098 800
rect 118422 0 118478 800
rect 119802 0 119858 800
rect 121182 0 121238 800
rect 122562 0 122618 800
rect 123942 0 123998 800
rect 125322 0 125378 800
rect 126702 0 126758 800
rect 128082 0 128138 800
rect 129462 0 129518 800
rect 130842 0 130898 800
rect 132222 0 132278 800
rect 133602 0 133658 800
rect 134982 0 135038 800
rect 136362 0 136418 800
rect 137742 0 137798 800
rect 139122 0 139178 800
rect 140502 0 140558 800
rect 141882 0 141938 800
rect 143262 0 143318 800
rect 144642 0 144698 800
<< obsm2 >>
rect 1398 109144 2446 109200
rect 2614 109144 5666 109200
rect 5834 109144 8886 109200
rect 9054 109144 12106 109200
rect 12274 109144 15326 109200
rect 15494 109144 18546 109200
rect 18714 109144 21766 109200
rect 21934 109144 24986 109200
rect 25154 109144 28206 109200
rect 28374 109144 31426 109200
rect 31594 109144 34646 109200
rect 34814 109144 37866 109200
rect 38034 109144 41086 109200
rect 41254 109144 44306 109200
rect 44474 109144 47526 109200
rect 47694 109144 50746 109200
rect 50914 109144 53966 109200
rect 54134 109144 57186 109200
rect 57354 109144 60406 109200
rect 60574 109144 63626 109200
rect 63794 109144 66846 109200
rect 67014 109144 70066 109200
rect 70234 109144 73286 109200
rect 73454 109144 76506 109200
rect 76674 109144 79726 109200
rect 79894 109144 82946 109200
rect 83114 109144 86166 109200
rect 86334 109144 89386 109200
rect 89554 109144 92606 109200
rect 92774 109144 95826 109200
rect 95994 109144 99046 109200
rect 99214 109144 102266 109200
rect 102434 109144 105486 109200
rect 105654 109144 108706 109200
rect 108874 109144 111926 109200
rect 112094 109144 115146 109200
rect 115314 109144 118366 109200
rect 118534 109144 121586 109200
rect 121754 109144 124806 109200
rect 124974 109144 128026 109200
rect 128194 109144 131246 109200
rect 131414 109144 134466 109200
rect 134634 109144 137686 109200
rect 137854 109144 140906 109200
rect 141074 109144 144126 109200
rect 144294 109144 147346 109200
rect 147514 109144 148008 109200
rect 1398 856 148008 109144
rect 1398 800 5206 856
rect 5374 800 6586 856
rect 6754 800 7966 856
rect 8134 800 9346 856
rect 9514 800 10726 856
rect 10894 800 12106 856
rect 12274 800 13486 856
rect 13654 800 14866 856
rect 15034 800 16246 856
rect 16414 800 17626 856
rect 17794 800 19006 856
rect 19174 800 20386 856
rect 20554 800 21766 856
rect 21934 800 23146 856
rect 23314 800 24526 856
rect 24694 800 25906 856
rect 26074 800 27286 856
rect 27454 800 28666 856
rect 28834 800 30046 856
rect 30214 800 31426 856
rect 31594 800 32806 856
rect 32974 800 34186 856
rect 34354 800 35566 856
rect 35734 800 36946 856
rect 37114 800 38326 856
rect 38494 800 39706 856
rect 39874 800 41086 856
rect 41254 800 42466 856
rect 42634 800 43846 856
rect 44014 800 45226 856
rect 45394 800 46606 856
rect 46774 800 47986 856
rect 48154 800 49366 856
rect 49534 800 50746 856
rect 50914 800 52126 856
rect 52294 800 53506 856
rect 53674 800 54886 856
rect 55054 800 56266 856
rect 56434 800 57646 856
rect 57814 800 59026 856
rect 59194 800 60406 856
rect 60574 800 61786 856
rect 61954 800 63166 856
rect 63334 800 64546 856
rect 64714 800 65926 856
rect 66094 800 67306 856
rect 67474 800 68686 856
rect 68854 800 70066 856
rect 70234 800 71446 856
rect 71614 800 72826 856
rect 72994 800 74206 856
rect 74374 800 75586 856
rect 75754 800 76966 856
rect 77134 800 78346 856
rect 78514 800 79726 856
rect 79894 800 81106 856
rect 81274 800 82486 856
rect 82654 800 83866 856
rect 84034 800 85246 856
rect 85414 800 86626 856
rect 86794 800 88006 856
rect 88174 800 89386 856
rect 89554 800 90766 856
rect 90934 800 92146 856
rect 92314 800 93526 856
rect 93694 800 94906 856
rect 95074 800 96286 856
rect 96454 800 97666 856
rect 97834 800 99046 856
rect 99214 800 100426 856
rect 100594 800 101806 856
rect 101974 800 103186 856
rect 103354 800 104566 856
rect 104734 800 105946 856
rect 106114 800 107326 856
rect 107494 800 108706 856
rect 108874 800 110086 856
rect 110254 800 111466 856
rect 111634 800 112846 856
rect 113014 800 114226 856
rect 114394 800 115606 856
rect 115774 800 116986 856
rect 117154 800 118366 856
rect 118534 800 119746 856
rect 119914 800 121126 856
rect 121294 800 122506 856
rect 122674 800 123886 856
rect 124054 800 125266 856
rect 125434 800 126646 856
rect 126814 800 128026 856
rect 128194 800 129406 856
rect 129574 800 130786 856
rect 130954 800 132166 856
rect 132334 800 133546 856
rect 133714 800 134926 856
rect 135094 800 136306 856
rect 136474 800 137686 856
rect 137854 800 139066 856
rect 139234 800 140446 856
rect 140614 800 141826 856
rect 141994 800 143206 856
rect 143374 800 144586 856
rect 144754 800 148008 856
<< metal3 >>
rect 0 106360 800 106480
rect 0 103912 800 104032
rect 0 101464 800 101584
rect 0 99016 800 99136
rect 0 96568 800 96688
rect 0 94120 800 94240
rect 0 91672 800 91792
rect 0 89224 800 89344
rect 0 86776 800 86896
rect 0 84328 800 84448
rect 0 81880 800 82000
rect 0 79432 800 79552
rect 0 76984 800 77104
rect 0 74536 800 74656
rect 0 72088 800 72208
rect 0 69640 800 69760
rect 0 67192 800 67312
rect 0 64744 800 64864
rect 0 62296 800 62416
rect 0 59848 800 59968
rect 0 57400 800 57520
rect 0 54952 800 55072
rect 0 52504 800 52624
rect 0 50056 800 50176
rect 0 47608 800 47728
rect 0 45160 800 45280
rect 0 42712 800 42832
rect 0 40264 800 40384
rect 0 37816 800 37936
rect 0 35368 800 35488
rect 0 32920 800 33040
rect 0 30472 800 30592
rect 0 28024 800 28144
rect 0 25576 800 25696
rect 0 23128 800 23248
rect 0 20680 800 20800
rect 0 18232 800 18352
rect 0 15784 800 15904
rect 0 13336 800 13456
rect 0 10888 800 11008
rect 0 8440 800 8560
rect 0 5992 800 6112
rect 0 3544 800 3664
<< obsm3 >>
rect 800 106560 146359 107745
rect 880 106280 146359 106560
rect 800 104112 146359 106280
rect 880 103832 146359 104112
rect 800 101664 146359 103832
rect 880 101384 146359 101664
rect 800 99216 146359 101384
rect 880 98936 146359 99216
rect 800 96768 146359 98936
rect 880 96488 146359 96768
rect 800 94320 146359 96488
rect 880 94040 146359 94320
rect 800 91872 146359 94040
rect 880 91592 146359 91872
rect 800 89424 146359 91592
rect 880 89144 146359 89424
rect 800 86976 146359 89144
rect 880 86696 146359 86976
rect 800 84528 146359 86696
rect 880 84248 146359 84528
rect 800 82080 146359 84248
rect 880 81800 146359 82080
rect 800 79632 146359 81800
rect 880 79352 146359 79632
rect 800 77184 146359 79352
rect 880 76904 146359 77184
rect 800 74736 146359 76904
rect 880 74456 146359 74736
rect 800 72288 146359 74456
rect 880 72008 146359 72288
rect 800 69840 146359 72008
rect 880 69560 146359 69840
rect 800 67392 146359 69560
rect 880 67112 146359 67392
rect 800 64944 146359 67112
rect 880 64664 146359 64944
rect 800 62496 146359 64664
rect 880 62216 146359 62496
rect 800 60048 146359 62216
rect 880 59768 146359 60048
rect 800 57600 146359 59768
rect 880 57320 146359 57600
rect 800 55152 146359 57320
rect 880 54872 146359 55152
rect 800 52704 146359 54872
rect 880 52424 146359 52704
rect 800 50256 146359 52424
rect 880 49976 146359 50256
rect 800 47808 146359 49976
rect 880 47528 146359 47808
rect 800 45360 146359 47528
rect 880 45080 146359 45360
rect 800 42912 146359 45080
rect 880 42632 146359 42912
rect 800 40464 146359 42632
rect 880 40184 146359 40464
rect 800 38016 146359 40184
rect 880 37736 146359 38016
rect 800 35568 146359 37736
rect 880 35288 146359 35568
rect 800 33120 146359 35288
rect 880 32840 146359 33120
rect 800 30672 146359 32840
rect 880 30392 146359 30672
rect 800 28224 146359 30392
rect 880 27944 146359 28224
rect 800 25776 146359 27944
rect 880 25496 146359 25776
rect 800 23328 146359 25496
rect 880 23048 146359 23328
rect 800 20880 146359 23048
rect 880 20600 146359 20880
rect 800 18432 146359 20600
rect 880 18152 146359 18432
rect 800 15984 146359 18152
rect 880 15704 146359 15984
rect 800 13536 146359 15704
rect 880 13256 146359 13536
rect 800 11088 146359 13256
rect 880 10808 146359 11088
rect 800 8640 146359 10808
rect 880 8360 146359 8640
rect 800 6192 146359 8360
rect 880 5912 146359 6192
rect 800 3744 146359 5912
rect 880 3464 146359 3744
rect 800 2143 146359 3464
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
rect 65648 2128 65968 107760
rect 81008 2128 81328 107760
rect 96368 2128 96688 107760
rect 111728 2128 112048 107760
rect 127088 2128 127408 107760
rect 142448 2128 142768 107760
<< obsm4 >>
rect 9259 2347 19488 107405
rect 19968 2347 34848 107405
rect 35328 2347 50208 107405
rect 50688 2347 65568 107405
rect 66048 2347 80928 107405
rect 81408 2347 96288 107405
rect 96768 2347 111648 107405
rect 112128 2347 127008 107405
rect 127488 2347 142368 107405
rect 142848 2347 144565 107405
<< labels >>
rlabel metal3 s 0 5992 800 6112 6 addr1[0]
port 1 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 addr1[1]
port 2 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 addr1[2]
port 3 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 addr1[3]
port 4 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 addr1[4]
port 5 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 addr1[5]
port 6 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 addr1[6]
port 7 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 addr1[7]
port 8 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 addr1[8]
port 9 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 addr1[9]
port 10 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 csb1
port 11 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 dout1[0]
port 12 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 dout1[10]
port 13 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 dout1[11]
port 14 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 dout1[12]
port 15 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 dout1[13]
port 16 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 dout1[14]
port 17 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 dout1[15]
port 18 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 dout1[16]
port 19 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 dout1[17]
port 20 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 dout1[18]
port 21 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 dout1[19]
port 22 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 dout1[1]
port 23 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 dout1[20]
port 24 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 dout1[21]
port 25 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 dout1[22]
port 26 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 dout1[23]
port 27 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 dout1[24]
port 28 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 dout1[25]
port 29 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 dout1[26]
port 30 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 dout1[27]
port 31 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 dout1[28]
port 32 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 dout1[29]
port 33 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 dout1[2]
port 34 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 dout1[30]
port 35 nsew signal input
rlabel metal3 s 0 106360 800 106480 6 dout1[31]
port 36 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 dout1[3]
port 37 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 dout1[4]
port 38 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 dout1[5]
port 39 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 dout1[6]
port 40 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 dout1[7]
port 41 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 dout1[8]
port 42 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 dout1[9]
port 43 nsew signal input
rlabel metal2 s 115202 109200 115258 110000 6 io_oeb[0]
port 44 nsew signal output
rlabel metal2 s 147402 109200 147458 110000 6 io_oeb[10]
port 45 nsew signal output
rlabel metal2 s 118422 109200 118478 110000 6 io_oeb[1]
port 46 nsew signal output
rlabel metal2 s 121642 109200 121698 110000 6 io_oeb[2]
port 47 nsew signal output
rlabel metal2 s 124862 109200 124918 110000 6 io_oeb[3]
port 48 nsew signal output
rlabel metal2 s 128082 109200 128138 110000 6 io_oeb[4]
port 49 nsew signal output
rlabel metal2 s 131302 109200 131358 110000 6 io_oeb[5]
port 50 nsew signal output
rlabel metal2 s 134522 109200 134578 110000 6 io_oeb[6]
port 51 nsew signal output
rlabel metal2 s 137742 109200 137798 110000 6 io_oeb[7]
port 52 nsew signal output
rlabel metal2 s 140962 109200 141018 110000 6 io_oeb[8]
port 53 nsew signal output
rlabel metal2 s 144182 109200 144238 110000 6 io_oeb[9]
port 54 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 io_wbs_ack
port 55 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 io_wbs_adr[0]
port 56 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 io_wbs_adr[10]
port 57 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 io_wbs_adr[11]
port 58 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 io_wbs_adr[12]
port 59 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 io_wbs_adr[13]
port 60 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 io_wbs_adr[14]
port 61 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 io_wbs_adr[15]
port 62 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 io_wbs_adr[16]
port 63 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 io_wbs_adr[17]
port 64 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 io_wbs_adr[18]
port 65 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 io_wbs_adr[19]
port 66 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 io_wbs_adr[1]
port 67 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 io_wbs_adr[20]
port 68 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 io_wbs_adr[21]
port 69 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 io_wbs_adr[22]
port 70 nsew signal input
rlabel metal2 s 108762 0 108818 800 6 io_wbs_adr[23]
port 71 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 io_wbs_adr[24]
port 72 nsew signal input
rlabel metal2 s 117042 0 117098 800 6 io_wbs_adr[25]
port 73 nsew signal input
rlabel metal2 s 121182 0 121238 800 6 io_wbs_adr[26]
port 74 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 io_wbs_adr[27]
port 75 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 io_wbs_adr[28]
port 76 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 io_wbs_adr[29]
port 77 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 io_wbs_adr[2]
port 78 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 io_wbs_adr[30]
port 79 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 io_wbs_adr[31]
port 80 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 io_wbs_adr[3]
port 81 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 io_wbs_adr[4]
port 82 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 io_wbs_adr[5]
port 83 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 io_wbs_adr[6]
port 84 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 io_wbs_adr[7]
port 85 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 io_wbs_adr[8]
port 86 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 io_wbs_adr[9]
port 87 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 io_wbs_clk
port 88 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 io_wbs_cyc
port 89 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 io_wbs_datrd[0]
port 90 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 io_wbs_datrd[10]
port 91 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 io_wbs_datrd[11]
port 92 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 io_wbs_datrd[12]
port 93 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 io_wbs_datrd[13]
port 94 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 io_wbs_datrd[14]
port 95 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 io_wbs_datrd[15]
port 96 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 io_wbs_datrd[16]
port 97 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 io_wbs_datrd[17]
port 98 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 io_wbs_datrd[18]
port 99 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 io_wbs_datrd[19]
port 100 nsew signal output
rlabel metal2 s 19062 0 19118 800 6 io_wbs_datrd[1]
port 101 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 io_wbs_datrd[20]
port 102 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 io_wbs_datrd[21]
port 103 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 io_wbs_datrd[22]
port 104 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 io_wbs_datrd[23]
port 105 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 io_wbs_datrd[24]
port 106 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 io_wbs_datrd[25]
port 107 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 io_wbs_datrd[26]
port 108 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 io_wbs_datrd[27]
port 109 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 io_wbs_datrd[28]
port 110 nsew signal output
rlabel metal2 s 134982 0 135038 800 6 io_wbs_datrd[29]
port 111 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 io_wbs_datrd[2]
port 112 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 io_wbs_datrd[30]
port 113 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 io_wbs_datrd[31]
port 114 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 io_wbs_datrd[3]
port 115 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 io_wbs_datrd[4]
port 116 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 io_wbs_datrd[5]
port 117 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 io_wbs_datrd[6]
port 118 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 io_wbs_datrd[7]
port 119 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 io_wbs_datrd[8]
port 120 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 io_wbs_datrd[9]
port 121 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 io_wbs_datwr[0]
port 122 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 io_wbs_datwr[10]
port 123 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 io_wbs_datwr[11]
port 124 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 io_wbs_datwr[12]
port 125 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 io_wbs_datwr[13]
port 126 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 io_wbs_datwr[14]
port 127 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 io_wbs_datwr[15]
port 128 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 io_wbs_datwr[16]
port 129 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 io_wbs_datwr[17]
port 130 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 io_wbs_datwr[18]
port 131 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 io_wbs_datwr[19]
port 132 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 io_wbs_datwr[1]
port 133 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 io_wbs_datwr[20]
port 134 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 io_wbs_datwr[21]
port 135 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 io_wbs_datwr[22]
port 136 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 io_wbs_datwr[23]
port 137 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 io_wbs_datwr[24]
port 138 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 io_wbs_datwr[25]
port 139 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 io_wbs_datwr[26]
port 140 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 io_wbs_datwr[27]
port 141 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 io_wbs_datwr[28]
port 142 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 io_wbs_datwr[29]
port 143 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 io_wbs_datwr[2]
port 144 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 io_wbs_datwr[30]
port 145 nsew signal input
rlabel metal2 s 144642 0 144698 800 6 io_wbs_datwr[31]
port 146 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 io_wbs_datwr[3]
port 147 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 io_wbs_datwr[4]
port 148 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 io_wbs_datwr[5]
port 149 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 io_wbs_datwr[6]
port 150 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 io_wbs_datwr[7]
port 151 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 io_wbs_datwr[8]
port 152 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 io_wbs_datwr[9]
port 153 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 io_wbs_rst
port 154 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 io_wbs_stb
port 155 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 io_wbs_we
port 156 nsew signal input
rlabel metal4 s 4208 2128 4528 107760 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 107760 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 107760 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 107760 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 107760 6 vccd1
port 157 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 107760 6 vssd1
port 158 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 107760 6 vssd1
port 158 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 107760 6 vssd1
port 158 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 107760 6 vssd1
port 158 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 107760 6 vssd1
port 158 nsew ground bidirectional
rlabel metal2 s 12162 109200 12218 110000 6 wfg_drive_pat_dout_o[0]
port 159 nsew signal output
rlabel metal2 s 44362 109200 44418 110000 6 wfg_drive_pat_dout_o[10]
port 160 nsew signal output
rlabel metal2 s 47582 109200 47638 110000 6 wfg_drive_pat_dout_o[11]
port 161 nsew signal output
rlabel metal2 s 50802 109200 50858 110000 6 wfg_drive_pat_dout_o[12]
port 162 nsew signal output
rlabel metal2 s 54022 109200 54078 110000 6 wfg_drive_pat_dout_o[13]
port 163 nsew signal output
rlabel metal2 s 57242 109200 57298 110000 6 wfg_drive_pat_dout_o[14]
port 164 nsew signal output
rlabel metal2 s 60462 109200 60518 110000 6 wfg_drive_pat_dout_o[15]
port 165 nsew signal output
rlabel metal2 s 63682 109200 63738 110000 6 wfg_drive_pat_dout_o[16]
port 166 nsew signal output
rlabel metal2 s 66902 109200 66958 110000 6 wfg_drive_pat_dout_o[17]
port 167 nsew signal output
rlabel metal2 s 70122 109200 70178 110000 6 wfg_drive_pat_dout_o[18]
port 168 nsew signal output
rlabel metal2 s 73342 109200 73398 110000 6 wfg_drive_pat_dout_o[19]
port 169 nsew signal output
rlabel metal2 s 15382 109200 15438 110000 6 wfg_drive_pat_dout_o[1]
port 170 nsew signal output
rlabel metal2 s 76562 109200 76618 110000 6 wfg_drive_pat_dout_o[20]
port 171 nsew signal output
rlabel metal2 s 79782 109200 79838 110000 6 wfg_drive_pat_dout_o[21]
port 172 nsew signal output
rlabel metal2 s 83002 109200 83058 110000 6 wfg_drive_pat_dout_o[22]
port 173 nsew signal output
rlabel metal2 s 86222 109200 86278 110000 6 wfg_drive_pat_dout_o[23]
port 174 nsew signal output
rlabel metal2 s 89442 109200 89498 110000 6 wfg_drive_pat_dout_o[24]
port 175 nsew signal output
rlabel metal2 s 92662 109200 92718 110000 6 wfg_drive_pat_dout_o[25]
port 176 nsew signal output
rlabel metal2 s 95882 109200 95938 110000 6 wfg_drive_pat_dout_o[26]
port 177 nsew signal output
rlabel metal2 s 99102 109200 99158 110000 6 wfg_drive_pat_dout_o[27]
port 178 nsew signal output
rlabel metal2 s 102322 109200 102378 110000 6 wfg_drive_pat_dout_o[28]
port 179 nsew signal output
rlabel metal2 s 105542 109200 105598 110000 6 wfg_drive_pat_dout_o[29]
port 180 nsew signal output
rlabel metal2 s 18602 109200 18658 110000 6 wfg_drive_pat_dout_o[2]
port 181 nsew signal output
rlabel metal2 s 108762 109200 108818 110000 6 wfg_drive_pat_dout_o[30]
port 182 nsew signal output
rlabel metal2 s 111982 109200 112038 110000 6 wfg_drive_pat_dout_o[31]
port 183 nsew signal output
rlabel metal2 s 21822 109200 21878 110000 6 wfg_drive_pat_dout_o[3]
port 184 nsew signal output
rlabel metal2 s 25042 109200 25098 110000 6 wfg_drive_pat_dout_o[4]
port 185 nsew signal output
rlabel metal2 s 28262 109200 28318 110000 6 wfg_drive_pat_dout_o[5]
port 186 nsew signal output
rlabel metal2 s 31482 109200 31538 110000 6 wfg_drive_pat_dout_o[6]
port 187 nsew signal output
rlabel metal2 s 34702 109200 34758 110000 6 wfg_drive_pat_dout_o[7]
port 188 nsew signal output
rlabel metal2 s 37922 109200 37978 110000 6 wfg_drive_pat_dout_o[8]
port 189 nsew signal output
rlabel metal2 s 41142 109200 41198 110000 6 wfg_drive_pat_dout_o[9]
port 190 nsew signal output
rlabel metal2 s 2502 109200 2558 110000 6 wfg_drive_spi_cs_no
port 191 nsew signal output
rlabel metal2 s 5722 109200 5778 110000 6 wfg_drive_spi_sclk_o
port 192 nsew signal output
rlabel metal2 s 8942 109200 8998 110000 6 wfg_drive_spi_sdo_o
port 193 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 150000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 35449388
string GDS_FILE /home/leo/Dokumente/caravel_workspace_mpw7/caravel_wfg/openlane/wfg_top/runs/22_07_11_09_37/results/signoff/wfg_top.magic.gds
string GDS_START 1343554
<< end >>

